��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"�ԕ�!p0��A]2��X3�F/F��Z�`RVd?�lL+k;�E�(���U�ZvD����(�9�7��F�3�>Rd�v���"#�\�8X�����P�`p���k)W�1��z0Z���(v������.7OM8�2D��3�-�>�!�ռ��9�OTCb�ffR��SHpΜ�Y�������ve��fm�ߨ<K��v��x�5mz����1ǿ��ʀ+�t��.�����G=l#���H5��}^�y���t��$ٟ舯��*^�q:,1����l�SD[��{������C6���^TBS���n�s�ڝ�L�����2o5��t�R����0$�X�x�8ب��R=g�X��c[9�}�4�k��%R��_�S����Α�v��1�Q�S� �)\+�,�0�Hmʁ=O�<�����5�gtR@~�O�l��"�����檚S5��D�PBu�F?��CFn�X7 �w@�Pq9�Ɖ�]����E0�|I� ��q[��q4��N��y�7����IU���=��3e�R}��nM$V&]^i����.��9�#��Ѐ��]�T��rf95� �@�<�M}6���@)�m��#�1�y�6�\���g�~�����H[LA�`��L<�wB����чIz����Z���P������k�hN��N� '�j%�C���RPI�X�'ݬ5��ֆV����n�tG�F�K���4LE��0��U�It79e��{�V\Q��LȎ�P�S�d�Z,⁻�>���i&�Β��Ir�)��x�S�KE��$���û��L֜��5Ӱj���]pn�W�x+w�D. ��	�,u��xj�o�BW^1�/5��+f.P�;&�� ܔ���T$��>�h�v�_s7�MǼ^��`�i(����4��֡X��%+g+/��	��F�-�Hd�g�j)�>�L���hpy�+���mf����+��sJ.!Jԕ]PR�IK��(��^�Ǥї��X�*yih�����5^9_��	�Nbyb������K�^ H�R^�򨴉W9�b��Z��^C����߰	n��W'F�:��^���f�%-k�,-��l���sT���dTp�q�k7
�5~���S8�������15���h�P���=A4�=�I;���+���S��
��'���ʍ�.�AOC��5/Sy˰�x�iD���Ba��u�Hy����EM5�$U�5&�e����
�H���*	=/e��{����Co��&��1�v~=pQh
��AP���{#ތs�����ʠFW���o�\��*
�-+�A�죒NvA	�����V1[�A�}��C�UL���"�.�'#j�C�Su�j�T�z���Lp������6�)+���:�Y��u�qW"W�t=�a��!*�m��g�X ����t��W���.���F]����b�G���<��1]�G�c�AP�\�jڲ�����md[E��f�
,f��QXB�w�ΰܚ([?������f1ys	���(>�1���:�l��A-�IR;��G�\{�?����_��p�>V���ĳ+lC�)��b��G�	_(�U,�dV���Q�ŉ?�G��$P� ���(T�F��F������f�[ZT�92IQ����\��J��M�����k��0���uC��V��:�$Kb\�pݟz#=�6��wB�TdS�X�� �1w[���W�N��Fz~�����d����×YK��ǈ�H2p���U%;�A&J |��a�o��&�w#Rݲ=<�Y�{
2Ȕx�%a>
��<4֙1���s�r�s���A�.a��1�4�򂪕�����;q3������,��D�[�aɄU�{D�'ӫ�\�歘wa)��p���V�&���L��@�T�K�^��O���Qe�0e�K'�p)2w$��� s_Rr
�:�$���U�UF���ƽ)� �J�%�aJ'�˃`X}�n �^=ɃJ�U�^��3��9���;~NQ=0Մ�m��Q�m���*�ƭ �h%/�a<��䪑Q���r�2��o�p�<<&D[�O�h��������}A#Ot�� ��2+=�H�j�A���5�v6d����]Jr��'4"1�����w�ۏ��C�iRY�ʠ�����M�\k��_��j�{����
����P;}?�݋�Ș�7
W7�"�#웎��̤��"��\W��X��81�0�	#�J�����#^++O�S����y<�et�\!�C��9�ã���Tr2����H+@� *:'V��+��+��t�&( ީ;�H6�Tb�C~P�t��稜�]�_�n�F2WM�����X!��� ���f��t
���qajIu��; <p���D5aM!-m�8���]M'�ը	�"S��{С6>i` �$�ؑDxU�"����܁��y��hʶ}��Ph�?��ab�=mX{`�����§�M�L~�$�2dvݰ��WcQ��_��Df����Nx.�N��4��K����a��C�P��x�ŦՔrà�ۀf����+�l����2��^�d P�G���jE�m�a}7Em������\�!e̣Te?�6Ϙi-&���ãeｈ❻��24~��(�YN��Yݑ�=8���j,���e�Z�g+���x*��C��da{�����f"\�
	���V$u`K�[!�;��+��m��&�k���ySp��n ��J� �R��LMj��Vg|F���C\�y�(����w痒��_�7��>�r+���5����&����(�����m"��n7QN'I�6�.��[Aa���O��ҽzI�9� L qVl�MV�A�¶A.x��3j&����W�n�/��;?�C���#H�tʚa�4)�9�t��/��HH�{~6eu�5�l�S��|m�J�n�#Z�r ��6�s���^,u���eČ0Q[c.m,�RW��7FB�А�
�{Eg�[3+�%�Ҽ�W]5 �s��Yr�I�q��[i4��yv�!w��k)�oz������c�T��I50�ޅ2�N�g��I�\C���:)�����g�����P�U\�*�H~Kf!
�{Y�����͒�Ƹn�uPI��	ϱ�g�ѷ�}E�g/(+�ńO��{�Y�я� #?-W�(��v�#��0<-"�۪�V��A����Vwo�0�+�����V�<\���a=b�10B�c;O�A-�1u�^ެa�d[/��횟���ڮ��Q`ev,Ȃ�4��2<��)����=�Gl�O��z��]��D@<(�&�� j�)y�be���
���@:�t��x������.���H	x6���`{f`S���NH<L7;�1�!��H��>@�tJ�QnW��F�d���r!���{����l��U������	�˪ج�����qD$W��p�SaR�?��7��V8KI�(9 [w�\�5e�Y�V�R����<�f=n܃�)�i~�����O�������R�**��+�<Nq52�X|��ݰT7Fze./t�1^FrO��@�C�:����[�M%�V��d��x���c�"��g}~-��������ɣ2��|�߰�#t�4�/�h�?;j� 0�	dp,������5�W��R�!4%,lc����m�MM�˽�jІ�Y���˲��-�/5�&���rՇm�z�|�:ө�vה4 t~ !Bt֙jo��~h��X!y� 3���B�faIǢ�n��?Y&�W�@�q�s�<�'��˱@#o��-��{�/�1��9Z�X����y.2���N��;�e�톹��"բ��eQ������Ob�%'t[H��2=���֤�or������5�?f�3�u�镢c��hǫۏ��H`��]��,�-;|)'{Qhw�ɩ��m�*�V���P�8`�6"y�.�����B4ڰqbXIq��D��;%u8jD�&Ԡ�
��4i���$o�j�_W�:�a��"b� d�ra���6�Bu&���F�4����{�k/�����M�Y����ۓz��:�b
8��u|KB����p��:5�LW��}3&�$ӊ�E�R�-v�������9/ђ$�߉yj��|]/��r�.,:�& &IF+!]o�.�!�x�|I'Sw�f^.�v�5���m�Ք��e�V.�Ax�H�q�＄͙�"�*��oͤ��;7j�Ί��F�!L'�f��@ �q����è�j�^���Ҹiₖ|�_!;�r�"��Ɇ�A�z�����kg�V��6�BU/�" ���Q�,s�|����nآ��$���n��#IT�\�Wm/H��"gzo���(���]`)�Ν$]gX)6�S?Wzf����K�˷y��Y�mlfY�QZ	I}�#�)��W;��d�A�R6��ᄢ1�(�����,�x�7ͤ(�C"���Ye��,�O���"����yt+�4��@����n�/�-�8�0�%s�Ґ��y�{*�nF�E#���G��P���R¬Z�G���x��E�C"�L�Vo���P�����N��X��?�Gp���=��� ȋ�.�
����F ���J�O�:����X��/,1�!��v���� $�*AV���h�M�y�*+m�gr����4��s���g���|c�R�.u<Y���ԍ��+}E�$p{"���Ę�[����;D1e��v��o,AL]D��2�_u;njQ���MR<v:�3V�5�9�"����M@��6&wT�2���`z�d�&+�����'0��X��z�)�@ɾf���U�y� ��[�3��n��ջ��4{�,�Ov�D<҃�Ɩ��i��lϡ�����Ζ��?O%UA��Q��3���Dr����:*�Yn	za�x]S$_���Y�����n�t�+�;�ry�	��{��}����i�t_3�_5׏�9��ph��x)�мeI;a!?]��=��5U4
�D�f�
���k9�\;%�f̚~��v��3������l{�/�DXx̚��j�M����Q~��	�s	�d1��Hu魈Ov��[ 25���i�7�vВyy��V!��%�&WW�/r�,2�T7�Ur!�- lɎ��b����W"t���;?�1�>*f��bx��a�2�����F��$p+42�*v�����M�b_Bz�@-�Ag��#��BS<(�g���N�0���6��iʆ�jC+?���dۺ�!��������ܷ�!m=*NkztAp�ep���t�_�2�.����#Hv��t��Z�WS#�\�c0/ߨ��+�!�X�x����.�E�3�J��S@cxS�pB4�-vn��?��J`��F� O���mTUc�L\ ��I��#�w{u��«_�0[	�G��ծ�6����2r���*�xl~�����/����N�,$ўw���<����P��o4��k//��.�}SK]$�Q(H����8�	"W�2s��^�v	N��편�؃��c�LI�g#��D�)2����ڿ���g�<�]#�,�N�H�� ��#鱂T�kBS;^�_/�,Ǉ��qjQ�&��c|�Y��@L�İ���^^�=)E�vͥ����k�Ֆ)# c�Î��DҜ^݇�c� O��T��*j��7���)j%WKz�6�F�wJ�'��\�����̤Ԫ�C@����±G���}J���^��0T�{!
h5�E�v�R ǚ) 4�g��*Y�;x*�%2b[{��69�����:��:l�]�u %�\%z>�t.,��uY&�SL׳1�in�LK�f0��~%�����ޮ6
�_���b�����O��� F�,:��9���bѭK[��龦0�&�B�AY�&��m>��YIg��H�z>��¤��Yoo��GC�O�!0���ה|H�ە�&I�����"����=
�z���iRz
R����6�b��կ�w(0��$�X�n��}C�W�`j�Ld
Ce&t�Vϯ	�	U���y�Z���AQoGX���T��-��_�~�"jY/��)�f��0�7��.C4��:���_�����@�������F��A���q����5�*�lƌ}�iɀ�F�9�6�n�n��?e%��e�jlK��Z6����|j��.M>��B/�/u�����b}��:�<`o�6m!���.���6�\oT�8iX�7(�d�)��9y�!��_2�j��\�Vr�1�F'ؿV�+rG����وo6-������e��r��|�+y.���ab�=?B�u��+n3À	A8Uc�2k��![��-l�ܷ��s���q�%6l���6�BOr���K4�P�Hn��!߲`)����1�I�oNxL���Y4~u��e�e`�2����W{*�ߡ��n`~_j�6+慊uTA ���������d����9�}�TfT�T�D�.+G�-�ꙇ��&�'�W����BLm�_�(S�i!|�<�%��[	�;Q��1���&��]Ets�����s-�mT|�kj*> C��v���jh��c	1~�����H���C ���h� ͷ����P�����l�5�U�z3�þq��y��9;Aux�jz�w�m�'��'�q���m���(���c#ۯ�ɃY����s�kޙ�,H)Uڼ"�j_��o��&�������1�dk=`�u@d7G�N�r���<.��Zڿi�H��e��5�{�Sܻu*&�W<V���t��ٓ��r-ԍt��o�aXN4.����v͝�qQ��@q	zzi��ʴ�|-���om��Ղ���y�U#�zHs�¹�I櫇%�w�]+��-(0����ʌ�d�w���=j�>@Hߓ�����{�z8Y2>
m8#��1�Ƚ���Ѳ��~��̅ӣ�jG�����گ\��$6LD���7Ϗ��p˕� �k<���tWAeVE+/:\�C����L��]�]1�]���gn��>kZ�ZKj���'��7[P*1Y�@t�UX�.�_��jrt2l)�I@Ό��I�UHU[���[�'��#˺��r��)�-���ܔ"��3e�署�Wh0�|��b����B�l��B>4�h�����%�j�-� e+�m(;K��:�:ר���{��d���ac܃�q��&Jf���*7��{�2L6��s�[�w]���{�z�g�'�h��H .a�����FQJ����V�e&�j+:��~����:��@E�RQ���E��#b
�H�������eiａ`I�_���ᾫj���M�6	'��N�}Ӑ�Em�$DI�~.����퐖(y��s��BC���q�W���dQ��?
�kj�|e�oW���ǜ�q��s)�-Mh�P���r9�����*�|���k���{&[gE���7��|��fl�Oq9� �"M�Rؿ�ʽi�\Z����������`@���9n-#h���f�4��v��k��n�̊�Ԧ��rd��ьa�k��rc�LI2i�C]��K��Ɂ���B���+�RҎNwiy�J�����kHZ�8V_�.���t����]c�2��L��b�#(���}g���N�Y)�DcU���[t''>�j��
�A�I@7���«eƺ���x�xu�ߘ5kpG6�:��E��NtY��X��Jh�;��0�[�� ���o���0�@�s��d20|"���Å�C��#����cS�LTJ�u��N6�n�% �p��UFe�;��j?`21р$X���Cߺ��Q�f+Ѹ�#p1
���M�w-��9=\�k���xn���c�|�H �a>I5>��~�Y�>��Ԍ�gg�G�R���\�����h���X 5�"}� �V���S��R"��^ Z�
���|'F�Ns��KC6��Ue���K��,�;5E�d1Lj���]{p����m��.S�~�����Vo{�{>&uv�L�W*}d�ڳ� ��Y8������m�/�i�y�YXJ��L�M�2�3G���ʬ�kF�id�nd�6Bnq?,��\���>�j�������	�9e'G2yu�c{�[{!(5�U]�7���S�k����o]���Z�zg^
^��|��S\�<��y��(x?���S�[*~���c���2~��ihtnF�D�&�}����3���os��_�'='�1M��;3*�^�}}mZ��W�J'Q�f�TN�nc����'Xz ���d�۷��j����
72���7����'S��^�;��Iy��C�P���M(ˑءV��:F��pxjȷ �����gN2F3B���r��wZp/|Y�|�a�ш�ʰ�}i���d�L�Jv����x]���G���nL��P�5�#�%��`�c���� �7���8��l�E�H�
����{3�3h�a����!N� : &E���)9b��<I2mx�n�f'~"_%"�.��h��|w��piY�7���˵O�<�,��lW�w�r z�&*��˥Jy1���.��w�C��Bm�7h\RE����gs�JB� ��l�������_�;�|�RAJ,��ƹ.��qJ,)Nξzs ��!�H����`FZ�@(TZ�����B'�� Q��̫�AV*뮊�w۟�m��"Yz�^ASa���hu<��t�3�W�_;�سiçx�↟q�$WmD�Lv��k!r&�Y�=�L� O�1K�;�D��Obu{t���H�	� &I�����F��^�udt��tF>�����y'�"F�FnsF_��ɺIN̈�G�.+�}��<?���� �P�j*[���6���sh��wY�T�;G��Ft�j������Fu#,��81K���Q;γl	�K�i"�n�+���R̊U>` �	|��M0�2�	OEofz	B�Iܫ�/89&c�!|�!�x�A���F[���ēyM�D{�! ���QC�P1szE��(M\��%V�!1����]FWSz{( y\��$��6�S+�
�\k0eҥȐ�X佻;k�Z�1tat�}ɤ����R�g�-З���O�V7���'1����c�w�d	�������skt�ȧ�����v]� ��p�t�q�1�D�?ߐQ�D��#���Nc�t)��Ȋ6(� ���r���p/�1$5'�q���S����z�����b ����Y�l_$ `�<Z����<�]������$��n߈�L�'�E&dq�ȁ^B�.�,mŮKu�c��(��ڙ-.�CK����F�����v ����#��M�F7������}����J��G^���o^�H��R�|ζ,J���E�X���\�����3J�w��)�Iގ8h�G*�wm+j/�o4i~~�n�"��Wv'�Ζ8׻�pS`�YM����zv�jn �M�m��p.ι�y�l�M�%�n��)��% cl�0+���o��m��65�����*�#`��Ed�$���d�hf�=����×u�&�aSv�V?���_⇬�(�8��	���؇f��eև]�Z�e�I�xr�g�z{����ᩖ��zG��G�r}�g�5Fڭ�..H�؇z���L�� b�zJ����AG���጖����u��b~j�f��t��e-3�耑_E�����!����7L�U*lȞ� �lg
��nx�S�ڡ�n�<�h�a��?HLP9�xj{an�zEݨT�ҁc�B��yx���V��m޼�%Im.�"�9���ќ�O�*ck\u��<��,�\G�-#H�;3� �7��3�.��Ԋ���(-��Ȍ��<3�7�>Tu�z��'V�m�ɮ����GT#�Z�|+F���#ȧ�s��,��� �l|Q���Z�tm	��f9Xf��5�r\�祯��}�����!o���� ��5�YҤ^��1sQ+l{8[WJ��l�i�nR���˦����7��v�:%�I�#��4t�bq��#��%��c�u��A)N���f3*u|k��`lQ�8���E�  ��qam\��ohCu�4��	L�p�ڦ�i�������P��S8���D�\4�V:�2+_)u�ɫP,�V��}%O��ݘs��I���-��Sj�nc�>�g&�Ԍ��� q'��r�*�� �-���/����2���B�b�U��D��.�v� �8��D��'\Q��<����35
���,�U+ i#��(e�lQ:/�B���+�I<q{x+��p��ʙ���BJq�7"��ݽk�Z�[M��_6��/s̑�!�4�O�5��$�Z�>u�c=��������<էޣ���evrQ$�#.A�5�{�I�^B�;蔨�Ш���U�ds�Ɠ�}o��Ƞ����<���+�Տ�j�3n����d�Z�N"�����v^.�)!�l��w�V?���N�kĨV�	].D��w�1>,�J�w�=?�l��Յcc�lN�l��x�pj���kR���F|�a[�ӰD���s�
1������s13����>J4�x����5���kN]����>���FH�w�~�=o����I&�`�hf//)��+����D����鷤��H���nw��g�ފ<"�w�oј���G�x*-�������@���?���^5ziJߑ���P�����9M�1��f���O�*�&Ů�l5�/���X�z_}Q$c�$:Ѿ2(b�<���z���9�����ڑ�Pm"+��Ɋ"�X��xy;����o1�}*�PQ�>K��mg� �5eCGD�Ǎ��H�-.X���1,�bM��v���0���'��)*2�mM3b���{�Rbk�:�9���r�ح�kķJ�5H���m�x%L�X��b��^	��7����*r�x��B3���f�X����0Y�w5����C��*e�t��0:ÃUnQ�jD�i["������]�����"X���	7�X�Hg�U�JR�4�'\�1�/U&�`S�F�|ɉ�4w؀����N��9����>��\����; ����\��-dg{�5>}��4��A�x�ͱ�����$�U�-��J�yG���gd�#�+Y�77�Q���
ۧ09
�ܷ�
�E8���7�T��N�nۜJ{C�%1Y���J��#�ִ=�8�"�=d9�r���Kɝ�y�������B71��A�U!����& /P�2���)�`�$+�1�bxlm(j��jL�f�fIv�J�(k�W�:E�{5 ^�Zt{�5�55�B	y�-�Z�����u�%B{�2 ��n�b:�bȭ��_ªDƗ�L�|X�|-�TN\���"F{��?�q����گB��oue��]�|���4y�\�	VL��fዣ�7�uM\.Y��{��"�)n�S������r��ƅ�6�E�����j��E�r�+ڿF$D��OQQv�P�,�lHeR3y�1��+�f�r.�ɪ|��-
l��;Um��;�"����b����۰��� |�4��J/�>�����mV Y(���\���.�{x��d|7uZ�������Ě͈�`�L^&\���&ۃI�2�D��Ke�j��'O���0s怫41�,6T����V�}�3)
��͢7��T/�̀��pL���>����A5�]�-�Y���Ϸ��G����Ek2�
i� Մ�?����.)��ge�+���|�gT.�i�i���8��9oo&��e��-Ƒ' ��yQK7@��6���&M#�4e��U��"ͮ*�r���` ѝ3�ϭ���`L�۾w�J����+X~����'�Ed��Q�%�X��de�(�Ó�3�l����Q]���6�Pz���`�N�u��������P]Ț�~ߤxC��[i��t����԰��o��[����ɖ�KY�L�,�4��A1 XTM��!Pg��9�W��Ð��iC:ClG8���������ȗ&��/V�g$9�h]JX�u����m�_|16'W��d�������4�y�&rS�f^��D��݃\  }��h!Gu�-Gm�"2�?&
�KۺH'�m>_*�
������>�G���G�'1z���@}w��Gt�ɋV���t�!jX����J���	�Y��/ѭ�� ����唎ʙ���G~��k���U�n$~�#1��u�	}�T)�^�� ��A�ž�d(�QL�J���8���<�3!��{孪�����yZ<Kw�f<B����}��a݈�74���N:� � �w��G�+ ���y�^�V�	���.ɰ���i��d�t?�&�ҷ7�Fre�p��Ebbg�J��^S.7�i���o�`��>��B���4ǂ�'�pk[�e�>TY�_^m,���P���TRs��X�򡬅dW�K�3\�x�*��^܋���H��7�;�F���4JI��Ū��<J��A�F��<��Z���Y����Y<�R��6�|]_Ʒ�f��M++P-MN��[������)x@僢p� �{L�#��-W�e�j�4�����I��S���ۊ�.�Q������?`&Փ���}aj=Ȁ�
�����j-�9�M�Ȃ�8}�9���"��o�YA����*��[�c`�=�u<�/��#KDI_��';z�??���/�3fF���V��i��[*�P N�5ŵ������>��QMģ�����"ĺ%�F3�۰zB��/�yJ��-v1���႙��1�5���ǥ�f �F�#�v�r���D���uxpZ�3�"�Vk���@�!O~
�f��.���ڨ9�םu��3�m���� }c���/hPI]�,��z�ъ�f��;"�C��w#�S�6,������1�ʿ����jL��V��t�@J�k���m| �`e3�*H�N�i~�w�3�J��`�o�	���F�@���+��r��kj!�U�
����ڰ��q�1d [�h��D�+s�`?��C�/�xڛ�f_���˞7��!��3���֙�e���n�F�T7������	�4�넧�`��F�9��ɜ��Uo��f,�U�E�r��qm�N������sf����ZE�;�.����F����qE=�t����Ҹ��Xr;������4m���.�������ov�[�a���L��t6:*��(��D��h����8{@�ŇRU��6�����K�uAm���oq�� ���!� N±Á���c f�N�a�D�`����Ӯ�#�P:`̈N���#Ҟ��p�zÆ�* �T|Ģߒ�0��3�n����)��&✦��CfC�ėu�����]f��
��\�DIS�Ԭ��\�LD���hk&��i�,�cfh�Gd*f��f� �`���?��)[ό�Fڶ���F��2N�ʌ�CK���{Ϧ�=����\� �a^[�Uy��iLH�^�=������ţn&b�f��vm�[��XBZ���#�B�-©���낅���'K����֦�L��*�Qr�&�g���V��A��xs�V2���5ԍ~,e�)\1�z��GOJ�d�0�	f�yDtiw��z\F��e�M0~;촡WD�}2Z~~'y~X�AUZ�he�H� 9��>_�b�a�gh<L3dZ0N���5���Q�6Pcݓ�y|^�U�:���~ƿ�]S2�5�Pc��N���|:�W��a�s�)�`)�e������	A�E��DG�vf���,\�00�K,9-�@i����}��l��x��[/�I��֤(�|q�$ux-S�S&�����*����آ���Z
-�I���`+0@?@��1x����d�w*8��e��=��w=h'�&,q������c�f�\�,���������޼=SC�z"�N8�/�����nFgֲ��'U�{,��GJ��F�m��9C���FT�m:
3p����W��fY\Tt�r�H�#̛��,�	�R���ni�� �Ъ�
�[K��E�e�p��A�I'����$��2v-]f*mj�ҧ�,���a5�|����q}�I��Dk�.�*s���_�a�k��A\DzI4e��Ȣێ��M�5y��_�K�5̆����Jֹ��M#K�2c����{+}�#��n$��
���F�����7a8�GV�|$4��tG�w�'3
����j�7�3��~����,�WI�_��["���e��;�/�RN����"��F�΋�q�DP�.�=�ۼV؍�r����	<:%�LQ��?\WT���*�41���=���ݢ�/WRY�*,�b�bT����C�J��`��L���P�1�e���]��
�l$��X��zSXmj[�V� ��F��"ky~yS��o�x!�<Hs��\��ؗ��=bvW�+�D���+N�� ��b6��P�\�z�<j�ViO�#�G��/���j�br���@[�{�e���7�aL�H	�}J���� 	8�i+;	`�K���.b�z�x':۱$/����ŉ���!K�*Z#X +\rq3�im�/��������.��烺���K��r�]�>���r��~b["��.�ӳ!P�8�\O��E��G�
���X��:�.�A�00�����cv�,c`�׷�4�)ܚ���/�?�kA%+�_z�����2���Ⱦ~L��m�����U��7n�T<�-[�����aN�RY�ɷr�t�~��,�Q�ԅ\�y����T�&OqS�>d$ٶ�B����b��L��÷���J��������팆�ˆ�GA^_�ᨉXY��6-����-�� �\�!�ԛ"C[9�����KA,���Vy̔�2(3��ec���)�MD)={*�W!峻�S�����=n�;|��e��_����ԣ���K���-�Ԫ�����(��}�b�����K���n��غ��Wy �fY}
-5������xzѹ��N�I+���Y��S���[���Fy�`���gi���L�oE^8[^���ow����Q��7��F�O��X�6���-�lj���$^#�kf�/�*7~?���Zr]x�48v:.=��iX��b�<��&<Cȣ��H��1�����|s�U�x���.��;ќb��`%��dL�k�h@0xD���Z��HW]2?�z�0>>������\?�jԉ���{	�6�1l���l=���e��N��N�߮ �����|Y#I�_��:��9����?��و�`WU�t����^���2���E�?��Ն_�שG���u�m�K{��QRy�h�w�¡[_�����`X��f�>R��su(����\�e�kX��0���߾�te�]��F�䤿L����jiR����Y
|��G�@*�Bt&R.K~Ϻ��t��5�8��TV���"��)��ĥ�Vd�$1޻z!��Տ�l��AE ��{�\��P���i�EUﬄ����	�ۜ���"��e���l��t	C��.A�4�r��0��W,��y�rf� ���N��c��ۀ�ڵ�;<R$ vmuFQ'T�n��q[��������ڳH��G�H�S�t�Qdf�
���`i,-��a8C>t�R|�`F��_�Ci�C9�p��~4�&w�=xG ]$���{wz5%��!9оAʓ_����l�ȱ��N|u>��ø�Q�_�\-@�>�*8nz�eW�ɽu�W�J}�U���r۸h�D������dϜ�T�\h�����m�`�N�A�d�W����4���-��M�<��{�e���W�z�����ȫߠ�r|����G����'�M�1�3�5�V��`��|C��?WŔ��Io�\�Q��v���v�Iu�����R��E�ź���W���]
hV����M���04 D�G�t�>V�+R�R@嘃Ǝ�����#"�<(�N�bb5}��|J��E�t.�
����, ��@�Up�\�T�\ۗ2��`�p]���Ooiڕ�ܼ����H�H����u��G��[��85Gl��Ce�~�\�1[�`�Ŀ���^�`r���jmz�օ2zRdw@�
���
@�d
,�W�9��o}�XM��Z��c�R�njm��PR��C��kL٣��̠u��%��t�̈C���T���I�����/d��R��۟C����\W�)X�fU��^�@�*LY���W?1�жAs�Z�s��a���	���
+g��.�! (�;� V�	����ړ0��%�Y�=㡰ŢpJ�G��N�e�9����{�p�
f|��k�i<�(J�vB�?J���P�-��8�űȉpۃ5x�c��-���s�30�Ѥ��T:Ntp�*,,��ߨ��f9�]B����)8�+b�|�Ĥ�J|7���#�<��Q�j������t���֔Ѩ��F|�R�2�ug�2��\gGȋ0'���������_�]/���S��wK�/�JR�Yʟ���M�B���Gs�T��H�
��6�@l}�=�JeB}v1l_<n���M��r���,ϪI���xMXS�Q�ʘ:�G�Z���#ai��P(��;�WH��n;�\��:5���ZU����p�	�e�����)/��s�+^����V�J��V6�����O �h��#�f��}��@�^�{8�H�6w��cd�<�=_�1ڭe�2V�e�++�����$�@*�xg �5m�Uo�=�s�N��W�TB�Ɩ��eVg��w�%3|1��3c�<s 2��K��C�Mp��zF�EBJy����&C�'.f�ϳ�+��_����q��R��_%W���}n,<�fhҖ��"o,����� |{�F:{�j]����X��T+9`�>��g��_�l�[�����V�nɟ�|r=eտ�ʺP����(���~P��XS>�����跲/�ī8�w/_�JF&D�	A��ڠ�AxS��9	�%���ŧu\m��1Q]b�UQ n�	[m3RO�Y�!���+�$Ǹn@@f�f���Ǳ�."��x�1&`TR�1QR��!Y�sC\N�4w�ju�e5�;_��W�e�8����0�tQӚu���`Dr�H�4_u�K�~�X�s���/ٖ]���͆�E9�������!;��ug�Y�H-��Ώ��6���5��UB�B}a"�p�����FD�6��MiF+D�8����X�k��aB}�|�-)O熢0M����:��L�ķ���/8p�9�d��(1�ʏK�|���$	��#�Ͻ�u^�ڳ����,�~TNlg�q8h�NȆ�����&8t:�0��UJ�taz�>�K8OQ)q$^{ ^���G��Q�0�� �5�˸�2p��U��`���&��͘^��D0�TS�\�u��N��L
�_���mCEs�!gAm�'ǫL �B�~�Z�
�����2���5C��==ո[o�}M��m:s:<�?�ir#�f�S=
}�z�Q�B��i��PԹ��"LO'.tc�3K}�f�,o�($x�ɿ����k�dݡ8֯��џ@�I�� ��]��Pҳ~����ş�P�Lt��hi�h���?�>*����,U��ԏHa�֭�,hu�.��C�[�r�,71���ɀ6�m����f��Q��MO���BI��y�3[��9&;�$�vn�ىQI�H���_:G��g{
�fH=�G�����[co��-�Aj�4.��7��q�-޶`���;D�
"}��L܀0?��'�XՔ�в3�]���(�k���oq�Y��K����d��!rz���<P/y��ZN ��E<�i��]RbE��F���=�e�
���7	p�@�d��k]���2�>���� 뙝$,ӝ/���\!��܌L���.�`��=cˆ�h�,R�E�bS1���Ӿ�,�
�[`���3y���U��Y�Ó8@�WOȿ�ѷ�q���M��"��2�D؁�0[���.!8�@���K������/�w�����끵�\��{4M�[�D�����d�%{q��DJ$�lݴi]���
�[R%%���Z����$�vI@+%���.���л�1,��2ށ�3t�%�&}	)Mt���g���6@��_9���xr���r��cx$5mH�:9����ƾx��={�Y���LK�M{|4��G[N�r	4��2-�A�nJ��@���QH���t��o�����
T�8��NT2vW.�0D@��ə�T���&i졃�GH�l@0�q^���0O3j��;��^�ԯ���vꢿ����8~��bd;t���čS<>�IsQ�Y�����I~E�e�L��ؐ#� '���: -p]���xe��#����g��l�1���Q�6�6��]ו 7$j*l�U����=|��	��6�X���U�EXc�Ӌ�,�g?�+�ڴs��.Yi��y�)�AGTrM��E�d7��\7�9ȁ����O%�g�K���[e��yX���a��&>�\���P�VԔj� �N�E6�3Z	�Q`K^�ڱ�н�bARk��>��%eS�����Y���*�Rx��~�0�hUn��<�T�~|��1@!��`��p�*Jl��'�C�]waH����{��9���F
�B�2�R�M>5EK�ʬ:5��i1��6/��j+��7�}��dYd��x&��>M��>�����^��5`���+809����g ����6�W�x�623�}��:ڌ!W��"	�i���r�ί.d�b[ �E�������5Jf��Q�`����F�:K�i���� ���'��k�Ŷ��<�ZG�L�Ҹ���l��O���Q&a��TN%@�ߴ�n�;�9�H)��6׳��Lf3 ��!�ي�?��)m���Y�Y�m��]Z:Y��\9&�V�$�+[r��0{|���C2_$����&u�����1�N\)<���q����.��A8`UA��Vex.���(�$�>	,�!H=���$�C�s�9%Q_���;�fU*���x��-�ؗ	�)�7y�&�i`����Nx ~�̋�lrZ�ZE����o���s���P�H�D�����f����>�ߑ����;3��HP%K�zI#F;o��)Z�-C}��T���e�URzm�H��mx�A[Up�|��n��,ѿ۳�֓��t���gS�c殛-�J���V����Uo(x�I/��<�O���e����/~c�w�љUn�V�&*W������W
:$���/B�����"k߈2<۴��f�8��/Gk�H�$i�8;��m� ������zD ���y��E!)p �7����r�
܀�ݓ�'��Ӈ�� u��Gￄ���٫�����?�.���������}J��א��i��!!�~{%���aDDi�8��4���6���05\^���HHa`[;^o�~Gl��{���,{�	�If��ή�
���BM8h�Q�P'�}���nܣσ�z���G��@Ktz,7Bf��!����{�Z�tX�4:�z�fdA��(�B�K��+w'�ky���(������QP���5��U��YR��m��
2��w�<��A$��m��f|���8�G엿:q�^���}9�F�2����(���ʵ�~����L�3K=GD(3��N�.%�1���,�K�� �0��g(�u��fA�6�)]���J�c���i�m��u��E'��y&n1��<ҎR�1e��}�<������<�B�0)��#T�4�
ly/�U?"�}Hػ�y:?���^YW��٦D���F.̏�-�oY�I��)�U�W����ס[!����1��Wj�؃���g�Ԁrs�zq��� �|���?��F'�r��rU�w�7�!W �)� ,����y�HH��R�a�B�OY�4�@l`�)*�c�kZ��V,���A_:Γ�u\�7��8z:���K�]!�~�"���e��1��	�=���]�9���	5�mg��{k9lZ�E5��0/R��|����Zu[n��I������K�AB^x*��~tH�@e��P�?,�;0[/���ECO�N��r�.��	���&�G��$|�@��J��y����}"��(�n��T7n�Xt���0'#$d��|Z(G�������ӑbt�ų`��Qט.�P.1t�Q�i������v�=��P�U��mx$�p��%��MɜF�����_�'Ֆ?L�4�ʂG{���'�!�|��{!�.�.:d*����Yaboe �;E�|���1���>'�:�`�F��ٳ���=��So
�{�*��=\P?�@��ڄQiBE�����0�VV�.E�+6������ɢDI5��T���E����"<�0�S7�Y0�*��L�x�4�2�H˞�ǜ�I��;#?tw�v���������w�g�e!>W�9S�fE�X��L��"E�Ku���^�z�Y�]���M�]�t}�y�X���Fq�Ԁ��z�7܌Wm�5���o�/�����H�B�n��Onè|]�췁Ғ�F���d",
v��mtY��AG����}y��Qʵ�Ɋ>����j�rQ5@�G�R�W
�&�(�ʠ���O�j���:�R���D�^Zs�ޑ=�s�P�utl�"�3|�Q5�d#+�Z��sa`�����Q����
]{Ҽ����$�?��Q�]F���1c&H�{E,Q�0Km#��>� 9q״�2"o*�I�>&��G��sJ���(�R	5���,�z�����h�L�R��.�~{rk�	'���Yq�*�:��BF;5J���R̪X��7�����Ԙr�<��CM|��{ڭ���9�C8P�Q�;-��Oڥ�&sa�9Z��Ȳ2�d"�N�ne;)<U��J�?�]�4[ڴ�9v"[�E��bi�Ā��@hxU\��K���3|lȩ����P���!o7ʿ���H��]/bШ�؎�R}�����h����͎�g�.�i��R %@鏚�9 %�*I|,5^��7���%vq}�K ���-U(�~U�,���g��I6w�� J���F�����+�7)�O$��kWsQ��P����o����d�$���_b2��:ݘ�R���9kZ
�XjT���2@Ը�Qkd��v �ע���(zԦ��}�9����(vGu��ILp�q£ep;خy`�z��.!���b��X��\�<�w��au;�k�e."�+�"��'����Q����5��w��<��7$�������v	}]�6i�
�dt��ye������� Dy5���g���6V	|���;	��=dsPΐ�����9���1$3��m<!�J@&�km���$]������r4�u�A���O�GS�֊r,�D��Lp��'��Z��b��'a�����0ݠ�`[�e�x2l����?|C�"wO�'^�3*�QN��UKS#�P����Խ�����)X�70��������ɡ�����.J��` �~M�C9z��:g�v��͵M��;�j9ņE�\�k���.�����@&��& �%Xw���M�P�@�GX�D��e]̦�Y�4��}\��g[�1|��*����"Q]M`�z6'���VH0
O�/�(��) �P v���T�MDp��6v-�����ls�bDM�����5�/S;X:��5	��j��i�;Suy��sϩDz�0^�
��<v�I���~|�����3���J(rK���4Q���4�c��nܳ�p���ɥ�d�R�`Z'�ayln�
H@q�^�,S�-f���8��&��9xoƴ�F2n�����C.vi�k	�#m��"�KD�'8m�6ZhŦZ�$�u�Z*��*;����ū��.b��o�M_���S/��LR �j�(S���*��`�G�m8+�V�yw����f6y�6�i�Me�+>����l� -*Ef^2���*!)U 5��FCﾻ�퀶D�i&<e.})I�ypt���f)
F�P����(`͡}g�̆�_�Ez����K�EB��4=�O�Ȍ
\���c�]�FcƄ�-Z)�'�r�}\��~�`���A�t��X����$��&/Vd=I�kR�c�G��T@rc�$'Ag�vau)��
� �&���X2���fdpE��|��ƞ�}�&
}����Ą��γ��/����k��@�E8�:Nq��S\�1~��"�T� ���z���"��cJ;ٺHa��4>-����W��rl*`R\����%�!mcbE����^$v�@�����Y�`��
����%���������@	y�����䋊9�{3���]/՗�6�ˡ��[:�a�"u�dl����i-zRY9�]%�Pӿx�y��r�AX��T=�ۡ������EFɩ=R�f����ipvB�V�;�T1_-`$����,��ܾ8T�9�7��tl�~v��gI������m���p.��˥n�	���jwh�h��T��kQo��~+զ���t��l��R6 =|�p�]D<�����Jr��L��g����&�o^}1������N˶�d��-����|�|=�Ae�]����*�{/s�Z2&����R:Rki���Qfw���c�䃭jϡ��'�se���K2�F�-Vd�=y�5`�8�!��1U�)^R�Z����9�nb�O����w��#�,p)�#�Y$y�P��Fg[��C�c�4 Wʷg��r��v0Րsd�r�:ܦz1��VbY?�%_O�2�42�a��5�1`�@m�l*^ 	'�7�Q��1�+Y
���;z���ɳu�Z���Jni�jS�M"��f�S8�:D�I9�������Z� j힊<��Q��0w��㕀�7]�i�6�eS�
)�\lw�O���]/��ʀ��M��j���尾Iu?a��Đg��nqvG�[ݪ�a't!�]C���D�{�k��Pp���JJ샌"�
�	�TK�q}�A�Bv�))��R\���[�b�m7�V��v; dY��eFR����MZ\K��U�]�DX������ ����P�'����ESfik|R)���c�i���)��!\H�}r��k�KC�NW9��h��NC�����5�j�<G�0F�,�D3���8�QLZ�/en���P�������rO������Hj��N���-,I�{�JS_u�I
��G��Cʷ!O�b8X�f�d���v��ۇDO	\D��n����-�v��G�.M���X!?L
:�6i�eu��.H��+��Du'[�P���D�ձD��ss@$�	c�m@���@f��=����ΗNe.L�$�]M��^�	Q'���_����`d2��a�2K(-����/�O3QԸ`���\�g��5k�G�7�����p��n+OJpBܔ�6���ߘ�ĶR�́g�7j_!�N�P����2�P<懀��������M�DЪ�K`]��Q�jL�$7��q��4�]��Y�NT�!�/(�RU�F�w����Иէa�6Q��j�z&[�6:, �?�6��"O�LW.���#�����H���ϪHW�H��gO��]V��y�.�h���ݝ�&��P��V�Vü�2h3E��Y�@����p�]��s/B���d���/��X�c��_���<j�`h�0/]7����ٓ&Tr�I��%�;t��ﱴ�Tg��k�:�S��G;�Tsu�1/�����UtI��B��]U9�"]�Z�ȡ�� ]��b���ՙ1*�򯵌t;�+R��M�j�|�9����QM5ة�K��9D����"H�+��l�~��6w�Q�|���d�v�(�u�3��Ř��WzU����؉L��r��郿k!!u��N�9��r��ҳKX�W��� ����^�
xD9�4�������8<L���O��s6�=G>��9�w�e�3�G����|@��pB"��%>���8�X�fE�`�ל9�'Yx�����*�̫��)��(�Ҵ�R�1��!�	#�C�&^��8LH8�n���(쒐N����a��G�##�X^,)@;��:)e��굞;=��gjA'�`���i^���K�S�:��'�� ��?���'��z�̟�_�J�oE�X��ؗ�.�:�a�'򢋈a��������2�rkiQ�i��/0�}:���G�)8��[����u>�K�8� 2K��4K�JRj;߄)���	r��BsٹI�%m2��q�.Q����jF�.�~�7�)��c|_�E�w��&*/0H���X�-��2y�B���xigZ�� UU�Iv"�l���[�����v�y����-GG�����"hO�By+c�Iq�V����~��Vm��l͏6�?��nW�1�����_"�5�D���Q�l/+t�Tn	.�R�H�J�X'�rO�SBdP�7k��ѡ�� �ū����Fٴ�ͪC���Zn�Q0��;'4=��rL�SO��x	u$BH���h�Ȃ�7��щЌ���-TR���5�%�M|\I�{r!���ɗ��E�H�J��6�&5�����j������-G\SYB��n%�T..M��+����䜀��1�����_U;r����4ibԚ���h_�o�-Ac�1�_f�w�[t-j��}�{�}��k�� A�%Rm�U�Ƈ�K�TS#��ι��Nue~��/�˼@gEL@�U�Lؓ���q���,X��}9.o��� l�EƦ��v���<�/�f@�������ذl�3L��o���\?ޙ���)&���U��@�ŋ�B�Wm�^� �É��T@�ۑg{�lN=G�{R�V��T�5���{9�����*֨�9S/�qZ��n�7Iqc��{�,j� ��{����d�7���&�1��rb(*�.�&���^o��#�X���y��ܕ�d����,�>jK��N�1���в'}�1^�uN��z�T��q�|`�\�`:���mZ={͝1k���V )<��O�Pnp�wk�
h�,cC�f���^sK�s��g�*Q&ia�U���_��r�_!.��REK�J�>�u�3>��"���LhO�f���8=(��1�|�&J���f���\��w�N��y��f1�4�\���:ON|��k�(R#��X��g���_�r��7[p�S\��>;������<�S.�6YK�Ff�Bfc���*����᝘����S��'$��-�w��wf�M�D�o�ز���FeuA���; `T%�Xۿ(�{���!���̇�!گ_��#���34�X���
|:0���B%vR_N����F��K���WJ��f�,���!�mxVU��J�mrm�ה(�?������^�����);&]��n��?��%N�0d/&L��rS�=Q���-�Z X��W�ԌK���
���h��!Ѳ$��ƪ�%��*X�t�u�d3jw:����,��w#�;egG��R}������f��P�u�N���YFX�^��'��i������8\���X��!c/�͜�7\�x�t�'I�\����31���ޟ����wn��[�O�?V�U@9?>a!�kXo�B�`������C�li�����Ǡ��y�痡ER����:�� 	M ��H �������8�4ƮTec`��2�=�i��(������˲��?�uk��<�,b�;�6쾯�(#�ȝ�P&Z/	���E@d�� 0BH�y�S!�`��(3֧$<Y��O@&��=ڊ�'��+���%����l���.�~�<��� 8X^��T��a]/�� /\IF��n_��o �[,ɖ������cO������p�{�}X���K�t��/�t���vc2�,��M�]�i5.�bMbb�$�&WTv��	Ci�q<ʍ9���'�l�Zv�=�y�XS���#K�f��2`�b`u7�`�S� 2�cC�r��T���S�v��&�>�"E�`/��0��`�~Un�g��
��4���9m�:]̾h�����ُ[����3��_5}���VB]]`�;�	.�z7ng%��*�F>_��� ���T�U�o�mP3Prm�nٖ��R����D���f�eTC�̐���a�7�?N�0:�4�by��N���i�?(��U7��xڋG��^g��i4T��,1��,�R�L-�_J�L�ِ��T�����v�X�'�je|%U�3��O��>�|O�f*C�����N3K���t.��҉����D�<�׽����<8��1bOX|E��yp��p.t���E>�?����M~���,?@�x/E��+����vӔ�
w�b�V��_�ӀH ৥�r�:o<OɝDi��Y�%�DW!�i��
�п�؀�冩��@�E��@��S�v��<m����=J�;�J������HR���Dԏ���>�V[�-���?���͗�3\���������h�}�x/�Mʶ��T#��j]��E�z ��t����v����Md��p��r)W� yH�E���p��\#�5d�yU���\_���c��j��J�m�f'���� ��E6u{T����轠K����, U4������O�� 5�@|���&��$@�l������D�n������te��F|whA^�.��Z��á��ǭ|
�ʛ͇�/�0�c~ER���yׅ��M���T�*f�.aXN��4Lİl��$��2�oW+~S��Ag�>�d+x��o�u+�\����/����Ɇ��P�W��۲Y�M��I��l��]U��B�]Z��q��v����ϲ4׹h��Լ~h�S$o��|���T���ܕ�8�>|4ȜIQ��?"Z/�Y�S���Wz]#�ϰr�S�s3�� �׿�9��9>���C㾮DN|B'U�+8��7�er�4F�G(�wQ �����]�עC{� @�DOU2��*k��nS��p��3���E��6Ay���(�< f�� �7w�Pf�7�[Tw� �qe�&�d
�p��z�e��x�,����	�U��@o-��Ԓ6¡�%^{ꥲ�D�5'Nt�J�@_7X�!}ʟW��p��p��=MQ�w�g���S�f��	�Z�~ML{�W^�xq�A[��PH�(��%i�=�"��ȃ7�1_���7Ǳ�ub��#
�J~�Ȟ9��v���
�
�"e�K��@,�3�ׁWD�<3���7�s߹%9G73go{��a.2al&���˻KBo�4C����.��}�e@Qr��ߒ�=KygL�S`t�A�w�C��+��/G5�p����4�k���!�/��_�/.93s=*����M���)��h� ��B�����ώ��=��ǒ&0��؈���J�(���N,N�G���+�<X��4l�E?�h�����=�����WD`�
 �JFE��}�o~ݓs�$-3(���Ea:���#�l;\�1J��D���y�M.w��������t_:�Π�B�*�[Ey�BզXT0њ�u�ۗ����m�z�6�*���|��铡7�'8r?�YIsv_b�d:�͆��b�4����+��8����]�m����\6��8*A>�b����[$D��v�3���~Mt��H#�[���$P'��}�i;a�""�gA��`�*���i����=�qAv�������$�81�_�:�_�\�k 6W_F�_������6�Jɢ���J����
P�s^���ģ�/D���!<�	d�f�L@7������{�jG�C/�T�΁�cȴ�<�u ��I��d^�13�9�c��Te{�j��T��DX2z>���D�������8�V���^Ǡ�Fo���7k����+�]������R�J:)UGj��ݩ52Y�v7'ߌ�qe��1^�g*%�
)8؂��v�nUE]e��
� )��`!G�F�#fL�A&�v�TZ�˵�+U��e��(A��/��Fk�V��i����s������	9���� ;�Ş�i��Dd���g6��ۤ#���Eh.���M&��؄vAn�.��N~��Ozc�ufī�R�U!�3�:��r]5,`�l��?$�5wz,����o�"8m�.S�*
��
0^4�{��Q��_`��}���O�S�Q�G�����AZ&8�s�ݜP�Rw�s�2-դ9p�:��o�Ũ���$��U3rƄ:K��?=~c���__I�l��Ug�D��fQ�<����4\�����ggW������@����wM�"%�qվ �)��0��p�nf{��rv�'1Sr#"�ݾ��k��o444-��f���d<Q��/yC�!\j��-����Z�O��+ג���V��SB� rڱ,#�Q�=�hpz�����xv�Ō�f�����A��oF�AC�<I, -p�Qn���i/8膢�ZeI
2f�A�J�^�ţ4�D���`��,��&k�x�ߎ�^�5���d�O��}�6Fl����Ao��}�k�G�	b6�	+w.!x$"eRC_Y�	�k���b��ȫ#��e�L��W�|��m<�*���b�/�q�����g³Mc�Q��EG2/�C��؞�{�H���2L�i�S$N��5C�P1�@�cs�3{�oF��p�E���M��� #XC����9w���?�,�	1&.�PV���T��\�}|��qD���j�a1�6O%cFc�~�g sGx$�+�r�S�Ϝ��
�Iom������K��Wq̢x��f�je��?C��۾˹w���9�z>�{��Y�KL���&:X���{?�Ah(�~��Ws��Ȼs�~�/}"�rY��!�T�����C.�ǜР8���m�"dh!�o�|�[�E�e,�9tr���⩱ǖ<e�l�J��zls�N}V�|&/b��I~;4!O��79[���=���e:���Ln�5��,�<\Ut���-[�xv�zGq��`�ytL��0ϢD�n�d�`&H�Y�f��+���aN6|.�td��ռYKv�cW�_8cɢ��m;��:i�'�g��>(�z�C:���í�MtHn T��q0��tZ��p-�mL@O|s�C�_�=�T2P�◺:�=kt�~�ZG]��	V���a���E"�����T��}}X�,��m��K����v�H�����������ğ�����AX��|�J!������	P7~�.�P�2O0a�d��vb8#�"f��SC��-���zƱԿ�'����-%��Ԥ�b��ޢ��T������g�8��75U<�ϼ鏿�z�<�;�^H��еm�d6�����^��(�lո���O�H"��s�݊�(�[�^�T'U�)ڰ�1�@��H�}�����M�5M�a"V���&lj�;�lu0sB,�y��͹̢�*�ۡ��kq;��Y�~�Z8�|LYM�YA�\�����bL�j�ʕylhP(����H~i}���#���UEƎ
��L�U>�gO�;�(
I���5R�sS4�5^&v�s$��w���:��r�F�
g��e[^wHc�P�G`KF�b>������s��hZ4Él_d�	�r�5��$��}%)��l]|g��.W�ZL�xN�a��#"��o��+�r���`�|�Τ��d#��·�B�Ũջԧt���e�llAX����4=���N ?�s@�7�Y�Uu��a��9ʤ�1����ߞ��*��J5�
�)�gE��,��!b��ǘҼ��NeAq���\��
�W��ɤ#K��n����Zp��B�Ҹ�'�ځ{OHs�}��#��f�E�ܒ~qw\y���(��fU� �����QoR��V�ɂ�"�z7{_)H;M_"�J��@䐺!�4���2�]�QF����4n' ��4��d�L���F�~�8�m
�uΧ?�_< DHj��9���1�1��n��T�v����|+q�e�S����%��5�q��������ܔ�W^�.�e�& U�M�H��N���+�a㽟�:ax5,ҮH��7�J���]��l�t�$��y�.#�W�``�O�=8C� ����"�p�`�#��ḧi t��_��O������hQ_O�췡'�媁�<xрCk�ª�wo+%0�9��#��ܴ�*��v���jb�����Ǌ��D�z(�68Y�od/�g�g�Ek��!��I5�֩�Ź�c���:4A�㲩&���hL�(��&��]+�5K'�Fa�Y�
B��Y�.U�H�x�h �e�j�W4���B�>f���U|���H�	�|�Q��Ô���D��E�5<��G��p~��h|:�D�i� j\F��:D��)����;P8�v><�6���$�"2�����l��H�� ���[6/z5�h������ [�$�!�]�<C���������q�A�O�^�sh��<�������0�~a�(�v+�n��]C(т�;��mQmo��:�]G_z ��K����7~F�@r��ze�8�	ADY���^�2Ej��j?��#��n�e��$�g�e��F�n�4�a�6����P։:(�F�|DB�"�.-2k!HPJ�
R���z^ɀ�<��
����P�u���6l���^S\�%,2�X����p�+uj6��a���Fk�J�qu왦	4��\#�iNjU�q��/u$o3&���K�����(Lv�� �zX�۾���N��� �#�=�tH��H��ƞ��|6ƒ!����X=թ睷v4�V�H:�3�Ըh~�'�KV$H����\�|�"�`אҍ���ǒc�R��V�eO�ҔZ64��K�n��!�(�^�Yc.�8x�z�Kqu{,�]gudu�/u����e�Ӄ�$��C�IR�]@�c�I�(�ƴW�2���qr�	��D�Ppg��@k�L��v|�����v�kk3����7��o�#ƶ:=jVBA1�pZ~lz�&��B��%E79��Ů��)��2�^ugw�B�������x��r��]tb��⪪�^9�	��7���䠲@^�.Je�z*��m'��A[wk�P��ۄ�d�������k
㏟�����hPe)��+jE����
���ʒ"�M�0�';�X �f_�!�����������¥!]�L��m�*?�a@~=���0��Z���+v���mǙ�Krء�$� ����mW��3�@a�M�!<2��EU��E����
�z�E����*��)���_F�oE��c'�s�D=�i^B�䰹}�䠛aYI/�f�Q���r�~�EnB:ٺWv� C�+��}���%"���c���j�-���ܟ�2�J�Q�?������f�S@\�1#N�ٛ��Jb���/�QK�)<�������$���N�3�=���ۣg�2�gW�]	��HnVF�sJx�21��C����b�|m�Ѓ�O�٬L�%��L���j ����_:���{M�x%{�xNQ�__|�	�[�u����E������x�Y��ҷz`iVc�ȅn�?��i�4A}�Us
���zK�ojP�j�)��-�r���iqI��Avɽ+���d�(%�����.ʛA䧶͎$P����?��m���m���Ƞ�^�?�.)������[����Ȼ�x�cM�Y�*WA-=�B�7aW>��J��K��p -R���j�/nZ"�YpD���]�H>/�S{����Q���9q*�����.t�1)1$�6��E ��a���G��B�do�!^J{�H�>�4�L4�ޜ��2HX;G�-oh��s�V���������m�>,�aH�w�`���I�ݿha�.�2�5�����{	�U�v���O��b[�9J�3���C������>E��lZ'�:A���x�=��q�^R�u�0����AR5��춀}�-�p Dո���R�;���˄+�L������~�v���2�����NX�L8y~^�;zrߑOMw�81)pa��+L��툨��m[��� ��8UY"P���VKE�`{��.��Q���\W7�=5{qb���1Zb V������oC?����àCx�Y�?���T���0ߜ�1h���GU2�<��B��k��]0�gй����7s�t��,�<��hF(��'!�NЇ�"ӆ�	��7�$���vE�S8L���a߲x.��÷н6�?r���z�s"�S����RC�'���À�:{]{�krt�P
F�@���YN�-+Z�Q�ںv!���B�/!��tg(|o�w��;�Eor٘��IgF��0U�|۸!%C������x�����8z>��%s� ��U��J��Qq��P�<�~�
'�nZ�c��
<�s�������A\���e=IY�?�W>9©!��NdN�s�	5|�Htj�C�))7؟�T��@M�8����n����GCN%qk5��~��vlo��$e0�߅�~�\��2��{�Y�`��h�-�l�<g��j�3������$\*K:l�3t�G.N�3�¾4 \
�����'�i��7[��+^�Ɋ�[qwc��r"ط�1S'�6���p���G�>�-O9?x��B��m�jwӄ@��fRr�8�r�I�1�jd�l+v&���b�E[���ʟXF�xk��F���`}��r%���uGh�X|/���ӕ��=�F-��xW��I����Ȓ������h���� toj>�o?�
 \u)��W�]���ޱA�^hz2���9�!��)vo�v(9Z��gF�#�-�����0a�#��v^��?�aVd��1bt��>��[M�P�V@J�.����)��8�UB��I���d?�������'8f!�4ǆ�����cB��.��.�b�sumc"����sh{a����Zl��J�X�fs�f��
N q�<}���<]�j\bT�_��7_i�-���ToŸ�9<Ft�������A��Xu�ϛ��Ϳz�����M��{K��C���(��&)�:�iZ�N�r��n����������q薪��)<�8��:�:U����P�-dq����wJvC��o?'Βr��)����I�`�߮�gxԄ ���Y�n���0�)r�D�и���Ƥ�;S#hM����H�VZ���3��r����|�KoI@���5dn�z�Ⱥ��fڱ�d��f��Y1s�[��� |�5�zv9R�K@�ÈmR�<���
��|��c���9���9����5�)u����Ve�#�S��ոa/@E��9T�r("M�;��K�w^����{j�vqۂ�Z�Jy{ ��ų���ٝ�ŝ��fݖ6*��}MH��/���q�� 1j�Oœ�Uu��{XPX%�4v�QƯO�k+��}�Vb�&�HN�c�M�}]�}՛�D
�t�V��%EN�U�OQ�I3�wr����`���Sd�SO�j9�sg!*�(�8R�K~���I�D��N�uK���D�>Y���l/Oo�6���B��L�Clqר:׆N.E��,����-���^m�Q� nظ!w&��q))Rw{#%��7�q��)fWݗ��nv/ذ%����,��hh{��<�x4�Z�ΘČ�@�R&�#Q(�~�-�����,��o��<���_^��:�L��Lc�lo1/��;Cx�w~4�G�q��I�̢E�zT�o��z1o�T����+�(4p�`l�p</��/3�v�V����S�z�vi����I7s�M���[��a�Г�����Xu�#}����D����2'[��e��q����vi�S�����z@�=@��Q ;(m>V���3�"�"|�}��e��������x�MJp��5��u��yx`\��{�C;���3��'�uN���\=�S�)i\��ց�*^S��D�q�sv����)��e{�@������m�S�:�Eq���$c�r-A\��t�_xE�[.ϊ=O��w'X���p�0mB�Т�q�P�:��>�I��WI��q�rE|)Yô�.�
�ϛ��Yv	l	�Y~�G�S΃��W�ӧah�l��W�_x>��TZ���9�uд",.k7<'�lxhj��%|�����UJ���6����J1�mU�bׇ�h�����Ȉ&G��ڜ@���t�%�����&$kA����@����Py[fՓ@ �G7\ o��MBi�DΞuE��i���X�#�����_�!8?K��K ��@��W�j�`S+bp�jo\��.#�r:�����9J2���ܼ��7�\iO"�������/n�)$w�F�	[	��i4>2�U����m�K�d��w�n��F�Џ�:!�������VOm ���;?d��u:+kL�Ƙ���02�U��̡k��W���&O�9�:	�|��h�xm��9>sG{���oC� ��g��]�jz�N������wqv�X����?�tLٟJ�'3k��R���*>�bh�m�D�t�D(�=幞��s����m�[�V���.A ��VKN�7'�ؤ�s�I2V��Jȶ�B�/��)�_C߳��▖-�~q������i��Sr"������u�ANS�56����x���:<͵i��4r��(F�b�M���7;�3��ço`��
MyG����B�nz�ZUI�MV/T�װ�oڇ�N�����y<]�d,��ڨ164��BBw�V'�|Q�%��h�H�z�%��c��П���t���Q�j��Oq#w�r���ͫN/݄e9pĩ�_us����`5ɉo2�� X���>hGHK#Шϩ��>Z��������٩liHت������¤�
�>����O�?--��|R"�M�,�+І_�Y~(lx3����R�8]vq����VO�5|x�BwoGػH��.?	H�����;�1�
'�d��\��ȝ��-�T���
�&+���A�qt�,���wm��ʿ'�'����۽B�� c<����6$��qnE=�e�)-Ӵ2����f{����]��zqz�Q-��]p��D�9���S�}���f>����IO݊���Gh��.�7�����(E")ևJ;Ϛ��6����7,H��}a9u>�� �*��l�1��}��������Bߺ���wD%��_�G�g�� �c�R��@Y!F&
I[8�����tcBO��y�i/x�6���|��4�Zf�#���>	�RD_7#N-J	��e��Y�$E��¡�z�89�}�v�#�лTjq�����w�.eHaF�L ��%���1yrG%�O�.GS�U[EZk�Sﬄp�x� ��H���>Òǻ�8h���oY�ꉤq8��7����G�h�z�P�>H �����^ZesY�-w��}�	1T��u�G.��ܢf�`ύ�;Z��Z�c���a��!!�m��S;��~(o���c~�+-�+�$҈ti��Y���1�?bS>�����ȹ��4�r�����ZC��^�T�gV�wRXf���9�`�A_�mBV�Aͣ�Y\C6�z� M$�]�}��4!�?K�Y��4aGP����< VM�C(�f���\kJ����Z�?؁��]�_:��/�(]/#͊o��r�,�޽�VU�4� BMʌ������v�j�`�Bei0�;15��#4ԆHr@�EN]K�
6ۚ&x����m�4�ĉh���lp8�8O�q��tO�"��SȞ�l�i�(�67�-L�R2���d�?�f ��%a̗8G��i�s-�tiS���󣿶Bd��L�˥��ׄgd���Y�9��Ol9��-�������-��ߎh^�7�=	���$���D�a���@Q�X?d�Bz�'�67�U,�~�3����V��x�!�X�rD���ݥy=�BI%~qÕ.Z��V��N�p��T�KL%�����[Vgz4�5	�n��/��d6CB����Ϡh.��i��A������p�C	|4��N%S"�o�&)18�!�-��a����� �3j�B�u��
��w��'�n��*�aሁz�e5I��n�_��T��ou����� ��4�����O��b"Q���Aj����h$t2t�w�.T��c4H{3�<~�/+�����i�ψKA�>a�#�������H`LJ�I6S汦�:���ܪ:�����&I��'y��:����rC��c=�_W����V��8.�3�Ӯ2,Z����͔9R""���r%����Sg4ʟ�gV2��uQ�����V�b��KcN����ҬZ�9'Awg{p�y#<���T�=O��.Su3C�.�VUt�����[�[���!!��k�f�����7�./57�Qhj��w��4��.}��
h�㬫��giϝq������s#G��|�n���0L�% ���ϼ:�%��(dj�����5X-��VXsf�D��x�_hQ�Fr7`]���%LL�79��݇�Q��S�/��0r]��pg`�iJ�$�>�T��?������hS�����iڑc̿��<��5!>�����,��k�d/}�q	�y�2UW����	�Aܺ���������1��!��jm�څ��XC�bQ"EJ%��<f2�@��S��U�HX�.��G����(�=?�#|��s��p�Blvw��&����2�XB�W���]~����c���U30��l�I�u�q5���^nyD	��g��郄SE}�6�0Ӣ�S9\�� RN
�X"6�>�+�-�ֶ�)V����h�]Wg�tN��,5��`�����  ^܂9w�dp52��w��!C�P���+���q�Ki���D���/�>��1#�h��,�)�q���|[�,����Mi{Y4�"�K�ܭ���ї���u0��;�����5��$�=�����M])׹ FMgLk���e�Eb�0�|��}��(7����P�8�5�P���K�4�Jk&T��~.4�U}���&�)�|����db��mzki{�BA8����h�T��$̟��+~�ũa���	2���������8/A��|�Dv��4y�GZg�h��{D�Q��)��WH`Sg\�WiZCD~������5&,zW�#���_?M�8f[S�iԳr�>p+��u|��E��S٩w�m�>��C߿�;�Ñ?ڡ�;��!W��,�H���PTG���O��P����ҷR3�p����JW�2t5l�V�|�?$)�Pp�`I����� �]G���b��F(!:��j�i�f=�TLlMR�t��!�Wi��p�=ݬ�f�1��^�0�N i"�U�;�h��̲ȟ�s���}�f�1Ց�������0#��F@��������Z;W&n�qM�;M4��&e<�$k6�0C�ё��S5��N�W��4 h��LB�[�)*c��ByY}N�c�':��C,bä{Q���*r8R:��۬��z�7zx+Aɫ��;�B���1[�$�L�$kQ�R��g4u���h/{�����j��aTo��(��[����z��F<��U���^:6"0(��L�`�~�"���m:|�bq�PPG`�797������qր2�=�9>5� �@�gF'�'�X3�`n<��c���+/�۵���>���^*�����9�h��������ef3����t}�Duy�S�6%nX�V��P��`����>�G��o[�S��B�^b沊�%�HJZg /�Ϩi����^��j���Xi9 KL��h��?�R(���d�#�������o+�}y|����L{b����@R�l�ѡ;��#��:���x "�ـ��Y���)�7�]��rb����[�5�������j$
WY:�,_��x��xG���A�(���y~}�uRU�F+\�z���G����_��ko9���Nh9;�]���ã|^濯\*�)_-�d&�ê{�"�<o87
��gF�g���f��q�y ��q�o��՗V��D٫�:F��O������<��H�e3h�QAy�S褪ɰ�l֭��E���������5����7 �^��L�&r;H�s��ƞ��:AΙ���i�����U����`��s��
Z� 1�&hѩ"��V�ǈz)��:��q��)v(��!�y��N��ҳh�\�,�K��bO�A�K�'�Hu���Ě�zj��[�jU��fI�t7��UI�	6�r��ݺ���IU�P��W
Z�GJ�� ��	A@��O͚D�'Uк}0陌Z�Kt�������ޑ��=GĀ3j��}Rb_�sR����H�D9�� hMD7���h�c����,7v�0f��i�'�um��z$�oDO 5��uv1��DO�0���n���5�b)qhk��.���!+3����z,{އ:�|�����^�"������NQ-3D�����s��pۭ	�4NAv��s���m��o����>G�����.�}V���و�̔�Ph���hv��j���wI�����=��u�[�.��a����1��:�>�K�s�-��P�2'�3mh����I�T�n
4iU���1tfbٌ�8 7)�+���;w*)h���n�9U@!|d��<��|�� [��!������JP�'eT��[b��r���0���+fа�	K�{V@!�:zP5nG�E'��3G/����1Ž @!�~�k)���W$c�Mx�e[.�v���ia3�{V� �~�7pA��w��PM���Ȓ[�J�%�L�Ĉ4ء��2�5jG��V�����u���Ի�)sQ�8�R���JqYlnUp�l�qbge9����+��$�Z$G�r�՞$`~�yT��Ip�� M<���%�ԃ���I��ߴ�'��mE��h)A-I��2g�66T��T��u'�S�NP�?��˥���g�yů��>�n�W��0��0��AIQ�ғ���u���%����	�U����\�Zz��-�?�΅;Z4�;5�R,��y�!٠ώ�'�PғΗDgB���*��R�O��E-����&i-$D�[��Z��}~�ģɫ��X���v������=�͠�,��[D�oxpV;��۷���r̝�J�0-%�4�݀��������)[�@�9�l���Ѿ�n��'~�B�Vldϫf9�@^�8��*<{��S:�o
����RHe��.�pV��x]"'S��.��^��;u4�,�/���έ;聰���S'�h����Hp���]8k�Y�����S�c~�z'ы<]��K
�kG�*�7�Q��2����QrH������\S��N�s���bsZ���gVW�[dw��c��2��5qKxB\O�[�<I��投yQ��&��ކh����R�ShF@н�m%Z*i�F����{�-��"�K��3���<%0�1a�˕Q�\���/�bD�*�&'����@Q�!�U�냠n��fDdR�'��z��#G �/���?.J}w*�h��W��Ms�!8����(��A�NK�J�1ߤ`^Ed����Y�\�16���	��T�Ԡ�F8�������_m���	������&�)���s�J��S>��]	��+�m���$�J���0�6A����$���¤IO�t R�"y�'� ҅���G���H�����ԲY�����-+3�7�����8*DNW�j_zMl����Xn�������]�,G�xȅ%�`*�՛�HX��tAj�QO��H
7vbgFD#�p$�:x~=_�_e��5�$<*x笈0�u�7��l��� F+�5�"�*��0�D���3
fG c��_A�r�,	��O�KT5]+�Q&����L�ۻ:qhܩ�l�����SM�ǡ��"z�4�NR��\�*���P��u��X+X��oo���͈������Uŗ�r�����3�/��B��0�(B̺P���8}eBm���r�8�2|��sT]�	��sˏY�N�σw��iȘ��x��i2�t�GQ������'���>JN2�h�6��r؍�{[?ѱ�:j���*�V��K	������>�c��������Za)#���J��C ���%��/�6j*[>]L\5}�O��0eMO��ܨ��J&0<���d~�9�q�F��q��R~��W�5B�A!�d���<�8߽��_`F�)cZo�k��"���!TY���%�[oy�v��}?���b�$20�!���>����1q�]~�����x��!VN=8�6�B�$uGfԑ��Љ҇v��K��V�g��V�g猐\G7iӤRmɧ,:�3�Z&Ԟ[1����n.UK^��WC�"&��N��1<H���9@`Z�^��Cр!3���:@����!�Xv�ք�h�w�����R��z>"�G�*�a�mW��r1�ĭ�k~�.�q��h����[m�梳�9�[񹫃����g�q�&�B-�@����Gͺ�6��D���j*%�F�?-;"����=i��<B_�q����F�i�u#(�!g�+�jF��{i�)�X�!wT2_��e�Y�M��\[�6%	�XiS������뜧������C5�a�K8�p��������5P��$o"K����^;ӹ����̆�/�Y��zJ������-��9 eI�z1_tIf�s����K��y��h[̩h�@�w���ۉ �e��
ݣ�.L�?c�I�q�h�gIcV���U&6DY~M��x����Q3�
�Sk�	N0�;�x�˃���ro�U�L!�떳a��7�jTf�I�
�sj��iv�i��1�5,��Xw��|��p��x�AR���x0���)$H�㋦�c�}�	t"� ��C��: �`Ԍl!�P�m��LdG���2����v(�zk)Mjǀw>/��%�{����w����z�[qYM� >� �ͅ9<�}�O�>��@���l��:/��w����s'�����S��"h��+�v��#�p���,�]��G�J�V�񀬞7(L@��1��n���6%����s��u����Kҽ�F���-������ʫ9l��-����)�6�0�܊]��,��W�j�{,HQ�l�r�F��at �דg����k����Ƶ��j�1/�K��dO<決���)�Q��ml��t�i�|\)\�#*ତ�I��km=��4(�?�IhD[��!@�3v�&�m4d]$�aU �	*�gn{]:E�X��3�x!�[;]g�H4�dpI�эx������c��a��{P�@zk˺�Th]��9U�hA�c�a�����A��������'�L�Bm#-�O��'�ĕ.�*�HW:����L������\��ڷ;�Bt�����g�R�c�p�VUξ����&�+�P�)�Z5��<u+�C\��'����fه���0/����^O��ۻ�쫐М{���o�Ĺ�U:}š����}�vH�=�]�ú�@���zQX������Dl��ͷ�X���y��N\�"%��������Ւ�Q��(#����C.ߔhy��F�{��Y\�]�d�B��۵��b� �|��vd޻]mh"�D~�Qe���i�f�Y�V{a+�&XA�y1fl�$�A�/q1򧵌c 8酫�#nl���g��L�I�g�N��~/�v�o�1բ�.��L�,�j0�A�_��t���=tD��Y��k���I�Af�n��{��jzrf��\眆?��{IQ�f���f�v�`j�fR��ă^*����ZѺ/�0�&��A��o1���ZP3�9�+���W�=�`:��UT{�>~۴�LF1��7����'�-� �GP�NF2�)<3G��4+#��79P�Y�7�����?�?���L�(�D
r0Ϣ|��&!q����d����@~Cn�#�e�� �.�� ���zW8�5��j"�J9��X0T����@�T$ق�� �𳔠���̗b���Һ�\L"����-E�/d�a����j��+*��=�,���r�ܶ<Vʢ]�7J�A��̦�;�R�(�H�G��t�],��޾��s��A�{�ԁl܌|�Nٗ雠' UD6�~)�K�K��w���G�]d����`�KC�,��C�]�Bꤋ����)���WxZ�qXؕ!x�.8����*�y(��_�}r˔�<�{�o��m����a��Y�.uE*�'��ngJ��I;4���Ȍ�@�iw>�Z�Aس�I�o3�%۽��I��&��W�Wi�~��I�f�#�F{�>�����ŊΝʦ�����o�l��+������pS{>iT�v�~ ����3H�}��lF�U�ˀ�R�,��\�g�8��^*����VV"��Т�ʬA3p�y�fH£?jǲ�A�r��ڏ�����ψ���ل�F� �� &��o�=��C��m�8cK��brf 7JS�4���tKB��=�7�N�c企pOb/ώՆ�	n�@̇�.eq��>�h���Rd��-s����^A2bYM���.�	�l�Xv�h��}5}Da`ަlT��3�Kq��EL 2��1T��J_��ᒭD��L��X&J2f
�3;�����Q����(	c�w��yRQ�e��KX}�uV��
��݈��k>�X�l�kI(����wQ��BFRBN_���0O��G����t�~"ͅ=/B%i�~�u����������̗�]>��|Ns�l#�Z�e�'�� 9���c��j���$�b�蛟Hm=�`\~Ua�p��8�ˇڀ5��8��w����GN4!����Ff�KiL9 2g�����!���2�ONn�yW�ȫ�5D7)hn1�\�hy�n��vtS�VzG�L�N���.���#C��������/���� ��CY�~�k�>>k�N8Y����]���B������Ƿ/�w/���9��.u-!{3dz���TO�K�8@��F7��%X,������^�#[����n:�_q�ҕ����!!�C�|�H潇���d�m�������P�AOod�������Y����Y�w$�28j2F�"Z/	ȱ�jC�IL�,���eq��tR:?���{@��	&�G��� $�ˀ����;������,��@q0�<+>���Ǡv�V��C��-?߸8Eo�x� as�/!��4.�e�\b|�rͪ�ҕ�����9����z�lx�	�it_bEqb��"�Ux�1v�pu�՗F�r��ٹH��UOHHɢ�(�E��Ϗo��RA>��P3�As����Z&��n4���c�,�ҝ\}��ZN�����lrB���гc�[d���K�D�.o�ǵ|�D�9��S �؂2!)�o�A�#���{�3����w�� 	��e�x����
�	c���+����A"z�Q�ɪu]��>�4]�l(�z	���ϡ#��F����Y����Sə�$�)������k��-��@	ӊ�#�ʤ��LT�jF�`%���Zu��sp� ����:���!��V*yt��ޒ�-�GM[]�	�ĩp��#�=��W��M+������Z'�`oK��vWp��]��(Ac�������^��rؿΚ�I��
q��}�P@�E��;��'�ϫ���Wh���7ӓ^��dW3-Qjk�����SwW�{P��q�T��H�\��٪4Ǟ��R����Seひ?���?�x��7�7x��BBzC��$���IB�C�Zof�i7��jJ�<�V�M�����:@=*wG[��nTK�����Ga&f��"�x����﷡��7�p;C�\j�{�d<��C�'TT���>gٚ�@�
�u��A^������|�g5���0H���"�[YofWO �G�Jwf�ϵq�q�Qx�L���ճ��J�q��x8M��N�z��^��$��ǃA�"�W_�<尜�W�)���<�Ն� ��%��ߔ>�T��c���{7��~�L�R�n��Tg�k<F��7Vyx@�,���zt&y�;~b�]�X;�F����5f�|�SG��uM'23�9�T�/!ZQ�.�SC��| ���Uح�\�K��Ҋ3a���*���{&n�p�C$x_�������I�rk�j����ϰ���-�Kd�y+�'ɺ�����\�<�<� �qE�S�EVZ��Z��S�y���!�#�κöA�!"FT6�^4m�|���L�� h.�u��~�Դ��i���ßcf=	.(.^�r�6��-���֏nSzt�ؤ�u��W��6ji�/�s�5
�;>��Q{z���L�s<��� �����1�e�K�y�dB���(jBLXzK�#�S5��6ˉ{`?U�;dBX��x���^7K~�9	I��,�`�W��
�:%̈́_v��[����2��,�k���,��j��<��� 0;N6TvT]�����s���J�X4=�H�''��L�9�컚�����X��,I%׽�_��vl�%zJm�R �ޗ���U��K�����<���4G��g���	�Q;*�����(�! ��~�=��F��(4�qk��1 #@�X�,EK�yM6$X&���]�j˄f��]fV2����R�A7���^s5���ؗk���K}#Nի���F��NU���&��^� 
W�k^���������>6�!m�kO�`{\���w��`���yD�������b�ٙo����s����ƍ�����x�]���N&w�V-�S:;\_��Ab�A|�p�Q[��Z��E	
Ʋ�`���9�}*������o�\��@?�To�m�����3#2!W�iO덿a{�l$��ۖ�=8�k��/h�N�ϲ��aǱ�P�˕�dR�ܚ��*�_����~K�܁�����+�6δT��b�����EN�j��e8�>�^����P��F�\2��g�W�=d��l˴�M��u�!߰'���###��cZ��R�@⍔��_�/s���Db�B�a ��;4�X:����<F�� �h3�&��|>���1e��Ώ0~�����߱H�ݮ�)0���k=����(�w��I�iq�A��z5�mw:������=�n��b��I�*��b�A��C�b/�����q�F䮆I��v����Cc>~��;5}V^����!���!ӳ۰9�g��9�%� �Q��������u̅�[v"?h��?z!��lVս��|v
�b]ʇ�ޯ�5d���r'g�\��?����P�tű?/oq�'�LhX� ƕ0v�d.�B���+��2��@�-��L�l�eq��w����	9 /�/���},�-��x����A;�N�����ޯ�pϮi�����5���lc���9���	�w=�k~3t|���&�=�|�Y�CKk�
~�r_̻6S�^�s�^�6ע�v��3����&&Bv�&)�l}s��5v���ۋ�T�6�ٸ��Dw_�Y|�n_&L8��|�@�Gʖ�m�����N���z�>����R��x���Z!��@����
�
S�=�P�蕍R6V�+J�9�F�T�)OBS|��\�of2��a8�G��)?�'�Ukuu��/���Fˣ�On�+��=cV�tY�rs��]��I#	�nͷҷ�XT d��Oi|����.�(�If�9L���*��p��ʑ>�ls��Y���A���;�ow:f����&~|ޣ�_E�0fzB�Q�!P��j���q����Mh2�F5*����cx��S�k��¶�����������8;��ҫ�,�N�pg���V��W����,#"e�'��2Ot�6�t%Лh�\s��p\��0���Uë��Z���>��������Y�4��2&�$���`D4pۣV��Vؼ�����W��"7@�u�Q�<+�!�/�[D�@����2L��RGn�>n�2?m���4�g�,��"�mޫw�E����NŖ��X�N��%�Ǿ�R}��ԍM���_��*��h}�n��)p��W�U�<Ͱ&g����I��)!S���e4{��<^.1��G����
�M�1��Q�:��w��|��O�U g���S�A�c��?&�_e
m�>>O��� �z���ۉ5�C٘\��J9����L{��Ε�r��{��i��fkϿ�+τS��"�����G���$�F��lSEڿH�Ua�.�
�o�L����V��>�ΤY��[t3&d!�o��M)2؂\�1?����}'��z�%�ttҏ���g��jq\Ţh^W���M��n�Ie�rx�g�-ѥ_�I��b�?�@����^��~��CFť��|q��Ǆ$!�w�)�$!v��Ȣ;G��B�3�S vKC��Ȫ.�}�4����Y��jM�q#6kIjf�	B��L�WL�Z�Ql]��Dȱz�^Ì�����M�J���ڰ��%.���g�GN���������Qu��;�����OY|+�������!A�W���+\L�B���:Cq�g���mγ�"�=�Ȼэ:5eG�M�O��P�ߙ�����1���u�W �%W�b9��_���^�듺��WTĻ��}�yR�S��.��H�:'#�\�<`׌�R�u�
.|��k�}R,͓@_m����+���Dxt7kXi��[��94�#؍�L�N�&;"Y�f��c/B�b���"@�xK�	\�*���f-�W�d��G����>�C�(s�B6��߬K�]��>5��6��N{7htԩ��:q�G/��J�����|��Bbء��@ُ��͉m����D8���>�&nREVC;a6z�r���XD�۪�s��[8rR���M6bb/����-��t��O 7,��µ��à�����lѾ����X*�x��/�H]kɸ{�1�{h#�i��k�����s)sk��D]�� o,	���!�{��p���~�´��8�d�9v�?(�"�<1���\L�?�Oe	�ڏ�0%b���w��ҹ��{F�q�w�C���p�d{���υ�������A���yߠ�A0��a��H�֒�\#7Z��͗����AhH%���A��_p�A:�J�,��p˝����?k�n. '4��p��L��yT�����;m7��r0쎭���y�����Q->��q�{%�M����c{��d5H��49'�nX�����s�d9�r�߶��v��Ӳ�~gP9`S���m���]����R�ڀOAǃM�{8��
7�����h+~Ұ�@�����L�{�l$l[�"k*ڠ}#p�֜F{�b�R�l��)�O��n�~��̍N�?(hnn��>bJQ���i�`T`b��죚��f���;�ç���%Qm��"��X���'Ö���� �,���ݟ�PP�68��ˠ����5��\�_9�z2L�گV��v�3���/�	��#�ܤ ���gTW��ۊ�W�mX ��A���u���ٺ�1wMS�j��{_)Y�`�<��6TK�����y�ߟ�����G����	�D�7����d�g���veouL2r�[�w��pD1��Q�t�x[��<��ECja�<�3/��*�M�?��ƇC���dd���S��e�p�i��cuY�jt�-�$��n}΋Bg�#Y@7V.���Xt�ߋ?Pm� +���������;y�{Bof8ΰ�!�J1�F7lx1��~�d�s"�f��Je�yx��^����9r�����m�U]��i�NO��qu��=i�4Ж\�m�����{m�^k��@�9�a�0����2.�۱�2��4FS4��F�ci�7`S�0����uGG��'�� �R�'�cȮ�fa���n��֐�l=�� =�%��oG"�0d�h��-j�{��k��X�,��WB�F/��v�v}\
O��Is���Խ�dZQ]y|0�|n7c1�����Ĭ�b���Dc�B�A��D��s���ˤlP�_�A:�a�1[0�j���b��<̲T/2 ��b�Z.Wų�Zb[�uvG�l�nźa�����u�t�"X��H1޹�0��T)���	�bp׎#N��Y��y����q��I]���_K)��C#���S�gzmQ���*���"N��ikyݺ8`ɺV�3�nV�3��lѡ��'�6R�ll\M�m�ҭ���=9�I�?�y�$u�_6�!��z�S̕k����x�9ٖ�0w��B|�ѐ
��EL�T�5FO�^'A�������Qȥc;%��
�Yh���H�5��<_w�3��_B��,��2�KGP��O�Y�։�6�mI���@+�,�:��óF05{6��c�N�=�@ra,k��c�hQ�X��恕!o3��F7z��K�-�t0�nް��t���[�^X���g�@�Z�-2}�s��f��ۘ6��ƥ�΃� EJ� �yw��F��_+���\M��ut~#Z+��'/k�bH[������Z��'z8H�����^�����O}��we��B�i����N(���,�����p\5�!��_}�.�/���ܶԦy�/��템n���r�x���*韲�������)I�]�0ˈ�b�,<����կ%o;��ůXb.�LM����X�Ӱ���=��-�y?2�U|s�3�i�~�=�.�� .U-��h��ii��̇��!�B�\����/vfh�,=�~��)�{7�hy���5�U�
�u6�]w��y���gY(�@�sƴ�j��O��82��j.���X~JtTm9�kg��u{�Pi�r4.���<�I׏����� n���R����lG"��Q�x��6�o�v�	+��Q_y�޳-Q6\�P��a"ْ�d:�m��͛����/Q�H\�l`%԰ug��o�!J�������Q�Gf�����ݬ��mK�@���r���!�{ѓ=yӰb'; 0p����:{=ka�~Ͽ�Qr`!}����J�4�)�T��;ø���s�i�D$�ai�Y,Ra�v)������I�1$���/�!�C�#	O-�3u��w1�������\�D+�.�F���N�1]}����̈́zi�Q��7�R�l��P)������ρUJ*�Tgp�K�v�{�M��f!���}�,w�g��KEI��{����y�Ʒ��'� oeZ v�׆n��u��ъ"K7Q-0���r�f!��N�AQT��I�Es%fF�D��@�_�F��?3z�����������R��9vJ� �$���o٣�õ|������)��N�8I��H��j�h��[8cv|�Ѥg&�y	���>�@��4��x4l����q�(T�ቕ���kıvT�o��!��ڞ F���YO*`n���`T[�K	���H`_��Ѯ��L���&�^͟�[����l�N�݋��cgr���!�Y������2 �a��������w�X�ӊ͖���[�$���}�/�^@���U$,�Kۈ������Vc��z0?WWN3�x���j�^e��l5u�b
����M��J4Ɠ�aG��ɧ������oIه��7�c�]�?Č6����������@�b������Ѫ��� ^��Q�5���G�٬��33B]�Po��D�B����$e��U8���i'ݓ�7���r�����np��s+Ll���_@�7)cV̏<yFP��~FL^vJ��H���q�%,��c$]��L�4�����0
qf5]���'���gB>���р���s6'����������]��a��Qi�!�Gn5?��L��r��^cV���[R��Z[%#
�Ӣ9Ԃ��η�ʛ�ޤ�u)%D���E�t�M��|�miƎ�:lbC�Vg��p��z] A��P�D�+�OG�{,�1B��n*zb�ߤ����q���k�=Y�I;�oC]"�A߼4�p@(�{1l���/,c�����
�[�qTfH���r~�5C�rQZ5k#�C5���`̉:B�[����#������s��߹@���:5�)[�Z:�ĝċ�<ډ�cU�k�i��kK�[qqDHz��.�X]�ޝ�)��~i,i��i��r������?�1Lq7`����O{������ݞ�ʥNIlU�wgÌC�ɹz��ֶ�}J8��_���>zSv�W����2��_W�7�o7��t��^�;ؐ�"Td�e�{lIp�l�kq�[�b�������b�{��-x�[�O�ɱ�ցeJ���ی�籩�?R\M3S.HKo�6�lF"�����%�k�� ���D�uٲ��h���f'4�UGd�8�E�Ť	{��_�oӿS(��S�kY5\���/5��,w��+�87ZPE�=��´����p\~�u�ݿg��lv�E��P�� ��JH��|��%�OɩE\=pvP���f�������Cw�:5n��P�f��mH*����ut8� �*���fm$�K����HZ`�J}r�hxf�a�*>�D�Ld)H�~�k9:��_��O�}�M��`*[���"��ġp�=2�!��fɃ�!���+����y���X�"8�	�$��k�Ϗ
�U)�3�I�A����&#o�t!�q�+$�FAأ��3O����S���X�H�S[�o\Q��xy�� Gt�]�J����> |�@��<Z��}(���~N��	�^���Ms���G�9|�D��?�:l&_	�,������yO�S��l�^������*[7Jg��]��hqc_�b�W�=����s�2x𦑘�ы�lt�`p�[�u�:L� s�;.�wc��Tt-Fp�5�BHu轻O C���%��Y���?y�7�n���F����}��m�.�.��|:��\+�˾�/��|Ɖ���Ù]��å�6]��3�Cé�M��L���k����Jf�ƾd�75ڽw��w�5,̵"�hMt�&ߔ<�A�n�*����&�=$��(��8.ڿb�B��?]�Ś$b(����I�#z.2�9�l����P|�=���
1"��'~��S̴�U���z��N0��("W=?�||���V$�J����̓�qn?1��mUa����N�V���>��f�מ�g����̜�W&4Ҁ�ۭ֩$��>C=�KzM���K����KR�y� �qrSf	���(��7���3�:Z`o@��k�]^��u{����ΓQ��4�B�ГՍ?��Ǳ=�D��d���|0-� 1�_�4�����w�� 7�pr�d-�E�����h2D���O����;������>9ӡ���r��Ly4��=Bw�V�������E�<3A�}F�&lh��c��Q\����������kT����r�{�#�=��Q���)BJH��3q.�U	W�R��uE_
�:��J�6r�nR��vQ�����oȍ�C��Ϧ�Eq"�P�:���T��3�B�	�&w�� )�K��n��-e���������h��`�DOڸ@Ģ"����Tz~���6'*�eM�!Bݒ	h����M
������h6m`��UF�{��̭^�����Z�(��
�A3j�*Ȟ.ƹ�0�¨"�ـ��������\���^���3��\��WBV���V���d�E�P�a��i�5H�h�N��a#Ƶh�C	Kc� ��FFC���l����7������
�Ю%�-���"���h���0�l:����!X��Y@�s��,fo����C�䕾�����$�IU&����h�L��d"��\�9��e�#aA9�ީ��W1B�T@g��Je�đ��B�C	ZP�E\�r(b+�!���Zl�������&�����~Ves���p��mq�×����nQ.Ld��%��{v��u@�є0�/E�@�;�^�'�ֳ|'Ki��[�*$���Pq݆�$-Jk#X��v�4����5<&D�FG©r�C`{<�Y�������1��v׍Z��M��Wj�*7�AC�E��r�;�������W�Y\te�P�g3�'��K��N����k�6"\�3�W+Fa�?���ޥ�irW������[��`FΩ^��ק�t�� 9C.Q�~	 �zh:��sw<�;�ɔ������]ۘ��gì~�݌� _������e�y�(bz�EǙ���*ǂ?	X�9H2�v`ǈ��PSOmJ���?�ņn�:LK6�	��0�X�p�E�v�ϡp+�S^5Rb�.�7�F��ˆ��՛�ĩ\rY�3T�t�l�ؠ�u����JV�z�]�����W���^�ӗ ����5�/�簢�qKka�[$q�ڎ�9��KOx�H��3�У	7�p#���ς �vs
��ze 4��M��Y�H�@̂�P��,�n�7B��c�q�|���E\s �4�4���f~�4z~>x�[�~ �d���7s���!��=�}�8uX/ٻ�̳G�7��g*��݈f�����g�*	�}cVP��I�L{�t�r�e�qlw#�$����|�Gk.1=;����9�lL��tBx�:�l
��0�*��2	1)$
ֳQ]�r��.#w��ȴ�6��ڞK��`��-#�^>�m|tG��zH{���] K��wqe=�ئ����r|��V�7���#y8 �U��2)2FaN��k���N0ō�|�È���Eo��|s����W�2��AL�#��s-��|_���ѐ�K `q�`6L�^�~����3�������B��dU�K��Hr�E\U���+��k�2
��s��d�8�b�1��ǝX��w&Q�0^%����%���i���M:6�8��qVi��
D�p��b{���U��(���d����qs�T�g����c����4��Q,:�O����v���&�o0+�@t��|�'S8<%a��a�j�Y0��v�e�M��0�+�JM%thľ+�*���6�kU�B�._��v�ᚢ����]��S�յ`����g |�����d+ ��vF��J�|� ��XIX���?J��S��i�̖8�?#c ��L!Yء{�i�x<���<"�K�*٥��z�E?P>�6�nر]����b0ά�K	�g�y��6��y�"_��f*#n4�7Y;�EI7� "��̃D�7�i��I}"��A�����+K0�ɶ�������2>��e��p��=�ւ� ���
�K��_9�
V��Q�&�qsQ�
�d�k�t\��p��K�RK���M[�PrAg6�m��CH1+n��<U�n��=��w�ܖ�����:�}:�=�<��F9�B���TD��u������!q�]bN�|�\�ì��׬��ᯖK\sˀO����F���״�
G��X�:���=�K�z$�hu�ǅ��O�+��F��H_�����ѐ7X���٦ύ��g�57��r��"!�E4�r���L����2��!��"1�����Oq���� 8�'jW�@L:;3�#�7D�����}��Yh$V�&;�!]Z<T�T�$��a����s�R��g5j?�T�K)����#^�
M�n��0G��-	���K�O����>�?@�BC��ȇ�_W,��xJ��j~J�F=�Z_Ӵ>��[yFh[*�gq˰Y��%]��h��KЏ�)Sh9���IR�r���wnP��C�$}����R��Ȭ��;w�:�RA�>�y��U�8�����¼=��h���W4?���Ż����� ��G���'tI���AP� �EM���'�ǳ�����8;Ogϝ�¢��=�z \8k2�QI:S�GsK=�a�0�Z��Ϡ��[^�MPJ��u
R]�H�+0�J9�xE�h��NG*�
��hղ�R�ܴ�W ���7
@�D�_�o�0��,^�|p���F����Oq��ա�G ����⌍��  .�聨r?��Ј�N�n3�pYö*ݞ���{��jc20��}*��9�̯j�*=�ln����j��_0��9t�|a�K��,�3;۩� �Ll��z�a�+����Q'ı�����-�t�Ƞ��B�WA�I�Ǆ��ӚAz�	��F@\ơ+�#"����T�7#DE.��d����7i]��bwxo�T��ڵȨ?y����[���S�2��o�TK�C5�A�s�y>P�mr��G��\��.-�H�e}�1X�r�OӇ�ǧ��ݟ��/�d��pqۦiZxo��?I�O�����oL���d�_}e8>�d4x�JT'��7��bl��֪�/�n�/	��U���a�ט� '@)$�2�K�R[�-RL��і�M�>/E�����ߴ�R�O'#7��N�I�
g���ƲRf]��W��[�Μ�F��Kq��cPA0 s:�	`F-�C�o�R�FvBa,m�[��
�O����ѹ����+�ޒt�T]�+Lq[kp���O�K�:$8���p�#D�Rt_p.9����ZP�����M�B5�)��H5�@}ٖ��<��@\P�+ڶ6�`VT[}Q��O�NG>��:�\��DRr%�U�g�)'�tu� Ci]�iz����Z��)n��ay���$��3ۧ¨�W���F؃��)(v���s�#'M�5�+J{x�V��|�۽�9x?IsI  &�qITL���{��Q%�eQ����YZ*l�E,�L\"]|,��a	�����A�z#�Gy��/���	6�����Z�A��.��"��a������sC�^@M�9���b�	�Ʉ#�	��B3�g�J\;��L"i��wܹ�Ƅ�p��K�]�����2�D �a�ETy��Nq��ı%0�g���k�qn���snS�Gpi���f���<�L��J��	'GԢ���Ch��%���Pq���d�Ϡ�y'�f�=�*�#�����cW�*�A��(���BH� ��5c��#���D2]zG�Z�y׬ϗ@E}�Έ�"<���X<P�-o;�i|w%-.��b#�WB+}��
�Ba�w)�YF�C4��A�������A�ĵ�߼�:[�"�����v�F$A�G���v����u+��j��I�-����fڼ�(<��d�Rz'P���Dޘ��/'�).>liŮ� 2�U`<mXMK(�U�_�R����F�ld)�f"�<U�&0($���������+9C��ZX��Z�.�	����2�(	1|G�
���Wpƽ���k�
_��bK�x b���am���ÿd{m{���7Щf'T��f?�MĽ2���+Y��&Y�ؓ �Zy��1+�e��>L�׭Z������	�F��f$C��)�/kԡ�1���qK^��������1戙[X����Y'�\00l�}�g	�q�8��d��-���o�ې	\��	١�t�ʱ�9e�ݷgK�ۇ�-$�h���*G�SJS���H:���"Km�g��zU� ��Z ��֋��U+�
&d�`��e�
QD�m���9;?�:j���"1�N�/b��#�~+�x(0SxC���n]�_�=�+��cA�蠮�������Y��P���T�l$����CE9s8�L�=j����z/�n����
k/���h��E�����OS^/ �=
u��Ǝ�D��s��5�im�K,�PB�~���y�SEHmM��3u����|eGi�S�3�XL^Pơ+t|�J1 O�:��~�K�ED��� ���}4F��:8�����ѼP��m���fG���'�q��ǘ^1.� T��ܬ�"�|�a7'���[" /��g�@��'%�K�%�d��e�>�̈́KP�����h��	�N� O>! ^Az}p�"�4�{`~�e�0�S��h����G(�R��qw��n�Z;����-3��C�B��ژ�yF~t)�R���Y�F��	��m�2L�͜�@_<6�=�c��Ps������϶R�< g �V6��d�S!߬֍�wF��Jl��>%��I���E�;�����D�K�h�*�%����Z(��2(�]�w��N.�	��Tp䎰	!;���p�xw��J!4E "��5���6/�[�=�o3�H �Vw��{`��#��E�s��~�zR�;�(���<��㡷�g��c���\��>���n��ꝿUBvRV?7y�{�T��-�p��8�*�S,��?����u�hw��{��ܺ����a3��~�ڏ��ܞj@aʸg�� �Ukh^��o�XB�*(���Vأ�� ����z�k���ko��ZʈC
���3�Z�Q�:�܀_���@ѫ�i����)�m#"`%�?ˏ�<������qEC�TW�,�m��g� #�n�'7�m�ƾ9Ɗ@��]	�b���_}�BV�$������<�%�{��{9Fv#�vXl��1Ķc��Ԣ'��u,���Sdw��\��#�Ϫ�Ö��ےQ`��ʁг3�j�)��Ĥc�?~��,s���Q3�?k��,4#AF�1Z7Ԍs%N�}��Af�A��Bw�݉�z0mv,RL���H3UO�]�����>Ѝ�y �6�h�	�B�&:�/y��0��$�a����9
��"��?��L<9q1��E�8�~k%��X�{w��!=���4���'Hq ��$��%#?�x�
ew� �A
�x���E%�ߘպ7A��ER��k���+pI���LU�b���Q�ءҲ�h>[~�'ĉ��������t�_O$��Ā"�p�l�;[DqY5h��{��$��J�K>���:3�H�L��}��a�ɐ����H�����ǔ�D}�mHq*Y�1���(�����o� aq�V���ߩ��;TH���}=R��%�W>�_c�Ѥ���M��&�:�Ę̄� ��q��5J���h�����ۖS:t�!!D�/In������=0���G�F��������S�Ի��ol���~s^��d<�&�F�H�V#��l8E�h��|/�g9��&�GG*E��k�����N�@F��I�z�3�1�z��P�m��F��t��Yy�������6����ڱwE
�� �;F�A�0bl�l��H���A�:��^����]Cv� �
*ot��P͋/�!����Lf����v*y�Dnы^��ϩs���oX�)a�}��rT�3~���Y0(���˛�k����6���cכ� 1�� *}�#��e�$Y�9+U����%�XuO]�~ub?�L �����/�nC����c�h {P��E5�*�^������11��n�8*����A0��ǌ�ARy�1��H�J5mS>h��ơ#:)Z�e7f��e�!_>
��
9�����T=`���V��mCk��;�W������*~ԅ:�Q�����`��%��_hZ8���&������QE�����axPu�\�$3k$�TW�s(��E'�?���1�mt�
�v�X�mo3}0D����^�V6�sʇ7&�;�P{k�FYF����*s�T�}�r��{d�Ńx�>�T�
.7<C�����	����I�'mၽ#�?d��f�4{�mTWw(ǩ���KFm��>K5R�R����C I�"\
s�z��ա��a��04 �n̻]*J�Ҷ�8y�!�My� ��%0�d�_�<�RJW$ f�|�H��5��|+J���	� W��Am�.�n2�Da����w��a������D\�v2.�� �&u�q���n���e"��-v�� �xb;�Z�.��2ʱ.+��L�)ۯ"6P�%���[����f푷��X9�ʌpR�{����@T/����.P����!kbo����xݍi�J�Kog��'@SHi�=S��Ƴ��3�+�w��(ɐ��h�����P ��Νf%����V��G�M���6�[:�le�d��'��������c�����}��5�	��G$u�Ɗpĭ	V�*��`��^H���@n���20����#�^�<�HE�U�!>4 g�(=,�kH���)����TW�w���7��6͙����Lj��!�P�2cPryu��n.}($h��%F�5&z�I��Al#.����:��6#u]�1(\���F�S�֟A������k�WK�-~j<K�k@�N����D|`���wF{�՘�r~	�I�y��ā�4�y��;�0�_���M��u6�FҦ:�WkC���w%���]q�au�:�mir�4���\Љ�H�	e\3߾P�n���Abf�'�?�8����?�q5^��(~���k��n��\^����ڬ6L�ݡwgCe*�+n�{;�J<��EW�v^��H���W."����&Q:W0�QY�E�@ӹBxeL�T���l���׶����k){�թ�֖/+�t������X3����� a{��(Tō����M6�+PlHPMCpz6���V1���
^�Qa���DF�/5S�Ek���1�y�%���cL��M�`V~��R��*�[��`"�ج��#G&USڑ8�2��$�!��������
�BPy����qf��yi=(PNq�����e^j߈�rִxg�N*=.#pu]�#;�U���-�S�S�?f���uK���2��S��B~}�_������vM�;h�
yV��	4[Vs��ܴC�Pj�
��'�9]LKeb�N+*�Gœ��ߔ�H�H:f[�L-u.
�-K�%�k����F��M������l3��w]`�L�}�a�]K�E�Ve��N�ʐн��d��>��~���Il�W�8�U9� -�� �N��o�s]�z� C���y=P���0G���r0k}9H�/Nd	^G��G{#��Th�c�UK+B�u��X�޾�s�DS���24[�Tr�}��Tr��'A�Ͻ��S�G$-���{�&���T�ȉz6H|�M\����;	HN��R��v@K�J��O��I���)�:_�����}��^��e�K��s�J쭯�i�+<�����W1A.Sҧ���8opM��k��7p��~zeU �����r�����tq��]b��<!Q�UP���C"�X�����G�0s�w��el�W?	C��i�'F%�;�.�_2���90���2MCj��aЌ%�X �i��>gg�|x��Ҥ�Ԏ�J�I��AG�s=��7(LAJC��0��YX��Ck0]Bڋ��uڮ��D��9�$%���	fP!#S�D�.�2��h63i`��������ؿ��?��"��NW�|�Qh�s�������^���<�)^Y�JtG��{,,��Ũ/���g��Ф���7F^�F0E0��#�k�rVO���#��� I����E��z3`J
��B�S�AFA�]��ڍ��&�!�xDs�Ɏ��.V�K�eh�"(��.r� r$qX�h��6��T�`w)O-��K�"�!BK!��+,�-ѭ3l{��n�����X�}���*5" �тxDN'��7�j������ͤ��<ةR�*
�B���g�t�,`�
�ߠ�
Ґ�}�G	��s:$�����8���x2�yy*}��y�Ҋg�	�P]m����Ȫ��^�uf���r.�?�Gk�&�E뉖�i�]S0��e���
�okE���?KY��E��J|b@��F~��,3D�be�	��5�>�uPH�궠�]X���1��i�����r`s0�}�	N�AE2�c�� �W���eE��'�:Y���OY[vx�=������B��I�̄)�j���� w�R��b��z4ۘ{u���j5`�~&��*�m*,uZ�ゝ�����-���߂*ϸ+�.���B��H	����S�zx%��)<�Q���g!5� b�m���+�$��P'�\l&e=d��D��X�mA���^ 5��2(?c��yU⡩=���!���S2��4��>�Ӯ%T���L�f.d}<p����)�Rn50�?��j��Iu�ȋN��<�|A�T�\��4)Jk�R��/���^�*	���
I��m�u��Q��*gb-CӮ@�%�.{�=����(9uWW$~>�V�´ù��;<��@-�j9����R5,c��� �Wuc���LC"�_�_�I��9�`qۦ�oM�8��#Cwp�V�)�Y��M��8��Y��	�Ok�>��0�Qv`#G"��?h����:i[(Fh�6:J�g���'��Q������8����\�!�~�C>�5���h#�"�ȋLp����_� N�Z1���J.�������p���5S�x�[kVN�#�
�Od[e,<o��hP.� +�k�)^&%����/D{Wǚ�|�N;��_�,�VDڣ�eW-]J�Ǝ�2zF��J ��9q����I80g�i��N�j��d*:1���M���b��_��ە�j����S$<m{b������h��}#���jܭܜy����x??Q�W�����ca���^9�g��Ǝ?��7�=g����r��E�IwZ���=��T��t[
�f��u�7�~��E*��X2P@ZN�.3�7Y"@~�������Ai.g	.�=��}�����%3C@I	-�s�}�H�ʅ�`r4�0K/(rR%3Yj���VS6FE�=�W�:V5�F:4���qD>�K
��nI�Z����+���r'����t�)�E��5�0�{��.�A����Ϯ�q%c�Ž��9��o[*7�a�	t�'ɬ�k=l;�8��3�:~�!��1��� ^�N)�9�|领U��]�ܝbd�cf�y����Uѭ8A���*b����O)��������p��M=d���9��%I�&]�jQ�rs*���\�g��R��U=�q@X#�\��t@j*Ԝ�uHL��~C%����=� n�a�$�2Ҡ�u!�\�����o���[(��j�c��Qlm:,¬fmR�ثr
�y��*�n=�2�?e,�E���@��Qѧ�[��x���.�@D�T�#{Ea�yD�p��6��&��k�o^�>�k��:��/NUy �5�t?һƦ�hًom"�=Qs��w�tsyo�G��Rhw~�\	`���6#�����y�лhs�0�{ ���h�W�U���.��-�� ��DB�m	�x�'�q������_���Ɯ���W�Cb������E�ܷ�L�b�^�> S �ʦS��T�UUK�G�.���������j����(|�X���l���C�]Q}�p|�!ԠE.[3��A7��֥#�#�ȴ�@�[r��0ˏX����tT�����.���;�+�E\=�X4�ć������^v.F�I�sq�����O%��`����
�)-\s ��do��_�W�ن�1q���ۡ���14=�?�O���o��F���!�˅���G�����V`��-�z �-�þ�����e\����wD�h�sιE"���6s��1�,�����m��-���3-f�p )a�ra����n�x�l���a�~�7�
�lA��^E�;�c�v��{3Lҫ,ː$y������ا����X�=�.}e�9O��$�>3O�ڃ8����s�o����g�i��nLadD�I��Jj�_\�	�ڦ�zo�^�FLůN�s��p~����ڈ��j�N��
W�c(.�'V�($�;�l��ƅ(�%���ђ¦ />�m�1VJt"�["��i��>�E9p!�e��z�K�d�����p�h��hx���Nw=u{,���o�G:.�s_�YX�mVa[rʀ�R2�_p�:NυN��z�v��&Ŧ�쪑o�0���j���-��Q�m[�A{�A�-��kRj �C�X��p�cݲU���\�����⑕c���d�5�1cD������{w����5����]���vm3{N)�d�d���`���H�"�S�@EFk#M3�f��M�8{��H&�gƍ��b#X�Bm5��:����A3��h7k��$sޫ�0%H�l��#A#���}����	^f{�~�}g{�v0�6�t5=���s��1���u�;��E�XA���I3#�Xx氟��3dϔL��v\ H֌�](
e|�>C��Q-l�Πm��m����"'���E7�Q�j�1��&z����9��QV��@�ژ�[�UnVH�&�Î�=DS����S�A����mmH��1+��lY#�{}o���X���C���՞Q.3�B�ԟ�|ʛ�����&���a2��_���e]�!���O!��G�"O��-3>I	���;k5T. \�C~���J=Z�#���$퉱�$�dBU��R��Zx���bk���c��*"Jy�"���7�1?��9�b�g�?e롾�e�~�0vLӀ��׸�.�74��ZS��z�")����i�ә�u#z����٨���RN��0�i�#�G����CTi�e�B{�e�@���`���ʌoz�`�tL���޴]Ŕ��iՙ(���_ٞh���l(XU$��R�����*�8�,�滄cW�)���l.�{�[�i_�9�j���W�O��zw��!qջ0�������=h�n)lT���V�����چ�C2kC%a]� \p���>��;K�5�!�Kd�N�.��YY�F�p*P�J��ob��À�^h��X_L]�J��-��LO�63��M���\�̽���F̀.����M����4IP����_�����%턽��~FZa�J$A
�W)
У��}����h9Ѫj�H;$`�>�� �61J����:��4"�[�{�a��VBL��.D�(��2��I8T����&a�T���Hă~$I�y��	�����U�iN�iI�c���@�B:"�T��������pnU$\L���B�����#e#)Ź���p�h�ؤ������(���Ԛtyq౾)��y/�-Y*�XE!�#�ŶO�{�!�-ވU*C�\����P�H�|/����.�7`~X1��_�m~����,A�Һ�KW`�Wg�?��^�[��3+�{S��E����eKZ��P+Zϸ��S�l����G	���X�䟈5�]�~3�n^��G�7�y�}����y���x�	zV�A�N�+Tك`���~�2���4q���35,GF*�v\ 9���mx�B�7ǘ���a�ՁgnP,�������^�c�f��v��N��P�dY�ꇅ�h�f�p`��3�e?��)�=�8 �v^�N�xӴ��V^�zi�&Kv�\f��S�����Ȏ���-���]��'�0�<���Ջ������U�-�
�%da]�ؐE��
Q-̧�I�z!���e����B��̻�xvG���m�M�I�W�����z�i��p�kz,�:��x�T��D�ڗ d���� ���=�L��ꇃD���*ˣT��B��sԳ骥01�N���PG7���92�]1�/|�����������.����*f�-uβ��� ������~˻��C��������@�oh�g�N���M��>+�&vA$%Y"�R� }���5�)���;І��P���P������\�
�n�k�� v�t3�,����c�T=�9��$���� �����2�L�L�������+[쳕���p����Z�[ϠWvd�ڰܖ��A��<�G0�ư]�⧷�q��!�e5|���ϰ����쨨aO(b`9�qe�MJV�-}^�Z$���%���1>ǡb��[2��6����3\����E�a|HS:C�_&\b�T�6����]=� ~�`+v3�Y2�����J�=O%�o��oe� �N��0����-���EÐ�O5'������G@ʨԝq�C�w�g�}2ď��;���[��p�˅�_
��N���
�6�ՂŢ��\���g=��QWVoA����[�����'u��&�l��bK�k������y�H��
M�M���'�j#��;�b��%�ů�KL��(y1+��r���  ����`Z28V����0���i�ݓ;U�0��d���ӶP������560�*�y��%'ԢW���-`�A�Zh7GMį ���W��ӽ{E8QT��Ԯ
9$�WVJ�����ZZ 6�}0
VD�"W�bC[�� �Գ�������5t�l��R�%�i[�ge�U���q����!�1���ڃ; f�Ԑu/X�K�;�\̃�K^�c�I�)�c�϶�F�����x'R��l��	+J�1��Ty�-�?�=�"��}Q{U�d����-#�_�-f�I0�bֶ��e����m���	7��5�d��ϯ(ë��#�xO�"��Yg1�Z�GDFG�9������VL��&N��ꪰ���p����X�9!_� ��d=�ϐ"%Ri(6�օ�C��c��.�i�6�aԓ�w;�78Ee;_rE5J<p���{��v�z-2�ԌC������m�j�\��%��~.�egU:&��]�� �����#��N��O6`~�%�t{iUݗ�B����Kv5��Y���n����Ǹ��[,7+�/5ٗ^K��8j>�G�)b�"-�w���F�碅`����I\QQ5�B�)�Kk=�ZIQ���o:'kͥ3��&��N�ۨG����
�q�1�C,.#YA�aN���=g�[�n��k���%#[��z�T`��/��6�s�׼z:e�ﮘ�~�c��PFl>٧6���V"��Dz:G�݌+�<6�OT�۟@3�k����'�`����p������q��$-ߥ�-(-�6�X+�S#rZ��'K/ɢ�5��O`݉28�3؋�����e�a&v�r<}H�5�I��Ѽn~V��gnaű�L���J�T=�~��A�\�V묥��w%:��Z*�A�r�1�����������_��?-x3ok��	������6S��jN)�ČR�`�� <��*;E�Q4��]��]��H���X2�-刎���˃?j�5 S�Y��t�~��<yV9_&BnY��C6`_q�_�	�mBb�.�~�:��2���;Ƿ8ze�r-R,���0Y�u�__��B�TJQM�4��܄���qĴ�e�����5��N�Q��<����r*M.�I���<��Ԃ�^O:4μ�UM�O���N���l������N�.��\�����4~�7������S%�\G��N4�1�B��3n�3�֒q�@#:j��p+��M^��/V=0���l�<��v��$���͂�yC�xS��"TZ�-0�wG��dy��!�䮚ہݱ���K�n���4C7#�20E^`���E}Ė'�pM��8"���>���M˺�&����<������X"�e�i�C����-�W�*2vӲ<(&�bx�
���h��[v��s,�et�dՔ�0Dm<+ܩú���D:t���y��J�i���l:���ó[s肎��EV��ɨ;�Kd�vS�
�m��o�z-}�w�4�Z)v�[3��|毨�vp֗�VB7��Q���߆�x�a���ErH=��&sʡʎ��5�J�EV����R�<wK�kq�CgA�՞Ot?тO���RU��ҟ{����D�{���x�./f���rI�Q^������M�j�����&k��"Sf�|�=�o�,P�w��,)��n����HO,��H��Q���|����Q]8?�&?�s�)���[��]��Gn��!�i�	�4�͕^
_P��ek���H�q�� _W<�*W)��SK���/x0�T�D>�Y��Q;W���8a�uj��JUo��2�؜ݝ'(�"�36�?j�0qӫ�\*�a�k'.^�Hh����܏�s�����&�n(�c �|����L@���w)=���ݠ���l��'I����: ���#�\6`����i�̆[6�4������6�9�K�E|����������
=�g�z��,+k\��:��	G]�_&��!&��5�,%s+z�*�*!�����c�]�!�t)������D���Lu���?��k�t�yJ`X�� ��iQi�&�*`�{f,ސK~� ݓl�&�޶rjUJW��Dp�8�'���,@����?�F�uIe;�~��K�v6�]��y�/u�R�颈�[�H����46�k�c�9�3��R��o�O�j�@������%E���0���~ �ؘ����D��z�^_<_@�<x
/���x)��n�!?�8�F�R�is���"K�����Xh��JdN����=aWl]!5 �Gif����u�>�����6����t*!��j��H?|�x�C���o�>5�ٳ�h�k�,�.�9o,#,�za��hj9�����b� �7�ֿ����cI��ٔ�� h"��*�}�=y p�������l���\�u��Uޅ��"]L��k|N:RZ	h�o<��Fx�\4���9ȝ�&�-�<���c8��t�@���F3-����H�����o�G�Wj����b߮�ܴ��ݛ#T��5�~�+�ȚP��-ç)NU���[)<��;LH��k�qABs��W���G�m�[w�A��-��7�M:�jOJ�M�ʡ���l1i�]X[}��k�5@a@�{@�8���8�r�#8P�͞���o/1�%��r6c�T�h���d~J�����gf��1�E��/8�ol�9Y(P�ḃ��� �!��	����n1��y�G����ޟ�� �㬒̍�����h�<ګ�&���=���[�˻[�U������� z��Nt/��s\|�p@_F���婽��)O�x�z�g��?a9��svE����f$��>�2�N�K�'P��j"V��d&�����?�/pf'�B,���i2���\_���탩�M�9��P`�J�\1�-�.���i�S����D�M �_�a�w��J��ynr�:��b���l����[]�#	����d����ȕ��G�����S�eϪ��ߵ3��>*�{�������,꘳!��[,��i�-u�УQ𖚂��;1І����>qf���W��}�՟�Ej��!B�8�x�M��\�)pPNO��ŉI��{	�жW�����DR- )ͷ}���̒"�Ń�;#Z��1j8���W/���d��\�N�KsڮĬ]C��؈����/́���(4
qWV�u*���
�L���U��@b�`�7FG��~����7���BLȀ]B@�&�Y�.��iω����s��7�Y������#oٞ���w�J)�
};�+�t����t@I�;���7[� ����k��~�>�@������` ϦD~%�����>�8��<]�O��K��5�^n���}��JWO���+����P��B���J�r���.�%
�C֠Ih?j�������\,��.=P���h�:�?E�ۈ��3� �,g�˓�:�ڛC%�&t-Tޞ�ˋ�!������@��B�WŅ����9r˘��؁a�<_D������H��{�ԏ�j;��rQ{�[�LM�f�Q����9��H/�|�+� �R)/�I�yt@#�$�U�RF�iO�?���q�wB���=g|G�6��n�Xy�:���B���j�Nl@w��Y%��_�#uh4�����D�N?_vΗy'O���jB����Klo���\�^vI���s(�,�����mh��@=�8�XI���칼{��ٛ�L��p6怴m���M������Z4��尮��yA`���4��� J��%��W�I�ټwf߮}w}�'���1�~I}����B�R�i՞��hg�غY:���{�JG"����f��q�*gg�h�p�O|����r�>��/�w��?��0WZ��G����I$��\�W��K��پ���8�9�D|���%�}B��M5��N�m�bn�2�>8i�Ծ9�Ũ�ݑf�o�e�Eof�f����7���h?C/��v�8���|1،"����q���6T���p�Xp5��Rp�]��]���noH�2�pXG2�s�k�UO&R���C��Oh�I>�vR�oIi��������,�eY��9�c���C�Jf�����b����i&d@��\�fN��x�X`D2k )jQ'�h�L��r�D͢����lK%O)l-��N}C�~��֐AUJ+�Qdt3��}r�hE_ SC�I�=�bu�sf>�7]�����SW��+����(3�mAֲo�{	pV����5A�,(<�t�F4;�����)G���ԳQrNA���׳�B�&O�6���k�Ys�<g#�~�9�E�x~�O�\}<py3W v�<a�����5ʘ,v�4`e3sH�,ݴk��a8����E:-����	h���,�|ɟAg&@�~�i�j������a�XGz~Nt�d���U��Pt�˭`�u�D,B�������7�L
��]�ET����}B��a�ml��k@!KV�C���EU�ڼ��;��ցO�<dJ�$j����11�ǳN��GC��Mnd�f�!���_R��C�I�R����i��Xk�����y ��dw�*I�}��p�����B��n 畡^���dG��㩑4u��	:s���lx���.�~���d�_dƢ2���n�q.�F��5�bE��s�{0�MGN�O�?*���/�I�rv�g� ��#�c>�i��h�U��؜�9���s@d'�&�h�z�?��y��A��"3cY=&U�������:#(�/"� h�)d\r�@��>�i�e"+Gjߜ^.�]�k}$�T���X��tiM����|8�8t����������=��_��c�[�|LZk�t��Q$ 4Č��
+�ڨ�����_W���}~=��Ch4��ˡ�Q��r�}8�0��򐑯����c��9���	���|�4��>�U�`C��fħfR2������V�M"���������o���['�6��a2J4�&�Ǧ Ǫ��o���e/4������F�0a"8A?b#�c0�� �ݢ����X�BM�P̏�';J�P��wA����M�5�8����-礅��)�����K�:����ӥ-���5&���N��hR���	,3X�)�h?x��?a�~y7��v��UN�Eh�������<AP��?�^�����  �hQ���\��GA��]�X��Ļ�%�ߓ^�3);|�՟��d�E����q��0��({J=�r�_��%�̪�@C�f:.�b��EsN�*#�eԟsi k����#,�x�=QW��v�%�4Y�q�؞%� bf�p�vhV�4����3IԄB�5��>F��X'��̤����t�rd�Ch)E�y�i�_࣢��1���Nu��~)b��k�a,�x���ڭ�X9kJ����~��*~�w��lߛ�̤��;A���-naIO��e��� ���϶�N�LW���+=4���7"a9g�M`"Z�Ę�v|�,�#q��Ϊ��/;D���阜�Mi�i�����w��P�1�~^v�&!M�R ?�Y�C���j>9C����\fA��Y@G�h�/�nwz�	뷕A����\�0���E�M�� ���SF��IޥE��SX�1��W@�ebYM��Pʊ�=�k�<L[S,�ɍyӪ��UCO�����HY��L��u�R�?1ڡ͗ɕ�gҗ�F�z���g7����ql��0К�[�l�$��|�/}�A�%c��T�L���j�匪��U(DAoy���(�V;e�X�7�;L�qkOu�[&v�4��F��Uq<�SN��Z!��V����-��}(�b�f;�����v�K↶�R�%[;<Ь{�߾�j����}<9��@�}��B����@�f4RҘ����$[�~Z�ڭZ,WQ�l���&��m-T�B��ؖ����C5j$�RTA�iM��q���i'�q�;k�ھ�6��X��������O��R�ş>s���`���)]��L��0����M��Bj�Y���q�	�C!j"���B�w��{������������2�E����ı�{oM�����n:m���<��Ȇ��o�O�&� �"��N�ѱL6E��\�W�i���V��ؘ��,�Y��u���ܫfG"�i����w�������SIw�����E���y+�!x<RER)���'X���p��j�� YGK�@g�a���(?�r�d�
W�I��22�C� �9��r%���Z#jկN�F*��8Ǳ����}�xFj:�}����>���W�P���Ӝ��ZO@��ku�V���,�v���GI�:��4�φ���e E���e�:>c�����i�Y��$�j�k��S �PԴ�1�/9��/��ۻ=���j���`�3���\`��/��o�s|����4��D������$?��ۤ���Ų3�( �u>�C��-j�C��Q9n�:�U%d02��Q���&��5 ڨɞ�<( ����x���7/�{�S��9X{ե�=���O�-96G-�}�6��b�{����FE��l���W� ֪�+ŷ~������Ӛjj�zJ�Fx�8���9��Z�6i�����Ő�6�I%_��B~��vE7���Ș������`����ϑ�"��[�I���46�X�R�0Đr*��z����YY�)�D�V�~�SS##�L%�8��υKA��#_��!#f�YXp���W���X��Bϖl��܇�=���P��J�F>���ü���0WѨ"��jLC����fA���ĶRpm\o�jYN�FI,��a���Om1Cڻ����~����X{B�䝄�6�,F�3���e,s�][��3pףc���f���WdkOE%\#p+���檙�&���0�k9�$��6&�.�&U�.20oK���h$��}A0�)9}��}�<�2?͸��0E�7:���<������h	�,�c��� �N0�{e~u6'��'e����)��9Z��f�>&��[=h�sx�'����K�Z9O��v|��@���Q׷��+0�d���9/���K�5?� /ؐ�O2��^f�斶�b�#�P�`w������"�!���T��q]���"���T�vU�(=U�mnR���Þ*���7��֓�ؙU'vԯ�p3�\�3��[�����)�mS"��ݢ)aV. � 
W��JO���jq����c�w�����*��(���Z��O���<���o����]=&
Q�����1�����@��c�B�.�O�X���-�u�H�G���ˠ�� jQ��ܘ��TOF�ωS�������i����k��Q�S\�=6ȯL�C�g����lBݷ�V���yU�Ua��ص���*(sto�gQ��@r
	 ;y2RV����*pW��(��恨	�>sIĹL_@."$�Y�h���x�y����$�e�5G�xt�=�b���{�A��Oi)!(�����u#Ž��PAl��ٞ��Tj0}������zP� ,��$��,�_�2�[��`�?�&3ju��A�Hxk�x+����5�����&
��0⋈�,9������|ac�<��dn6��'8,��c`�U��5��?m��U�/Ogؗ���X���Ek�� ��K�c:pM�,B��/�'=�جg�U�����k�E@آ"�*A�H-��
#b7{f�+~T�K�)tB��ctL��F���򩌇�=o]��v�&1�&OK�ްy��Z '���},�Un��dJO�"s��$���|h(a,0����N:[��$��8�3�������	���/p�1��{5�43���y2��q�s���(�T�j�u�:N���v1�Xq��O�r T��0��!Q{8`�X�w;�S)>-�䁁cpX࿀I��я
����Ƞ<�A�Hf��"1�����dc!a�3�G e>�,��	��|�'aʩ�p�"	�8����I�z;G�͌�Z����x�y��{�p�o��;�a���H!џ�᩻�ſ;�N�P��o��\�C�d�z����)+,������J����+�_k���EN͆S��9��t��nR�� �O�L'��@a�Q<�a`v����gz2�W�� ��-���H#��r��U�rho?��讘*3�7�4��w(h@�4燓����l�3�3)�̗���j�>FӼ���,���BɇL����ĳ !���u�oZI���TF�͸e����͖K���d�f.����AgT.�\�Ƭ��IȲ-T���]�"�U�_/TB��d��f��Y�64G��kti`��H��!_	^�V5?�ƩY����p��X7��'#o��j��{	��S���D�)�ª��5�*X��枍�����^�7���$U�t.����CY�]�-��'>eߢ�G�^�.Ʈ2��, �N�qC0y$k�Q��~D%�3��T^J�GT�s\B�|�rPm�~'����ִ��GHa�P|]К�E��TG#�/�HZxġ?F����f"���E���o�b�q��T�1�2#�.xǥɃuE�z��Ӈ�xv� ��dD}�Z�V6�d$mό�<.�
v��!\E�V���>פ��Ј��9�!Cb���2#��$ԩW,]�r)8A�o��2��I��ȲG[	��U�-��Zl�I),�Ϸ��3��x�9�[8�H�K�]�>�o�m[=��}	�B���(�u�D=Yo��2u�V�zp.��)�,u�8u�z�ȓǯ�7�\�>m��!}��ῷ.z�X�l]j���}q��@zdcŒ+�ګ���	�t��Zad�Z���BJ\�}l���1�����\ oXZ�I+�:t�{!�jF���W,�XT	d�#��K)L[��c�K���uΠ��������,�/�j@!n+��	�3����06����ǚ�h*��;L��Ml������ C�s��.�SQ��ܪH�u��^la~*[La ��/^a�S=�̓}y���2L�t>O�S�mμ�m�kZ]3�
��I�&�a�瓼)����9���xd��i��.��Q���S8��I��˥fXF��}D��6�l�h�E�8f�t�1h����. so�ЍFPy�٩�����2����n�{7h-:�n5K�1�!���B"¸W�{�f:<�J�Lw��p�u����!����-��]�?�ܩ>��vտ�a{fV>���BG�z��1Ҭhy/�ё�li��>ġ')���Z��YF���6���t5��;^���*̇�n�3��J5l$k>�T��e�
�5M<��t`gvX,��Z�e��?�ʥ�v*�3jS�j
�u���1�
��	j|k�N�<w�z���ߔb��LV��q�}M��qD������N��F�_.�ږ�R�s�hƣڮ�[���n�=i�P��-�^_�=~�p'��җ"�KE�	�������l|C{_2K��2P٧5��|���<T�ݟa�S��\��|�#�wRM:��q�9֊�wVt�m�wB	+�ъep7�~�{7��l&*� ؓ��,�od>�ڂǩ�躺��|{�0���ix��iɇ�D��{���߯#r5��6�h�:���\ݞȉ2)�1�k$����03$$ku�v|�	�D,-Z>�b
N2f��X���ƒU�����ȁt�����UݧH�҇pJ�8�J�� =�ɓ�Ai�0g����-�k�,s,�?@�z��j�����ٝ�!Ĕ�s�?�e�cVI��L.�!��?0�P��|�!^��9ŏajS�)������-��%�{K��޸g��u���X�E j��"ɦ�!Z�D[��R;���[����=p��?ᅇP�S?�)�Xw�|��oZ{����m�Ȓ�����,�kUcy�L����@�vg�\�^��R$ �_�8�� 9���I�r"�t��d��'B�aGk���R}O����~�?��Â�{�E3�����ߛÄx��;O�z4=�=]���E�٨$O%We��Y�`��g	/��B��\���l�Lf��L5���oX�-o��XLT�n��X$3�"L�Aw{�^sF}�����X���r{�&�G�-؟p�*k���Г�h�o	8�g�.���n٧�׸QF��ˬ�����{r�X��>���^�u|�Ke'�A;ʔ��!c`�$l��^`u9�%��X?y���}upΊ8B��-���]ckή:j. ��R�s��@4��{��[L�-t�{@�3E����ny�Q���7�S�L�(���E���*�$��%�L�%�xQ��q��ʺe�*i����>Z,G�e-�O�|S��*j�a��׳�D��դg݉c��/�#��nvXU�u���Y'�ߔ�������r�ˉ����D�~������ōe�' ��M;�� "R�"|b�mP�-B/���:r�o������ֆ��� X�r|��ˁ�+e��Kf"��@�J���,$fɔѸ��0��S&�9�&��_��l�Sf��f��2��駶D�M� 	ȓm�l��������)U��X��"�m��p�>�E��R��:'W#^?�x�hv�	}P@��&i�O��R��_�w���1{5!yG��5oH���ٳ���j��eǽ��gC^���!T�UKԜ��H����)�\��!����CN<hpz+D�۲_����. `w�[�D���b���՘�]	U��)Z��|z��e�p��x@�򩼸�WB����\�f�|�a��Հ�,17�9<�3Aa��8f�K����W��(�a�E�����^kb��~�3P�>�EH�@AeJm�������S�̊�ychp(�)
�����EM�����e>����N�XB,�:�ڔ�*��MJWU,|q\�
��A2�3*w��o���mX�g�s�ؼ z��& �'� �m��=�(j^��U	����{3�'�M\+X�6�jG`�%Fl?8�-���g�k������@�T�a"�)AC�o��s�ft7�,�E�G��Jל��	���9%�$B�d�NY����0(�EeW�]��knƞIU'cZ&Ò�e��궑�h�`��}36��O;#�g��f=��Ӌ�ޣ��,��2#N����{�������d���� ˜a+��z�b*�[��5�M4{!a�}�=��q@g�xd��zB;���@;��n|I}�A�,����H#)��������#���^�0�%Г���u1UBWw��%�����[WXS�� ��$v���ÓR�Q�:4�?��4A~��E��H�������J�8G*���[?��K�� �~7�i{i�+���Zb[$��� Hѻ!V��(�`�U��!���������	Η�I�<F�z�%I҄��0Y<!�H���r���%�*�q �H������y�� ��J��s��`�d>f�{���P~�U@Ѭ�$�=��P
R�N��M����]P�B�j$z�c�>���2�h��44�z�`���+��V�ʆ�~�[~i.	?zn�^Kt��]�8�^�4�1�9<A�;F�؛�KnZw���1w
�m��vu�|��;�w�f�$04�GǴ�y��dj*�~�I6��b��J����x�f:�з�آ�j�'���0h�Iyf<ؤ&��S A>��/tF����7���k��PnL⋜^ҁ�K��K�ts�%��E'��BOŰ�Zn��V�dO��j+ų!�-;���C�����=.�qjn�	�-q
L��*�t��� �[j#դk�4�`����Kw��˯A�Q��ڪ.9ë��ߏiKS�K	����|�?�?"�j�~������W�:΄���Y�0�ɇ�.%�{7������l̅=���s��-�f�B�Ȁ^b~�Y�Kr;[̔{9���?���<�*'H'^��}!fWT��/�v񞽚;<�qq�����$�ߩ��k!�
�����>x'F�+�-̝�,Ռᒮ�UK8������M��2�>}����&���=׵�� �/WT9��"��r���^�7���!mǓ6�יa�0�P�!=�N�I�(f^�f�Loau��䬕U�Z^ۅhX:��ۚbz,v�� ��x@�63�hry��&��~Cr�ŝ�K��|N�R<ڀ���P{=S�6�����5�J&^��L|��n���/�%h�Xy�&{>�F���nm�� Ϳ�.�F�����8a�W����3�P�����B�:T�<b/�RD��T49\ Ȯ��ؤ��EU�?V��$�����|hO�b=�V�6�>����6�_�֎�}퓚�i�����wv���K��z���R939�J賮%Mo}�����P�H0`��R28�ڣl&�^/`����s��cϏe׆�q�e�1� ��.�FM9̽4R[ 7혎� ���u�k)0�����,Dʺ�G�-�r�I͉uX�t����DAcD���d�T�vS�q�A�
�	��ұ���ˏ�y�|�p/���p+n:jAH::�5����iۊ�v�Z����|Q�kqC�.|Bp��˙���#�Y@0��@�ɟ�f6맹�l�6��H뙝	�)��b�e|��������ǯ�>ʧ���x5�/]zS��(ͼ6񲀇Xe������7b&"1_����b|��k������_= K���'��Ae�� �'Y����!A@z���1}�A/�u(f��ѹ�7�P��k�Z�v1�����	E}L7p �X�-��J�n#߬XL~��`��1��u�,L����θ�1t��F��u�����~"�K�	s��h��/;��45�^�딯[�rU�Vi�4E���Y@;~x����$��\���tk�dUM��B��;����v������s�k4Y	��$_��pC���(�#k^�I��t�B�q�=��	����FHJ�=�Z� �~c�T�T���Q?���vb%���c��������5����BG�i���x���V$��]<<En��
kN ����BS��>�a�%�3�����rz�hS2(�Y*Y��\3'+Y�]W���v�D6
RTWk��������*����g�����#�4�����'�Z|�$�%O�1��=�| e �wL=jU�`��*Х����}���篙u�����5�	�3�-��7��H{ku�>T�q��I�x=^[+w�)����6)�h-�!���a�*��r��$6m<<���G&�JQy~E�*=k'�>�bgN�N[�ͬ����#�z�bws�^ΝPp�Q�6)#����3T\*�l����F*9�r�$����*�U��XG��d�ˬ�Gl�鉡.�c��P�>���L8>�n���`x�(��{��s��N�*���9�$�/�`���}v�H�3�a��*��ŋ�S�<2�x��\j�n�V!;�	>Eu��> ����z����Iw��s��x�d$]���َ�@�4�GG�T��L���& meF�7�c��/��$��ۈ�ZXݑ� �1ϘQ)���1�G������NS}HQg�PM��Sp4C�<�NԨ����x�R�1/�F
xT׽�;�w���w��Uz��R��B����o�\�v�D�6!Z)�%d�Kj�k�KaW��#1�'ּ[�&=�@�gިm�.��6j�������pR���}����V#�h2|x��V�l�<�:���GH��鳹.:!�"@��g��m��}�x�8����V��yI���[_? H7�O ��۴U��ʨ�O�וVc��E���i}�x�B�~�0O��;z��ˌg`�X�p[�����8i�r���䔊���|y>o{q�A�L�~��֡�,
}�((���x��N��`2�1��{Ͽ[�:G�η�Dg߃�w�����"O�O����63yTԼ/�V��Q�>㰏�
 ózؑ�pC��4�_�n���|��wf�ň��LA��]*�����o�Y֏M�Y�)�P�J*Z�N�Wչ���U�Ow���g��S}��W2�B��O[�����ڑ +�6��0���uX����wc� �������>�T��3�rk�L���,�.֧��8�� N`	�z԰�Ee�����'@��@}D#�/w����&�4���D=�	�R�� cH'�֢8���n��k����}��R?�-��'V�_N�t��l\�����ּ.s��U^ձ�r;���1&A^�tѦ��kܾED�7���_�i��t縌�h�5!��Q���~򟘯�����k�qm(y�y�MF�<7�T����`��;}A�D�}w��s�W ���e�o]D�#A�3��4����Ia�s~(sȾ�Z�X�4�1m�<R� �\[B��;]�e����� �r��6�Q衭�@��s�;嗽E�8"i�'UTͭ�7{���n�8t��z�+:�5�x�ԧV���V����Ctm������G��u ���ذ��#��an�!6�褕����ze���ˈ�?t��#��b�"k���K���g��G>H�����S��i�|�+�k\W�w�J/Ԍ�ޗ+.d�&A	��S�"�)1��S�y��茎�o��n^�����v����NEG*��f9h�� �^ckO���'J��_S�;IL^�M@��$��X�C��S���y5��-T5 YR�yEX�M�7��o͖*��@�-܍ԧ���'zO|�7�3ߋu��+�8��S�,�IY[�������
�$2�"��3��PHY\/#���?�+��N��_,�A�O�����;��X���~�LgbV������|a�&'-�V=-"�]	����I�YA�k�ק��p�#�n�����wÏZ�\��=��竧[>ꠋ�� �7�{Ǔ*�Z1=�����������75�FZ�в��1掣I��,��_��:�.%|�z0|�����>M�ST��%7t�����i������S��\@P��l/��XV�y�c|=��	�9LE.K�x�ߤoWq̩����h�E�_a�n�L��:��L�{FI��$,-�2��N�I1z��k��y��/�������]��m]� �KY�"��ܴ��k�W�t��>OG��L	%z�c������O�"��@�b'�)JL�w�1aI _ѩXԁ=u�xC�0����7U#�5q_dŞr���'�ӼyA��R+[s����w]0́D3�J<1Š%q��f��
�8U�ݢ��+.��#S�Ʊ�Ga4�|M�}{�PX:"#%�]"6Bp,����C�
��֠>6L�/�ޗ�t�fD���E�hX���@�*���E���_���0�Ҁ]�{~�
t���p��m�¶*3/@�A����3��z�x*3�H��zrgG #�w\���C�d�~��� `%��o3Hũ�9��
#{��4bl��n��(���?"�|-22D�u�m�t��[�}�nP���^T����U�NW��7h��3PIJ5�N�{q�y/4wN�6���&A��o9/����M*=�N��}�:�"o�AN䯵s�=�Ӑ�Jy�8�J4�K�� �嫯�MqI+;�'���w�0��l.N":F�.^S��P�.=��r?�[���@���{>��{�-�)e�C�r�+����!X���j��z�ҿ8��<�)�4�R� ]��b�BU�'�������GBG����y�*���g���$d�?P¾+H���.u٘�@ϛ	��l.��kR|If���������^p��CzO`Fߕu�-+S����[��x6�l��"@͓���-��1a$��u��`�M��
��8��Jyu�s�O_}~C��z��5l�?D��*�W͠��R�[�<k���<ﰚI�_�ě�y���) % ��g����r��+�Ot��>��#�-B���j9[!�R������Bʇn�u�T�S�V~}+�+}��=K��Aw��� l�r\x?Ϫ�}Y�_��c|��6�V|\~{����v'C��I��g�����i0���}����O�Bj�/IXweC�҂P0 ���[�BB�)[�\�r�i>�y�=���K��F�<;Q�%=�Yq��߆���-q���"�tUK�k������[L��ް?�Z6W+۹��bʫ�*�|c)�j�v�K=.��"��i	{a``v��$t�P���1��E%LЖ�З\�އ��X�`X�*m\S�GBRl7����� ��c�W�1����,۲�@)~�w�iT�����yc��0�) �d��n��m�Z}Ɛ෇)}RI#��VtN�u���=�M�"N'^?�b'|;[�dr�iu&�0�G��r��1;�Zg&��L�d��`���1�_[4���۔BMV���������_y*M��w����f��tL(����F Ft �G�Y�19�bԞjș�JÊ��0�[�Z�*�����?�1gY�����a���#p(�ҋ�9\�8��ic0k¥�_����ݙ�@4YFt^���}��So-���s`����`�� }�|U<��j������ab+������Ճ�xt)�⢈bղ-h�<��<�}�!e�-���?���«P>o��l*/W�7���� ���l;�'1���f�l3�$�k,�r`�RL�`�Gl��~Ws����۬|�p�x'��T=������f��+�\�4���E`Cc^���gh��W;�"����Hi���x(��?�#� ~"�B����kď<C(�P*�2[� �g�b��B�#��l}���Je����D�)H>B�y,�^[�Iq)��}%G�&>���-\�5�u[��`�AA�{���7JR��G�] s�D��\�ԝJ>+M��v�c��-Ô�9 *�J����C���pIS-K�A��z�HTI�ƪԾ�$�#׵r�t���l*k;�w͕�#4�K4�ℛ��4���>m
�Q�O|-�V���cZK����:wǤ��Jj��GJ�mG-kD�-������4�v��%	�C��Q
�K>]����!90%�ܥ!K׾�\�0�r���Ǹb�M�m͎�F�(��{Vu!�¯&���\�����lҟ�R-���/|m��.�C�T<�+�c��p|,�a������I��*h �7���]P������Md������g�ܝ�5mD��zȕ�����z^*W�.�r��H'-���iڶ�}��zkƶT���.�)� n��'.�^����_�����:��~�=W�<#:���ѵ� '"��JG��q��}r���f��10���u��^�����*����d�]UO�v�����4	n�������Œ/�h��)��F�LՕ&����o����M�Ép�r�H$@S0S�.�b�d�P��5J�F�J�!����c��ȝ6�,V���&U���4Aql�,�Y�p������It�49�����
<����
值�F3�#����3��):�`S���1~�3�	�4�N�<tO�p�jKw�U���_%���6����z����Xn�$�ZA��1��w8e�������:i��<}�iڢ�����YGT�>1cB��<`�7�2C��}N�>_�(�C��A)��h ��q\8L�
9�@�1߬�tL䫍�yM �`��w)�0<_Nۿ!�|�pA-8|�Jn�5����4Зi5�B���vlͪ�
6������jl���k:�C��i/��yp�h�kmT}@&>�4��h�ض�M���z�o�Vi�
�c�H�����5�7��ʒ�Zt�4��:ݽA��0��4��RP�'Z����On���v �X��䩌���9;����0��qe���M�ϸ������=�J�ho��K�� L�D��o�(v�w��mHɴ�ܻ��Jj�Pu�����(4%fn�����Ş��h�k��rO����ܚhG�d��6�6Xί���ap4���"XbIvdλ����5���i���Fz�J[}�(|X�b�@���~+ꡲ�8ő���� ��H�A�:]¦6������3�u���Ś�e�f�Fc�!ꟃ��%���4!���N1Yc��?S���Z�K�j�\&�$J��^�xX���5�e�Ι}r{W�s��J����x�Y�<���J��IȈ�R���9��'.�}�A5��Y�j�.�p���VR�w�oq�T�<�P˿������,��s>�'���~�}�d�,�p�v��{��I�h�W�8i�㰩
��4��;����]|���+�6a�T�2��@*4;C/�⫁;��O�5([6��H�#�ɟ�9T9:�H�GC�xi���+}�4S/lg-H�}/	��LCK�;wZA7�cľ�Fe~~B
�k���������H�x:�˼k?�=����_J�E�q,��5s�ddW~��GhW��p8��(�� ��dm��;��zy�C�:��'F<�*�q�Ů����x��8$�CB&�)� ��Ѣ,��un�
�c�$J�>f�&��� �f {��LJ �?�X�0G[o��� ('>�i7![�U��CAO��f~������9ژa��1�&�A|�oÀC4�s/!����˝$e�L�Zb��d�F0��KCa"M�[V��I��M3пް�H�w@���8صx��� J~�'�*MO,�d�+�
��a㭐Ø���h������ɵ]R�[���<]C��>l���5fv{�&�f��Q3���Z��#8�t�)�����ʜ���l�7E�B�[U�V0�m�='�^��O�|-2�Rb�*8�����Xx��KW���E�f�w,��#P�O
B���M�|����7�����S�{� ��ZZ\�	͋'|���"�ZzطQ���e%~���ʜ��mj�JN3���HX��Ck�h\ng(G��}!V_��/��xq�h��bѓ�b�x�G����ǔ�6���~���X������c51��%��IDi��N�x�|3Q!�΀t��gF\~�ӕ秩�]���E���NBf)��42����0��'��'��C];�tfK�g�qc�>L^���S����`�hm/<Ů���&��*�-�j=�$�e���$���kbfj06�s�5��5fY�:`g����l`h9#h��K���6ǩ4dtx@���t�c�fH��ϯ�U��=[r�V���"�v�t���H@�x%:�Y�<��x���vЭ�j�<B�kŹ�!���ϥF�D�{�D��t��?�9��#!��K��� N[�ql�s�����k!�s����'B�	�7,�[�V���bj�L�!�{���v�4��KV{��h�X���M�W	����ĳK��Jmػ+V��U<� W��ę2R��`��{·��L�Ӏ�!G�y}ɷ��O�vR�Ié�Yc��}�!h9s~"Wg���4p4��X3u8�md�EL��`���#7e3�z�>�yf�x6��49/p�Rw�
b0����0��詸��\% �3n���<fɰ���3zW���Aq뜃��|�|qWB��i�S��+��6d��P�#��0�ڞ��Y[U���G��@:k��d*���L�Ff�%��x�;�bj]hn��_�g������T���j������}��̖r��Ӓ0E���XM��o���j��P!m�dse[�:����ҳ�sF����1��3;W�ڧ��Q�kk��mt�S/�av�A���ԭj�DXU�j�f�̥@ܑM($�'��]��m�l�ʹZ��5�]K�Tǫ�ݮ@�u]듕���0cFr����ڶH���(z���&���JVs�sQ�R��x%�A�;�k�[��/}�M�K��͚/ ����������ժ�v��F$�q&>��5��ԁ��+��?����t��y��e���y4�V�T4ڑ}}�f��7u65
�Wh�|�?Y�o�i�wm���:��A���M���m��Nݩ�N��}���?`�_���EK����q� ��$���OX�/J7�/��r�)��H���=5U-n��Qڊ��"�!?&ʥ;�7�Ր,�n6��"d�����ӭ����^_��Mh���:��`�#���]Um ͖�fCvN5����D��6ʠ�?�cl��j�|��dV9�EC�)3_��&��V�@p�x0���fL��ܧEHI����kG�|`
�ز����N>���
����`�/�˹F�U�t]tQ���mkS���f��"����S�]{�H"�1��6R꟟F ��¡CJ�-�t�FA��A���o��ˑF��K�����gİ߭��9N�ئ�*��Q
g��`M�D}�C#?��.������ѓo�U����O^�|�)�!W'��@��+��q���U�c�l�_ѫ�:�����2LYo&���tj�+6/�(���yf�V�;
����HM�Fv��D+2���+�t��d|��v�\ �ȋ���B��{�P�����YY[bW�ӓ �g�]��'^���#��ى��/�p��y� �ڥ��z���f��#�$ǋ��a�[*�k@�Lo�9h@  ���=��y��̯�4���)M�uEk��Y^�G����o�)�0n*zX|��	}�w_ZT	ZmZ��nՀ-�[DD(�bu�p~������������,�Ӱ돵*�A�)����D�'&l�s�X���I��_�G�uj�8\e������a8N��'�C�5U��{1��sê����,Kg�gd�����lJ�(�E
�s�7�����T1�E����ǔW�+���L�5&8CwQi����g�Q׎s(w+�(V�-�՛ʍ;*8p��V[�b�j�ŞT�{��r�����]��WPV�w9��lM��s Dޗ�}N2��h��>�? ���#l����9�{5ϭ���,%6(����6Ͳ���0(-�%C����Nsw���H���&��n��0�z �#������%'w����i�D(,�g=W�V#�	�Ԯ+�(�랎���VW�3���#,�QS�Ne�y��,�DqE�c�`ʋ��z�q�q*$m�N��n.vH�||�g]sD��kxNU[���h�P�H���5�����2T T�c�U�:����̿F�Apb$��LZ�ɪ؁	�K���_��=�N�Ȳ;|쳗X$K�j��6� �Ư
�؆�����N"iXEɟU��)ĬD[�;���6I�QR҃��8ng��k�y?�u�s�@�p8��mI^�C�sJ����	Ȣ���@��zlA�i͆��e^�h���DKX�g����'����1b�d���ݖ��CN�7S�pS2<*�V�Q)�.3b��6U� Ā_��XNm#����B̗j����+/a��n�S�(ށ�Д�cd��2��cZ���]����V.�Վ�/��K��g�I�'�<_��v;iƦ��	\��"��bI�"��A_���?|f�N�g�����x�ʂ�w�0gm$�	*�/��aHl��<��^��=g��Kٻ���#%�}�n�'�هuB#&�J*��w<���t`O��!&S1T�ޚh�s_��[����,G�R�{D�)Ub�i�nRmD$��}y�'}��� ��k3�Ͷ|~����qm�v�o� �=K��ic
���G��.�k�Ža��܌�}��-�K�a ��
��ƌ�F����2�MFx��k��B\�##m3�C��W��WKـz{e�����A��F��0Y�@�oT)42�$t�ÃY������es߹,#5����tV�[��l	�s��ɿ�Dw�Ć�0W�>�c���\DTŎ�Ho؟'	g�.;<�ÞxBwa�?��^Qt-�ycv�u\!�����_[×� �f\�ܺ��Ro�,:#9�ţ�	��O�I�[�%F�"�{��!(2K��i�nA�\J���cP-��V"Ŀ��=��˛f�*���MJM��yuC��Z�� n�+Rj��y�Y�}�@�}E���ix�[O�j	��X��]�[��C�s�V�v��!U��%�!t3>m"*�Ϭ����&I���)Z1p��f@�E��d�pL��)��j+}!��#��+=/x��/�+Z<'�y�%	�/*eEs��5��+�d��o!�k0l ���<m�p>B�54�<}K�� hWcY\J�r�K2�v��N��6�梷�`+�֛u�hkt�5����~a�#�`A��!�8E_lE��]ㄥ�b��Ǟ�^>)��[e�F���H���q~�r��i5����4S���TM!���U�E�������tK�ʳΨ�&4e���y�N��|s˭�����<gg�f���,�b0���Q�W-٢���l��	� �Tꡢ܁h4��VIܯ��u����#i	͜�P��C�w�|��̇�]���P,4�@��9�!8��c4U
(���6�N�p�a�F�|Ӏ�C���� -a��7�!<Q�`����Jk�0�����4�m=����m`J�@��.X �Kǯ�mR�c}D[�������W6�v�N �3��Y����yrg� *��>�Q�g�h	�LML�\&�z~��F}ӃMn(=����lD#� ��kFj/#oV�������8a2~�K�|����(���&���u�(ܖ���*;�> h  5�P�5G�c�'6GP8pXD�*F\���2K�AWyu�>���l�@��'�y������$�(Mfq&L�_�C��Ԅ$Q�l�8�1>�f
�Á��50{����AaQ�x��[��[����D�տ伈'���<k���쿱���b'��+�I��HM�-Eܐ���k� y��m���\�*%����Z<��"lٕ^0>��.���*����w@}���u�4���h���wh8q�]�}|^��S�S�b��G�O6�&yI���A�[:�S�(��e��\r@�¦	f	*j��;�1$Q�Gd9b��~�L� �?��;�,���Pp����!D���Y	m�/6�,�� ����ݝ�m��U9����qG(�FFR�'j��m}�l�ʈ-zҲEf"�NLG?8u��������n&5�@؞`<�a����k5Lz=���o�ʄ���I ���2����uV^�u�����Ah_��[�_��
�z����f�҄���A�lw��☡�ʵV�����z>> �g)/F�Ӫ�Wn;D�ok��_.{�����]Z���vVe��f��\�l�ژ*ʏ���7~mS?��q�w��>[�����b܊?�če�X����Md�V�9���~%�,sQ�.����؈8'I�5��~h�̾����F=>b������2������oM�s�i� ���C������E�i(L�D���u�'_f��)S�"D��n��IY�72��GN�o&��z�)�\���$�Q�s6��"	ǧY�����U��W�G�w(�X}�ȃd��#Z�zR�� ��$�E����S�mX������6�MX�por���F1���ݑ\Ps)8���b!�|��e��K �;G��%��{m����Z����E�Vӆ�Y�����kx���Q�����͂��j��B�N�F�R�-�eo ���ު@Q��]�*o�m/`��aZ��8�(��y��E����aq��l�L��
�Y�ȅ�Ýb�p��3���K�Ã�-��9Jn(��P.�����5��26�����i!gϊ��)f��f�^y�|!�x�b���$]��{6�2�� ���n�G�Bn
i$��_;��W)zΌP;<C�gI@�~y�*IO�C�&�
t�ã�ؽ�������q�1"�4�$UQԚ�6����΀������&�����o����E��t�����m��;b�NY���q��R���A0�t�(�%�Uѡ��<�K5A(����|�*X��w��,6���W1�s��.@"�w,���3PB$�>��-�x�E����3bR"�OQTE�a�c��o&ۛ��N)���ͪX�0�~�� U�j�q�0��x���IU��gW���s�\p�V�M���v����lU���r�\D�j�j5��>��@�>"I�ĖZ)��\�+o��EYO���t�ܵ/����z_������/!�a��呹�1&I�?����$�����MDA�*�����A[���m��x���?��=bK�>��}ѻ����
���t��������vqSA�]%3Ȼs1��8����8�H��Z��a(n��*�8���+�S��7���߹i,%�4��]�n�f�k�] ]DJӖ3#"��4�za�M���:�y�ݚX��k5Z�-�A��w�Q`��8��c�']k	ևkӡ$��۾"��6w.*.bM���B�[j�	�jSI�PH0�0%�i�4&��A�|b�^�q���rE����^��:��p�>��|!~�r�14��Qj��"�/�^O+�qq\K������'��ﴸ���&�P���8h��a-�����G�K%`TZ>��"�ή�vE&c��c7�a���+`!�^�8��E!�["�J�F��ZPe:��?&s����FMH�9�!�0�kS$!|��e��w�N+&�'�.�1%<�j�g�G��?4Fi}���]�������C-�Cʀ������Ck�2� �9�²������?����&����� Y���i7Իb���xy�޻k"yOI_m��̀	F�Զ� �a���G�MSsa�2���<��,��}+I��v�۳��2�aV0�?��d8�M��y��F�J�4��5u�����dHf8�yf�){�9��{�;KfҔ >.'y>�]}�d��Gl?���i2��V`J�k���_�q��faJ������"�+�_ҍKr���9$,j���ן�S����x	�+:^{�G�O�#1�����}��Af�Ī^R�n��Y�M*�������Z�`T�F�a-�⽎�d:p�ς��\�P�dB�B(�g��]�Z����F���mG��*��԰��;Q�Ufmp����_J�� �!fs\]%qh�4lp/Dz��.�@ZYy��$�Y�;�[?��9gr^.�ڂ�Ӹ��-�2�~�f�B�\�
X2bI�
�N��uO��#�;\�ew@�]��(� ��RU�?��"8rk��حF�a,��	�S�I2�]�l����?�]`��2��M[�����sh�� X��I9��J�2��`ғIQ���O�����5��){��.�㫤�V\�ͥo
'A���7V�P^�JK�K!!��z(�1�i��I��2`�0��<;��	��0�[�[�S���7Y5���l��}��>��������~9r���4����nR
	C.��f4Nj�q�-Ֆ�k����?/��u�H<A�3G�
����劸�u�d�%����/͛p�U�FY5J��ӓ6��h�e`�~���]��[d����a `r$��l���� �������+���x���Y�5F�A��@���}z���#�]Ç����[��Q}����������8[;|ܰ��J,/G������y߻�EE@���7�;���B���h��2�k���<�t�QQ���� նw��/)z��N�o�mKy[ T�ɦ�Eڿ��.J����m`'���:�-u�a�S�'q>J�o�{@�F��ۚ���?}p��ӬJ<u�X�
�w��ĉ}�vP�Ő���g���q�VW���VX$�HrsF�Z��ْ8^w���N�h�"?ߙ��E��A�������r!Y�mOH�2#7"jam�h<0���b�|£�·4��xe2��-�v�����`�)�� hJ���_��LÇ"�b�Y�f�Z�L{��k/;J-X�D�ZS6fQ
�{�c�$l����d6o��vV_W��w���������G�Q�̢��|xh���%P�ώDKz���g�E����Ɛw|�IoZ��v{�I�m����@�{4�(���+%T�oW?��:�/�G��D���/�S��J��#�ԯ���_��6^�,e9��OuR�7����A�)%��v�B�Bq��I.�������;jX��Г�7G�cB�>��o�R���X�X�:,�/�<'�uqPx$Į�ML����|12�� 곦���<�b��o�q���J�0j�N疧��!���Q�M�䶓I����]���v?ɩ谋�5���"��2l��,�u�8H�ؼ�r�K(�b�G�v��4��Y6�x���m9ڈz�k�l��H��`]�Cra�bkM鲓-
�S���Gf�DK�+Z����J$A4�|��nöB�*��T�����_�T����G����j��Z�f��Nu�%�(�e.�x}�:�8�N[n�77�4xT�:5=�me��hG�ԷK]bS�V)Ɗ�O|D��0(?[21)�I.v)J;��%�t�R���n�M��� �j�=p.����T��?v}����xaG�>֑�7�񘎷\L��p"v����Z�ʏb=�7·��N$��c���͋4�I���y���w��E:�`y�b&%%��d,�cΟ�ځ4��޻������7ɛ��'�rő'�b������Ġe�bu�&��<' F
уx>�ɫ쐊�@�M#�&�M�q�TWt�G��&$W��Z��w���HֱI�$��V@��؜��|u(��.'�$'گ���J�����.͗M�d]>�$J�7���S1.�A�|�W�n�7�oY��0O����O�>v�Td.;A���� W��%�nH);�YY�����9�T �o�
g�2L�6F8;AIe]���T9�l�o%�=t�3�r>3f=���H+�"r��-Bn�D�3��S���l(��M=���g�v�Lr��������������:���u}�4g����X���WjGJ��M��9�H�p�h iP�f���`Y�ٹ\���n�?t�`Apr�Mّ�E�[�η�3(�"�.]��� ��58̙�s/mב<0k��sx�N�4�R�R�;RL�rI���V���
��h�$��T�����>��(e�Mf�����U�@����z�n�R�z�H�}���PS�^�icE!s�$l��j7N`����׬���D�I1sbxl�UY��p�k�f����n23��"��K��B��Z����c?v�x�ˆ��v���]�A&VLVrI�2���q���#CdĂ0�QN�J1>6�4��\������mB�;r�,ef�:�ږ��y�SZe&(&8��.}��׍��=�Xvv˾�+�Bx���Y��Dv�Dja����џ�t�a�Hd�b�Ɯ*��c�>�m+��"n]��TS��z�i�z�H�u�9�Վ���ZRߨѵ�\ev?�l�2�@���SQ �כE�6������v�X����k	!c3�(/�^�`/�`����.ҏN�!�N�ؔ��0U�+��X�QX?k�̂:�����H �!�]���^��b׆�#��0��s+��_���L�e��{�&��+shN�3��2���7F�����s	�>��S�5`�����u��$�������('6u�\�{�%��O�#&�9�k���C��|�͓w����F7:Ҕ�nNK (l��WhL���3�dx�́ќg�w򰯌_�:T�
�Z�k�C���O3�LQ��@-f=cX{����=� Ժ��&Oڄ8��#��W�;-��0D,Y���Ұ��dp����� ��:�?�W7=j%��$!��+Б`0��pc'�<�$t�^�K|�*�u�D3��L�C��"b�!4�q��~@)�@��X�F@U+���ō��UD-J���֥\��z/ZI�dvb|��V6��KT*H�O���ܦE���^C�+�Mo+�2ͧ�S�pW����� �5/�1=�O�h��W�r���43��5��������� ��(Q*���=��7x��K]x��f<��9���}�|ډ`����2��v�S���\@_�e��df*�.�f�"fҲ�kʁK�c���8���E�9K���)��wF��SHg�K�x�k\㰩T���߱@�ɵZ�1m��8W=$$�k�o��3,�B��Sם6=��O��̦���cC~%��c�-�/�J�ٺ�R֜�z���׸W�.���%hE���fo:��L�Ɖ���W��?��`Gm$��(�-h��ʉ@ͯ_e2���
�߸�v�-��e/ zi�L�����a����?�:�H)����o	�D��r7���%9$�~����8Hz�U"%��*,���6�?/���A&�U�}~T�<#(88.�8mqPjCr�b;N�z�D�� �M��sΫ���P�����\��f��(I�/�V�d���$�M�'�2d°;���%�Grnkx�ߏ�k�e-��L̫C���#�(}=���li��ed�m�@lhL�����W�!�Jʎ�gͮ�����j�����e� ����	lU�Q����ҵ^ӎ��-�0�[O�(m���B��U��V����)����Z�<�#ړ�R�ɍ�&�� 0����L�iƸ7���9��̈Q��j)�q�8a�ȗ�0I+���� ��5q�2E�A�H�>Z��}J[[ۅEG�9�vsp��D�t!qoI�[]ll�U������1�ύ��
vȮ����W'Ͽ� �2B����y4�L�z���3I���5Q<�Fp<Oe7��+�Q�1c��y8=r��9e\�b�ɥ���Z�z����5A�`�{!�S�s !ER�מkj�Å������*���n�H�o�8�P;��U1�^�L�x�PaR��6O� �4[�0!�槥i(�蕖q�����$\hg�'��ǒk�F�����\��#hv��d&�6H��ݾXj��<g�c�[xHD�%6�*��`���$�� �-���ֳ>�Ȧ�%5q:���2���!OQ,�fX��)�K��n^KZަ���8��ܔJ�=ȃ�,�-fK+�acc�"V��v��6UZ��֖{������`�����O�����p &�+�|�k0Ƞ;�&i༳�q2�Vf��p9��� ���I���H��4��(�Df���+1�Јm�%��|c?��:P5�wNP���ب��}LY��a^��]0�q��y`�Z@J�&�!Pj���YH�V�	�W�b\h͔�5��� ?�֮�n�!�p-=�ߵw�}���Z��?k���A���f_��yH`�G�����)�� (J�r��]a'�(,�c�K^���&�ȕo�_m[�j�n���z����]&���q��p3��U(4̐z�1*�. �K����g2̊Ge�s![�-�Et�j�M܍��H��Ox���;��:��E��1&��Ӕ;^KF(#~#�5�� ��i�u��m��)-Z�Hw@bl7�݅_�wx�WM1�IE^�2�0+g�~`{c�>���<X�H�ǔ���mĘ+8S	��?�{NuҞu,�A�ȲE�
i�% ��9^[X��x��i�k�q�J��w�?��g`�X�ĺ! �h6�,ylܠ�?D�l�����LNUx;S��T�����]�r��Y�N����F<2�+��� �_�8��0���g�~�9��T��c`�{Q����B���f�>���&��Q�ڿ����K�e�2�ĳ�B������t.lD��dZ@Q�v�@:��{�7A�>-hc('����d����Dz([��D�c�ۜ��������+���6;`�1�|n��{Z&� ��״��j?�yM~j���5������zp�G����Ե���G�5&vv�É	F�<�����oȥ!�~�}��䗭�J��(�܉��mp鈬Om�
`۪1b�A.�$[dA��y�",D4�8Y��Q7�1h�`|���s��'�t����*�����X NXiAP����] �p��$�z�C��{�E�hU �%m=a�+�������*�D�#8-�"��@b�<��è�>I�ITz��*��Y
���]}�-���]H��y�)��"`��Zm�`�)����s�2cmz��N����ؒ5�J�����:=�"�Ui�pr����+C>S�H��!bzA �T�MZ�k\4�R4�� en�� ���~��1��C��U�cG�m�>��S����'���$ߣE�E%�X�G�K�����7B0J6��9C'g,4Bp���*��|�g�Zm8%1 6������*C���]~1���;n�c��O�
�%��w�~��8�:'�j2)F�6�7�v�>���t�A��c��R"�V0��dY�Ȝ""�܃�1��\ ��W�4��d��䥁,��_б��=zA񽬠"u$�/\0C�K���S�,[���S^����h�Ӟ�+�O�ws���#��Dp�wٻ!Tgg^Sw���~�x
+m�e-��ʓ���	����k��?7�v�*n�7Tz�^����~�K��?R�3��6k�Ƶ�5�#X���5�)�Z*ř�s�ВBX�3fRR�5��G�K_E��׀���>�J:�;K|����J~��(v�3#�g$F:�2�p�X'�/}$�xuư��a�*�,�ڞQ�X5b����Οgh��ē��������a��8�.����'�1�A
g�Z��c��<�O�7���%<�Q�r"�����~�<�«�]u��SN���a�:,�Y��X*��\
;?��3�.����37���Ж0O3Lea�3�+O��X��]�<u�O3�1肈A�������@�_VL[�힓��KZ߰��-�m��*�8��Cd���^%`���~wR��SYJR�K`�)�|m
*��V
�ޗ�O {r����c�#�5jO�tn��Uf��j�$�s<\3Y�p���<��H��u�b0҉�]}IN�����e���j�酱*9���A_f�sk G��F�vz�5m�rW�E�b�F{v}��'��������2t������b�-A�0Ӱ���5t�A�6����+Iԣ�4�h5֔R!���*�/ߎ��e�Y.��6ZU��=�a�Ar�'M[,m�,�S2���K��%��(�k��z�3�&�p���`�y�sA�	O��t?������ٗ��7����@��7��g�X�e,��,
X���}�3�yKdl�� �%��P�&K�[�kb�|<!Nȿ�Ơ������tkl1I��+?DD)a�2���)\��!�5���f������C�_��T�
J`
��p|�-n�,:��2��5��1�Pg���P.���q���"f<��|��bf�oۆ͖j'���la�H"H�B��Y��*���P}�4s��XVj�@f��A���^1��ѥ�u�g����b&*W
�9��e�0��#�ש����4{7�C���A���1�w��WÃ��l���P���lp�Q�S�)O+x�?�J���3�����lK�>�Z�-�٢�϶�����5t``L�_Ȇv�;�Ԑ�AL��<�Z��0r]�<j�a��՞I���v�Ǻ�^]#�{*$�;v���$)����6���ؤ�`y��o?�H*l��)=��]�L)C�a��y����A~�Io*��X�D1L�x���u�C�J{vL&K��w�C+n��љx��"Q�Hq�-�c(�8"��xE��^c��}��[hkJ����H&��B-,ܫ�L����0� �41��Dt\V��kG�����1�t��K?�!�Xn�kS���u��eV��6�xYR��N��˜f,�)K��磐*�Y9��[1���+hQW��}!�+��(*�'��al:	nU�b��7�������k��W����k��Z����������M��u뱵�0AB:ޛw����ZC' �O��+xf	h�w#�v;3���Vm�y �A�����?J�*%�!V]PS���ts���N�)�	�:����Ũ���K���b����g�~��W����kc��٢cN�Ĳ��-A��؎,zЭm+�̺���\�(��ߝ�9O��&�1��ݿ�&KH�8yXLP�j**)�2��f�^*�|�h_)Q� }��N���N$��zq,�߯U�kv�XO�v��.��z�4��Ғ��y?�A�"�?�����M�v�ͳLJ���~��UK [m8�,�=	�).'I���l���ĕD["���A��L��ߪq��~&���HT�;�@)��#���_'-��,砇t����?�uL~��䢩u�>8 9=�:+���R���E~Kf_p���dj�h�Z$L��b��9��O�TAf���wHYN����e�a�)�����Dn���j�VF�1�C)^���3���l,�nwfШ�Stf�F��alշ9g����|9���U��A�ؖ�&O����ka�"4=1X��J%2�X�� d���=k{;vw@	��-.�c�ˌ�!C�B1��#������KWg)T.0<�v�N�[e+���'ڈy�a�sF�m
�� '�p�aY��s#Z?����_goc�+��`J��®�1K�]��N��d��~dᒃNv�t�!��m���Y������C��`�\a)A�.T�U�I͆�
�n0�S����>?a���"�Ly ��jLa*\�>�Ĳ�6"S���N4�L��w���/�WPgǻF
QӲa�`�D�4�?�s�v�g����%���|J]��eZ�S�3eci��S��h-�Z�ʪ���#f����et�*
g���9����l����(ݺ��6��BGӖ�@�	�
�g�F5�вe*��ltWN�3�����g��X�	+�e��E�ቨ�i�f�bZ��nKT>�����mK���YT�tg偩��g�#�)���d��"_��N���L�A�0�}��6JxA�͝*J��*�% ���:�b4�9�K�g/�pM
�gѕ�t�\����biP~o�e��g��� Bڐ�-��JwϦ7���n��R�ǔDM�6�!��u]������t^R���i��5�?f��η=�77�t��`�z��|Z��YR��`����(���E�T^��v�~1,��E�j�1���U���u�_��� �.5hV+k�ӭ�xV�5�O��,�^A�p�G�C�����0n���'�D0�R�G-����@�]2�����ԍ�Ɣ*H�9\�b��Z��QT�:�J1�wv�r�w'����v8�j��~�	��Aqqk;�m�^������/�Ŗ���xR�ط��M~|G�'�{[�l7���c�>��=�%�ݞ&T��D�ۗF�t{�5�S' h�XZ�\�!�b��"�`}����0uC6Z��UG���aw��,�ӫ@!���=�u0'�W�^[�֥�����ʌ$B�].UJ4vqL.R�hQ3����w�6�iSe"����u�֫�����1A������	L��|eO�X��#����{��Lb![9�&2��� ;n��7/�35U"��ş?��h��M+�@�	����N��V+��4(Ȳ
�4�lS��KQ�jX�ȂS� ��pc�P�SYnHgR:(��+N�m�L�k��h.ڴ^����.�sE<F[du�g����c�Bj2#�� ����>�E��f��jM��l.�Y�1{rW4�\���"c+�����VAwo�~9�i߄��!�I��v�ki�kn;c)� �/�.[�����`����O�P-�j֠��	��s���[!�����J����F&4�Dd� �� �q��{萝���<�� ����86���u�|!Mp��%�y.�/0�	a�=�)�Ȳ
���K��kվȑ+O	A�7F��~ǽ�؀��?��[Z^"j(��4�MEP�3u�]ʎ��Q㽀���J~ІAF��ht�VТZV���� �օd�F�恩6�*�1>C������=�&�H�G(.hhP	�ŭ� rxQh<V�bFO�⻭��հ�LB�*ˍ�>�i��=�^BF�R3��&�#�{σ�u��|�B&{�"𜏽���{�v�0�P[�qG�8#�3����+}�<+� )���2ewjۯ�G�(!Ɠo[mo6���z�yD�`D��o��ܮ���d�����i4ǷV4������D�6�5��={�v��W+�9c�]��Ka���R��i)<�@�OBkk���ޖ?u�o"����L�8�}���R(�cD�e�]a����QQ����&��8���-U�׳��:���^�>�����_����Z]|�0��CĖ�p��+}:��7���S켍�0-N+@��� �<�;@�����7ǐ�ˉ�i�G��Wꈜ��mft��������d�8��r�?б�)|���f�ȶĂG�����:�<A��T�J���&�5�z�?��Fg���FP�,G�Af���d��{ZǕ�S.�I�>_o�+ڃ�(0����3�-iħx�����z��B��f
K0"b���%U8AJ�����r$
�8�q67��'��6x��<Yaq�ǡ4�Z �k\C�B�+��`�Q�i�\�
йW?�z#?�C���2�~�s:��*I�/��z#Z��TY�DX����F��~��>8�,]yÅ�H�'�{>QXx��J�j&+���)(�쭼?��%�X0�=���*��`�>����h���BT!S��e_�����[���-a A����
&3	5�s��^l���8��uA�$R�܉/�N�Fy���a�mi�J4n�R�YPfA`��EDݖ֪��³���}���LP��#1�9�9�i#;tP��ہ[�����`2�@C`���<>���mc)�����)8��7h�M��q���@��Szp,�v`�t��X>�k��'�k�Sl
m��s�Jq�d��੒eۭ�=qn���yi�Iz=��Ϧ�q�Z?^���O�;K�媷�V.��ǈK��<�AE�k롍�I��B�9�ʬ�y� ܣ�%�P�M�#�a<"B@�>�9��%υ���w99E�T��!i��R���#��f���_'pE���ȡ�e�JU�[uU�"�L�~��b�(֐牣s��)����HPj�!p�r�-�
�(a�
z�̎!8݈*(�କZ�� y�g��U��x!8�b����6��D�+�Gjj�p�H��5�h�4������V��Q�i=<�w�d�K��E�ܹL��k��V��y(G�/n�������R�qp��[����ֵ�X��Bb��/����� R���/�C*��Jj� �hU��w�%��F���
�5;3��RR�Jo���A�MN����q6�x2�l�Nh):F<�1YKˀ��8��2JI�O�;(��)�N,(�M	od�H�wD�W���(u���A�s	�p���¸�ۼ�v��*�l�ɭw
�1h��i��� 
����,:�FRQ�+Ⱥ���ZE��4�!W�o9fN�����@�u�\m+�)e�}��h2��N7_�̌����o&3��6�������2�q�����oPG�g�~����7�hr��ܱ>N�]��,�op�]b���=�MڡZ���i~�p�$Io��E#?��s6xQ�$*F'���0hM$ ���C��gw^[ޓ�ĿL�է���{��ť�Q�2�*��2h��L~[+z�Qgok�K��	*�&:۲�E6��:`����6
���:/_ }�����#ʺ�8k���?r��tG����b/�y�9a ��������!��Tr�X���/��(~��O��@ᕌ>��E�;��3.r��A��Y���7��E�r3z:)���y*�|�H�5�{��T�㛻]_u�����Y$iD��>�]�o՘�4Z�������L��l�K�r"_��_�gK�������?x���
~���� ��h�d������@�䠓�sS���F�,��Y�GG���Eux^Қ����;�gi?4�v��Aȗ�{9����8�7!���p���9n�����|~W7��2oO��F]N���\��v��E�#�N1��tc�1`[��!�R.�Hď0q���9TI����2e#F$4�F8,u��ʙk����R�կx֥iY��Ґ$HP+�6����s�|d����ߣ�T����g�O�<PX��Vh�Km����?�3j�E��v�z����dLU%������x�Ne��+��AF�l�gAKU��ĉk�cqY���B@4�>�g~���)�~�tx$�,�8��ϖZt��n�d��V���a��Y/2���c�x����\�B�?-����4�1or�'����Wk70����[x��D�T��* 7y�=D.�����R5�1�۴*�\_�Yo7Zᥬ`�V)�֕b�P^޺���#�&��	ۉڸ�XX+DR��2P�ʲ�Xc�+�i��]�Tq�kv�o�
(Խi�Y���*Iנ��XO��\�<��T��3t�S�V~�kƎ��DI�����<�x��[TuZ�Y���F�i_0�;�)a���q�`N��~�L6u�輶�����A� ����v��RQx<س ��gd�h�Qa�z��G��]8F$���5s��$��p�.��Ĥ���*�_�~�������� ��թ@��
^&�Œ���M'�E�c��UC�VH��to��C�ĵ,�����k�1g0fQ� "s���B; ���{%g��J$�	!���:a:�̠�rDOZ�4 k1����f�V�_�屉Ք���vO�S~��V�2�C�Wc��d>d�B�0��$��:9A�Zx Ӡj(��\�m�)ẗ́w����ڳO�n�/Aهaf��({���zn*��`�� *�t�Z;�K�V[@���*�U��[��RO���B�"^(�M�3qmƘQ�٭�����lo��oڍ����Lҩ���-�:l_Y�ll�rw�y��eo��H�2H�|E4�H7]��.핕^!�^M���eշ��w���[����m�ԉR��j�H����7��j�3��@���A��L�IA�\C�3q��k��8L�,�7jimw�3	K�p'"�[���{\��VI�xq^)aoZ�*��%a�wn<�{Eh������xN�J�0Qn��(���_� ���lo
"�n��U9&��~�oP��H��f��)MI�ha�� 9�����U	i��I5��a?��|W,N��{'�4ↁPb�6����òJ��T�Q�=����2Hc�|�����*���ڑj�"5�,�Z|����#��r��0�&��類��9G�֢��F��U�ˀ������꣛:fהy�V�"0�M&]�aN�Bق G��&K��	k陰�x���7B.p~�b�lF���Qr�F�4�9,�T�gDc��X��7#�\��ӯ�n��-PJ_g�L����`���̂��-��8�%��s�7T�9�P��<m���_|m�U	�P�#b�^�K�lj�6E����Y�)�M`8{WqPj\./V*n��-�r�´�{ޜ���ߺ�py��ŹM+�(=G%���`�縡kE�P�Ҵ9���
�E���ɴ"�ٽ���"�I���p�g�'��7<)��B�Xb����������Wx�vh��h���sDW�#~���`��ԍQ���w��y��֧0˸:Z��]�H�XE�K������Kԯ���-E|�#�\�H�[�.*�T]�㜅\Ca��=�U�W�cR �@��+��	�9��w��u�$^֚���)G����Sm���n�D)[�$�XsK"Д�I��4��ͅZ��E�δ��wP���r���e؜l��)��l���n�X��A,(0]�)�[U�NS	M��f���:Ў7*r�N�߃�d�ٸ��6\�CC�I|b�7�ߏZ�m���|(]6zN�(�v���(��XՋh~��9>�|�BɐX�����k1��Ÿ�9�=US�/�i?�rT�v�U�$u�k��ӈ���3y��ԗ��[):� Qv�zD���	mD~���$��-�1�@�<�(Y4�I��?s������Ҧ'��q��4H�)�.P����O�#�/�X�;��X&��k�b��qQGUHc��Њ����A>ޥi]^�*�������)�~����qT��؂��^L�:a��3�gΜ �R�ьj\w��0�2/�:�ڛ�D������γ|��F��Ѫ` ���֙�&�a����lM����ރ{焃�����j�D�ج���:ON�KJymb��G]Q����K����BR�]��L'�2�����IIg����'���f��iax}��s&a*���!�[��9����]�'w��Z��b=k����oY�qz����o��q�؈9���ú�����!ѰQ�]�Ƒ
"Ca�������d���ڪiC�j9_����B�p��Xv���=Z2�zo�?�����}Dǳ�/�j��NPb�#xr$bi��:.]�To� ��p��I]W ;�z=������ĊF��I7hrC�r܇xh��!�f�#X�vf����O�}\s��=�u��]�H�ώ�@�z�]Ñ�lUЈ_�kG�$��>F"��o=���D�˾�̓A��~S�Q�\c�ѓQ�(�jC�
���R�-u_2CN�AKH�by� Q�2�Z����H�꜎�\�J�9������|��ƴ.C�ɫc����(�z3��Si��v����KFt���V���Q�t��v���.|Vtڦ�	[8��k2�f�q��F|[��߻`d��%Xg���Kx_4s�:3_�_�v(d�|��;����rp����\��R�AeK8������+7�H� �������� ^e�	�m��E��VԎ��/��y�V>3�b���X�hi=̮o�G�>�	kU:X�$Q8�B���NϘb=�Z�&��x\��)1���
G�d&���0��斱k�'幚"u�Kxʜ���v�m7�Mr������oZj��:�ɤ����T�6�֌�zL�C��Nt�C/:C�@�P(>��.�M޹�����~�͏Rx���6���Q��.$�Z3d����Δ�&��nj?����.��c0�6s��<��.�=8�j��9Q�{�@V����.���8ji��%6��$���3�U09O^s���Ir5��7g�":ڕs�A��[-�:�4�3�q(ۿj�M�1®��zV*U�hY����z�Uk����S�Tk����#�p2R9+&V��g4Y~�@�Fe����g�����o��R�1F�N�VRyQ;ߴ�묢����:��(_t�����v�N�,����RL��$���O�|�;�˺�J�C��n�p���M���8��P�4�'���h��ۤ�/n�	��?\�2n��_9�H���96؈L�"8?���s|�z�<ݠ�\�zWh|[�h
�R�n
�	��.�V�m���qț0��6�Gs٠�m�a�u�������RT��л�/}�eG!��/"���L���V�-'���0y���h��AQx}����N(�<���S��ڳ6r2&�����&b�^1ǝt5�Q b��wS)U`���甑iI�+Ǧ��*e�W�rKJ�Zrt��9��Tq`uxU�O+�
��3��O�z�b��|qFm�6��E���\�O)����n�L��)4��s��U�;e��!�,�x�����/�����P2sZ��� \ף�X����@Y��Ɏ"`�G�:@K=�>Uɗ�������BD���`�&�	�(��/l����<�>z��',���h�'A�: ۸� �7�KO�>��Q�Z�5�b�Y�S��#���Q��]�u�K��L%=��j�-�CѦ}B��j��x�W$��"FcI�٬ͭ׃]&�w�\�ޒ"l�d13����Pa��/�� �>�.�����ZO_E�Vcz)�nF��?�.�"�؊<`�?�b/�ec^[�����i���4D���ѷV�Л�����jL���,1N�9��mCq��2�w ��jO�{w]Y7	�^�f
���n�zdOd.��0WC���|�ͥ�o0�_Z�&�aH��LׄjZu��e��}�A{�4ꓲ���k������$��fV�.ZCHJ���`Q��$;/��.d���LE3���}ШI��f��WJD��sLN�Yv�odt|D��ǻ45u�t%�+�l��P�^��ZL��_���CK]�o׏&��ng�vP�h�L���B���Tk�����p��Az��#� c�>��7'��
�[�	fu_g�ꡏы9}nd�!�m!_P��!\�H}�Q7;�w�[	��K�Q䅿�c����h�^ޱFl�?} 6�kg��$��z�nO+2+�$�P�#��T�5��ɠܰ����C{(�(��4\e�O��ٌ�1p����1ĳ��~�g����J�sO|�n�y��; 3�c���L6SR*B��и�;R~����b¾�^�^��=�����x�BU2f�z)_���g��L�z=E+f����O@��ƛ�D�C���BM�zKTEU�(���@��QlK�[ɍ
9��R�:�ʲ�qnZ��6s�u]��m�scb")�����2�mo7�ץc8��K:�{>�9���H(���w��#4�������鸭��b+�
������̆��ol���Sľ�����z.���2"��0��Zj$
��c
���!�&��1볿.	�L#���w��n�/�����(��*��1���Jʞ�M~�W Z,�f/���kpϺñ��r���+|g/Gc9եI		YO�1��g�W�q:(��a��up��Դ�ou-�W
�2�Օ��h݈���9�>��$#���������n���"dQl���MO���ζp$[93��f�v.����`
e�>�L��N�����E�����������]%0﬊��3�����j( �	v:�,�a���G�����I��B'>�h Tά�����*�(�y��=����H��x�0�V�A�+~Y�{�N���ӿE�
ܷ:��T�g�����;�2�~T-L�%,lb݌C�Z����`0���F��.����zF����E牻�a��ɻ}�>:����h-<�(��m5�f��gז^����j%�ҏ�j��@�Y�:c�v��#���0�
+�	��kT�`�8�|Ű�N�sV�`O�0�Q��i�3�N�_��gn�ݎuz����G	o�e�<��/l�L���Y�ōn��{gv��T!壇����g,�jus?������G*���fUȁ�����|��ŊIs���2N����
@�y݀
�Ȥh��O|d�9�b�:$��ۻ3�m9v�!}̕���6�s�  ������S.0O�ɹ�,���7��|I�`����U�QQ�i�z�4�-��T/x42tk�%�?�h�]*4E��T��'p��k��'!�V]�F���̧Occ��n��#h��W��A�i��R����/��X��4#�H�I�jf�J��U��6����YZ�I-��s?�C���޽��=�q<�w1ᝐ�������cڮ��S�z����i(�(k��@����υ&(�+���9�8OK{Lq�<��K������JԄ���dfI��/�� ��R��H(w�s��z��(�7za�o;��Ù��`�z(�3N�dl{����m�"{̼�h�Z�X+�_�]V����ҙ��qew,���{G.�I�K�ǎ�N�x����wh��_[U�l�w2��b��"51�V��n�ǿ�]�����8*��~-�P�S��V��"R�q� }HpEi .�����/��T/�H�1\���xщΗ6Fv�j�G���B�vhB�4�~
u�����n��mS�!��}I��u���Y�pښRR�-���p�*�ˑ�-��%��t�3<��C,�gf:!%��Y]�ne�pa1�O��C{'!��ʓ�=�BL��'"���!�n}:�`�O��������'|a[r�f���hA�^)/d
�T/�e��Ԇ�W3�@�LuE��"�����k�5Y<�K��t�+�/���2��6�G�NUp4�uAY����&����=䢻ZL[l�V5�O7��S�*�T@��]D�X�C�y
aF�8��;�Z5,&��s�r��|uG���S��G�?m��(���EZ����9C�I�G6j���0�wk�o��9i��ՠ���=�}��G�O�'�r�z ����N��Ł�UR0`����½��{�3�b_8����$�ݞ�e�w����(Rq_�Ж��e� �t��u�ӵ(�B�o�?SV>Hx��x5�{��v�.��#��枱i.���[~�x���2��`�j6q)�#�^v��q_��06ޚ�cT�Yĵ<p�����'�]z��j4[���#8	�~���! �/}B3��ܶ�TK�U��^����ީ)e�Mc��
����Abb�f���a�kQ���2��Y����6]k���?��$Vb=}�T���xOer(�%'	�r���ϭ� �����߇q��'<5ݰD����I��D����[W<���UIW~F[��.�頲���-�f3{�u���Ez:J,���}�A�@�����t.a�_�ڑC�˖�y�>�g��@�K���W�a4���u�l���4��=rs�4�N���B��r�B"�k���*=��g�hjt%��0��=���zF�i�v���ZS��L��F������c�0�RV��D2(Q6��Z	�M��?��X5�*��uyG�c�\4��#��X���{Gpf�<9� ��8�UI��4Q"��n�k�^�o�!��g�����8$����ժ���R����rl��'��g�VNǤ�����s��M$tAq�,����R���+�ti�}���������h1L�����v�Cb��b�-�@�.�x�@�:qC2��s���D���Ӈ��py1f�zL۱��n�(\�x5�x3�4��?�5�	��1,#���ح``������K �O�m���ګ�}�u)�����'�L�Ƈ�8/9�5����pHO�І�*J=G�Vc�i|bW*�o{�'w�!��}�{]nJ�`]��~�!��ئ�&5F���6:�����V4?�5�5�������Wv�ذ���H��q`�ֱ��:4�aJ��[��0 �7K�J���[��bE��N��m�&�ߦ�$���� �ǋy�/S��
�<ih���87�ڰƫV��nS�ɞ�y�tϔ��H��]�tJ�w��#��Q�qYΟ�>7�֞�E[}�}���bQ�T��p���AF5X>8I��o�,�H���9*���3�����{íLb�7�fS�?����$q��>L�����E����m����ͣ���������l<���s4Z2�ج��[꿒$�����2/�9���	��ΐ��{��h�3l� '
�����x��_V��Ɩ�0"��m�QѨ|������c	ӭ3x��6�j�%�,^g�����5R����"�' "0� ���&Ǻ�(����[|�tm����8G�����`���1	�>
[h��O�󽫢��f���&{=�1�B[w5��'�6���d�`�ֿ��I��ek08�̿�-Rf��JA�`�T��� ��O]Y�m��*��R�A� �S=V�\���y"D����ͭΒ�ʆV�����%/���!��^Z�"�&\�n]���`VT_�
{�E =(P��ţ�ů�[�$��,�'Y�G�r�Ψ��[�����M�a�a���ȏe��}&>΋���=��!`�y3Ç ǅ�i1UgD>~%=�Q0�� ����w�W��"�/�^�}���p%���y���ϙ�$7/���V�����	��kͧ+"A�,�k=Ê��*��W���l2�)���up�v�D[&r�~�a�\�v��7µJ\��u�z���g�v<�IYˌ������2ѣe���z��oF�[����ku�{�^�l �1x\��e��������	� ���~�,q_���Q��|h�GҎ#�GOU�� ��v�F��b�Azn�t!�((�c����Ï��A�_rh�۾"(���sr�|Vl)� l(�I�m�t�4"v�a����/���/�HL��[����Cᐡ���-�|�dp���c��>�W�&8��"
Q��գD^[� �lИN3ǟ`�t�GrjWa߆���/���g������ nz6#""Y�@��RQő��hq�����`��^-����Z���^�LǸ�PU��fg�����I��/*,G�0Ul�	v|�ش��#X�����[�=�F{�c�&}�\�fuG	��)�W�!�_pO�?�����i�X���%����������{��5e�u�/�	��|�V^+��)�����	�&Hw���;�d��!uJ�������S����7`d�S����x�0 Qr��g� ���\X�z`�`�~��y���s��$�^��R?Z <�Y�<�f��p��a��0�ƥr]��e���諍��Ds��N~X���4/ O#�T��S']lg���K�2#�0!]�|�ᩕy�<*y8����
�?U�N�/��$=��u�g���-5ZOZ�?����\�����@�sr0��'�߇ms3�0߷�0���yQ�{W�"ױ^����, �C�(6�uq����!�~�I\멄��8��*L��Zh�h΂&�2���MF�M䢣��	�v�~}�	�)�4����y�](��葦,�s�*�q�)T\�k�w�/�~Xز!��虥�<�=�*_C�B�Ũ����y��̔�;��/;�'�{�P:�]r��"F�Z���͂o�,��F������Q4y��Z�P���=���,���	S��t��ۥESJ��z�|�M��~�~�E9��dI:/�8M)7����
~z��QC� �Q�`�{`H�վ�o���Y�^��������^�Bq��r$���؄2#�k����<u�JV�9X&�� ����kf	��q��$/���*��.�����SV��?b}�?�M���݌�򀷫��(Q�55�bT�m�\��l]>�(�p8�X���4z���Bv��8��{C��5��N��r�����ƒٴ>����B��N��Z�+�сy����vi!.K�k�ҽ�W]��p����/��,\$�ũ5�o�<�:��b
}��֜jA�"x��~HQR�V�8)|�|$��Bv��d;�`���m*�-X�YQ�8��+�ғB�@ɹP�o�6�;�m��Q!����r�4�S��I��P���C�|��qZ~�-�i��e$S/'�e6^��vK}�_���������-%0&'KŖ�碜:o����#/���)*7�3b9�i�����2 �O�\�&�1	�x�z�7���{��Ï�ޢZ��PT�UT���N�[A-�.{�ł��x�Vtb`u��t�*3��ms��k��J?%��Z
x�قH����Q*ѽ��$�t�$kj�8c�:[pc�� ���Q����[�N*"8h\!4\�-�*/�-��%�HFFC��������-n[2V-T��	�H����O�\/2���i�vlq�q�}�x^�;���Y�~�Ӹ�3-�C����=������l���A�fR��UD�xٖY�ֿ�îuw�F\����=v�	f�К鶨
11���h�\��y���ou�I�Z;,w� �\
>L�k���Z����l�������!(��h�Y���ũQ��ʧ+p�)SN�1-��*��j%�m^��g:�џ�0�?]������s��Л-�k
B��I��G��-r�L�(.t�I9&ERU��*���z���SK�=����N-F�8�������&�X[�GsE?/�HQɘ�U�8������s���;��=�ŮP����M��̎N��Gj], ��L���_"5��f� VV�|�h�Hh-/���?���\x_O��М�LC��y��� �Ʊ+�:�l�Z�e�����*���W�<��PwɁ��$Qw���cG���L� H����(�����0\��*��
�Q����ڻ�[3�`l��6��4
Q��(KS�cZw9�<v�Ed�e�
�Gh.�`M#��r��0V.���=�w�U1�nQ�s��{�>��Ϗ��$�g9U���=o�0���Bv�ү}��*�c@X��;� #�cQ��l�)����*��� γ0@�x�gS��[T@��9U��	��v/?�zS����'N��k�p?�驙8l9Wc!���*�2��H=5e���F
��'jV �g��.a�PwǙl���_O��]<��3�LD;ȼPд ���"E��4��N'���kEh�F�����,�t���1��X7�Ѯ˧환������J$�7p�$Ơ �p;&ቀ}�;$���<��\���IH94��d�*�s��}���^�������p� �ҭa6��n~�Ae7���v�����:"�c�;kd"��1�������m6�a�@6�g�jo�p��I%u�\�#Q�X�Ȇ���,3 8��R�O�v�j��!lP�ƽq��B�_l`��r�kPdX):A�X��y���=�������奁(����̸ꄶ������PCL�z�d;�^g�[�/���J���z4p��_Cg�G��.�qi�����Ƭ5���#�v�1�� ��v���/�Q�ܗjCƪ:�_�<iåJR5p��A��!@�n㘱�I
~l4���yh���1������bV3z���Rs��i��0/���P�$�p1Y��I���bP����X[l����)
޸[L[J�ZƗ޾��f�bQ���藗��T��u2܆>0��ta"ݕ7��������rI@�N�Q3K.�t�ξ�OT<����K�B��rK�a� ʋ�ħϔ0���iґ|-��m0�'���8�u�{�0����K��x��֎��Ć��ۡB(�5Y�|��4\fk1N�aF�o�:]?�Vg2����Y���P�A��&���;����^�	�Q��h]_��}'J򛇓NH6�Lߣ�+q�Z��xC�r�Xۘv+Nc1��:���A6��J�U`\�`�&n�>O��_b+�F���f��A3?��K���i;˔a�&POl�'�܈�MSl�B{�9	�b)V�!LC�3o�Ww°!�#��O+a�۰zQ�;&ٰ
�ú�
B���6��c���h���?�h����S'6׹����̐���+f���W~�ZG{�y���N0���H���`>�����^|�KQf�|��0��g�Ws�3���m�H����H,5j���@z��4��!���k���68�}���1H�x��`�����d�7��0:-�.�Ot�jd)~��DY�M)C�����2�e�:�9���&�w�	�K˚��ߟ��j�T�zl�yT�z:��䌡��E?M���J�Ŵ�G�*�G>r��p�I��OC?�Ε�k��Z���	rB ��*�MC�Z����B��YC)�*�^aJ�⌸y^"r��-w�D�-m����<B�$�|2�pC���)�{BDIEKy�Q��;�������D�~�R��˪H�qߺ f����N�[����)��p�]�>�ڴ>,���_�4C"F��Ip��\�i�K��\�Y�1rJ��M�F �b����8q8݁5���>��U�X������>_8Mɖ�%%o��d�|��X9��7MbA'o�_^į���I�<тO}$RD���iP��֯m� p��\�P�g:K~���2�l:@��S����F�.�s̩�y�_�T�
t_�6���~O�W/�-�5b����c��e��u�3/%����y�r�_�G�IP�q&��.�D|�v�P@����^^l�M����|Y;3���7�6�ZY���/�����-�t�m�+IN��� Ƣb����N��ћ��/ڳ�EZw��9?(��HӣNIgy��مoQ�.(l�����g
,�j;J��qJ����l�s\8|������!A��:��}X���-�~%�"g��n�	���2��
5ߧL d���թ�a�E-.<.����Z�Pc��� �d(rJ��,n��b
	�"SՓz�����*+�]���ut9C�Y	���h,��E��x�M�s�٦�-3�*Χ��l�b=�D�\9�7��DD�R�^���NOr޳3ޡ_.�����c���T+.R#�?�%� ߡ�{C#�g��ʍ:jx�����-մ�@S��D�Ϩ���D{_xB$�� ���P"0�zP]c~.+�x�i�G�Ϸk��x�A�GXC��R��,�-��c��J���K8f#a����5�d}?L���z�nGp��g䕬@(�7y����3�������Bn���䡹�!�Ш�a��C����~=��V�Ɵn�i�	!|��C�&_q老yp2��4�S���Wʓ����E����8��m���K�}&�p�-����GE��-��(3D-�S{�F��vc��_G�3�f���<a+�����T/JH�\_>l�H"�i+ `���*��u���$s�E��+�87-�ˆ�x���m��=�ֶ�k��6�Z�T=B���9Qt���i=֑��F��[�6�K�*��7c��CL�1)]�<W�$N�������_��a�ZxU������~b��>��z��	M9g �{Mp�Z֠����� Aߘ[���)�����wcF�����p�H����p�B%q5l.gZ�+^�Őp�/���Q|"�)��������(�"�L�|c!I�^9o������3�>�C���ˑ*sr�c#��Ӈid}}�D7:<�9rZZ��x�k��}q�+��5������sVPI��~^s��C��^"�OU�sOU���A'�Hm�L�)�_��C��~�Q�tP?2��4��dU�bc��{ؕ�+���Z(���V"��D������Rn�/�����n5����l$�3t-��\$��]Iq52Vn� ���e�!�]͛��8wa`	��B��H���ʛfeU.��ݖv����e�TxJ�ӽ~v�P�؊.�}흹�`O�O�����0j_�^g��㕪��Q��K]�C�<;���s�ږ컚���(|�/a���}��	�ri�}h���${�s5��<׺s�"�Eq��5G�B�Ʊ�!Ξ�{B�[	���YK��]'��$=<Z��D�U�u*��'�ѻw͑�S���J�^�� ��66�C�XS�|l�.훻��&0.Y����odچ�N/����r��
����fhr�U��||�X�e�Յ�R��3Yb��s�A⾉`�+��Şp�{��aZ�3��^��8p�b���{������W���$�5�@�/0f�o��p_�:%>"�7b���h\�0 W{tl���}M�(��{ݔT��p��rjI��0h��o����-@�-����r1�ݢ�2Z�i�1�����`��;B8��p�����YW]o?r��N�|�oW�Tڬ*2��H�l�y��m:�"ԫ'���=vv��HW��'�Uf��Yp��gg`OQs�
]c���QOӪ�����e�}�XO��c��eNŢ��^���C���9��H����Gy�����B+5`����[X���~p0�T�z�fG��iKk�QX�*�����2X �G`�tȭ�A��s=�PpO
x�3�/�<U�$��=x,��p���G�s�|�߇̕su���v~7�i�~x�I��7�-���ZX�`��%>�3A���@��G��]�`�����s�/��sI�0�'l?��x/�f��6��<n-�����V�6��Ѧ?߹��L���W���R��}j��:L�S�6,/� ���񓊢�,_��E��dN^��+��>ܩ6����Ю� �q���\�MR�~���F��K���v>c#j�~����:��u寺 �+ *�ޯ��3�(nE�cBOf�/�o+�-0ʹ)�*vo���EJ�ß���"32�Y��| ���^�Xͺ1�� .���]#2�Ar�n��I�w�7�M�3T6��<v�c�� ��E�=�gpm�|�w����n"�6FJg4���.l(P4�����5���{�1F5�C�-�Q�̋d=8����pi���L��֤�Q���%Lˢ��=,�o;��]®�a��u�tQJ��x�ԕ=���b�X�X�g�-9�2�	zp}z۠�i�Q� �kD�����f��m�^DH���{��j�#{���R�ȼ��_�`�ې%R��<�Z9ڤv{�׌����&�d"7u2"���)k�	�*�x�q�&{@��ΔF�QI���������x���5�p];��H9�L(̗�$VӦY�u���Zr1���_�5r�8����>�J�"���%�+�~�j���x��FṤS\�������8d(]�M�(m{��@=+ݹƋ�l�,�uI� �)Nc�W�;r���mG�
!��W��	E �7]Q�ָ�W쩙Ax�^����`�]�6./٢z:��� !\g���z,=Z��ބ�Y�II�[ȁ��w���C@6$D�-ݤ�*��S�B�PS�I O#�z��L��7	�6�:�O��"��YXo�����*Ym�Ad{��s�o�:��}3K��F��s�*�ƻzeB��.k�X	�{�J�����rT�ѭ ?n@�I=��s��+l���Z��#�����H����:��-;�(*�v.�H:�\�g,�y<a�/�D�FZ�ڡ7�E��������YTc
i��r8e���r�i���i2��-g�z:��v��L��0;'ɆT����@���U钉���-�9b����I�
]�a*B88ܵ���j��m�$�,+�Em�řW;#�L�f��H?�J"�X;��%�#ci�5�p��6�E|ךX���?	> i[=�𐔝�aa��)J��FV/և��֡tT;)'	�.���b�����<E���ZLh����|,��N��q�=՛2�J��t��J��Ch���+�e���E�\����;&q��n���W�P��m�`�H;�y�G$��f�ɮ_xh?�Ea�������
����jap��w�I�ͬ~�P�N�B�g&��$j�� ��r��i��#�ޛ�#6�xt�n��/��oF���\�F�΢-�a��:(mPD�@U���2V�v	"����mDޗS��R���o��1�e�d��%��ߏ��c���&M�
�s,·��8%�1��� ����v΍�
LK�b��@]E����=��_ 66�����ޅ�� b�=£�ͮ��R�ƈ�*�ZkO��T��E�	๋~I`[�M��gh����t�j����xȷ��ĚF�5�ci<M��g�a�N�is�m�3�Du����1q�\��D@����~ݱs���1R_%6߆�؅R���;7���}�ۚ4���W��������+N��a��p�z�����䇬=������ߞ�H61&�{�
�̝bև^>Z�����מ;�I��>�Y�B�cÂO������Fm%�n���
X�,h~�xrh��Nj�
�������C�"�"��Fx�ie���^kye�wحL���;nZ	u>�=A��O�����6�2]R��^7c~����[xA�3��^T�{{�,�J*;+�����cP�	�Y�����\Dy(�M����-�#��{�2)�W�Cj3Frg1�h�NGᛘ�R�]���`�j���a��=�S�0.5n��O��H��F�r��*�;�� fJ�WâD�g��pmw�h1�E(˝Th;ѾxԴ�rb���z�����Ok�Ȑft�%��5�H�Ge�p?��`��#Iѻ/#��Ya�q���%Ud
�l���q|����P�dj �� ��y��
+,م�� ���څ�ڊ6�\<xҍDV�W&���r�E"��-���&���!�I�G4�R�9(31t��D	����ˋ���������+v�˿�i�^�yW���!���A�cl�,P�v���%^��/�j�^��a��s��Jn1w�α�����&�t����Ѹ���ўl;`l�O�Ѩ��
���B�ژdM�8|�WYD�2��r��Y
F!�vg��ԩ;��k�����ڍ/#���zh�N��K���~@ ३�)�y��8�A�A�0俦_�h��R_�0��� �����N���M��5YJM���N����Yu~��d�Vk�m� ��7���jt�/��4q!���X�u������6�s�����-�Y]�I��<��Js�ߑc���Q~Ax���D� ��d�ݵV�b�Wi�<������P1&�T����Ty��yd��7�x�f��Wq/�BsC��������.@�iO2�h��D���k�8�nqcn<v��5����9��:��M��$h��u�Ͷ��Lnl�����}Y�K���������y�~���	��uи�!mM=r24�m��O<�.��G���� P
���������q��PSq���*���3ap��7�Z����hl���K]�i�r�����à��$@ۤ��=��x�\�޺�y��k#K"�o�xq�ʏ� >�boxy��rz˛ʴ�s
��ܱ�-�BN�D��ث�mUZ�݀�(��"C��$[ �h�����xY��_7����p ���f�rZ{�̤ٺp�2g��a��mH�h\$׶����</s�GV$E�}�R��۩tWsz�h7(�	b���G�!�wKP0B#p����rK��;ɎT�ZsA\�0����eou� �Z��By���C��B�a���ZH��V���ұ��>]=�d�o�V7��=�iE7x��j5�7�8r��6nu�d�``Kŗ����ώJhK�k��-5�����P���{[bT3�S�n2��vd��p,�|�Q%t���j�IQ����B2����ѸVVFyb��Ci�_m��Z��>���L��x@PX���&T����@C�����jvTK�o�@E�� Lp�r[����O�hZjJ��I��I@�8|xܩ~Rě��@["n_?��UO"(�:�nnzO�\����b��b`�Rp�=��	�/uF�X	 �o�f�ۮ�9�x~G8)��ٕ~����%g}>)6Db x��SE���������+ )�Ӎ`���%=;s�T��Cu�0G����Px�8������d�'E��EIS�+��<<��j��0��9]���� �d ����{u����4.)X���Z"[b����o];���U�Kd
�!�(_�b>��h�\�,�O��ٯ�YOI���V�=�y�I�Ra��~�u�Lr���@a`62�uu-B ���W�P���ECH;i�N�v�����㩣Ge���/�
|]�^S:8B6Y���yj���ub�r��ڨQ�h[��_��o�m᡾��4��
%2q�j�n[� ���x}�Z~'��'ۊ>�^;��A:+�2�/��Q�W��Ӵ�D=��}�S�2�����#
2���D�蓋lu]�*��u�����	��E9u�[��+hs��� M��&%��G1�
T^!u�@"#P�s�l�V@�_h`��i���*]�cu��:E*T��HQ��S[[���V��^�+����� �٬A��?M�����W�^y�=�g�UW6uu���LC�EK�(TFQ��3���B#Wčv�Z���,�x�:�Y�AiLӜAm��)���Űfs;3�4{a@�{�3�d�p#�g���r���~��O3܊����с�-,�d�q>i)*o��|�3���)�u-9��f:�%n|}TPS�qO��u���Fb4}�\z�ߜZ_�NJ m:�0�r5���?`ծ��";!=�&ܺ$ޓt�޶L��Қa{������}4K9^<��p�����U�_�3	)Z$���BE�Est���y�������/����4}	v:�n�������K2	���h����?SS<��e<�K�����0���ts�y�9ʪݔzˬC:��T�٢Ώ�x��,�n�>�*�+��Q�p�����C��d1^,n�	�67uy@�=�a��LiH��HNVR6)M����Ѵ�)��nx(���E���_ׇ�E�����;�y�-�C2���~g���f,�x�x-�ҞV8C�jZ��F7���D� �Q=Ud>����B�
|"f���pS7�@� ��\X>�bށ	��`��4�9]0�M��I/����#'��"��(~�#�ސ�;�BJ��"	L��~M\�[#T�ڴ	Y.ƙ�j��[ꫠU�b9��E9d�A0f5�pX�]�fs��{\Ʌ.&6�/-[�y�'���|Ňn�H�hD�~����Uc��V��l�`;��.k��8��*�F$�v���. 3�x��*�s��mH1�
*�����K	�0��ɸ��k�K�R�T�o~��.n�E� �$��%b�����y�؟]�^N���o5�'-W��|�D��� �Aiʘ!�ޤ�x��.�����L��Y�NB�W8w�W��\II�6�´��b��Cr�}A�0�����D���C�� �H��虄��\��@yP��N�8��S>}�vcw����lq@��R
���2~l���ȭ�ҍ�?�� ��m���gW�����r�Xv��~Iօ�a;��}�����:>�K�:��"�c�?�y>UK�H�QZ?b(����k��Kld���bP���bx.�i�c%�Q�p���i�*�T�D�t�'���-��R&0�:li��"t���wy��;��A+�D�Μ�Y�t)��ٗ�iPB�Ay��1QA�D��En3��OsJ��-	R�f� !����<v����;}T�립L�=�� ]3IHx�A5�mZ�5�Қ�<op�s�E�l?}?R��`���,�bytޏ��F睕�M�ea��8����o�5-TԻ,r�������5z{ A�*�K�����U�6X����$�t��BdΧi���At� �����T"������Jn��[n����10�Ta�"��T w�MHR-����/O.�.�僈�����>�� ���)��X��k<����Qݠ�3Y��o^h�E��(�^�;��Fa�)s���	;k�+9���7�짤���Q�>2E��0̗#� �<��.P��� �/7g����؍X��0��;��*�� 0MK%QH|tנ�7�2���M���g�7�dć4��#[s���	��R[d��p:@���+_�����==7��$y6~��qI��R@z�����*����������7�"\
�,th���M�̦�&.B+�㮸ƿ�?�XR��ܩ���t�zaP�9�2�i%����/l+e~>1�X{���֪'��`h�9y�6���BF �%����OcWBߘ�����A�K^�y��@����x
v,��K,���&��A���V�e-O�1�&�^�,(�ǣ��gW#>jݞ�"�p���m<n�4fO1QIBw���%�
����m:�WM}O�^�Τ��Ԩ͛���R��𒣋�]X�~s�`*;�r:g�~�!�e�P��lqՍfgm�Ѣ����o��*qgf����M%As(&�s�p������Jq5{��SV���77���T� Y�I�{k�H$���Ȧ^nA���'��OY����̜~&���Z�=�
��cw���=vG8��*��aq
A��Ǟh��r�~��fa�!��S�k�J�IK/��5����\�#X9?����)3���D���JJ��	��$��)��c�䖢������ovc�V������f����O%���V�v�e��7�(M�j��fk[[h��׃/r0Ɖ,���)�D���?@J{}��/�Q�z����ƈ�Y�����̍���w�itXm\�N�[�6:xG]�,�eq����	�'��FJ�[,���a��##�фkU�sݠX鏷AP"��m
�C��
��2-N/��5�*=I� �f�j����e,�ڠ0�{�,�֙%"��:b��ׇe2��|][8>��H*}Y�C\&l����c�x|.�+b��&�=�wt߅*�������,��O2@��)
p���#�.��E=X���s�T̲7?�+����y�gd6���������)��Ւ"Ō.8+�rW�����B^~q��~?$���C;���f��(r�^l �P�G�U��lk�6^�?_s=r�dACDv��!��9�]%�����?Zl؋�C�����h�R��fg�H���QۯLP"�s~��o�Ŕ����
Mb<yެ�@���xB:03�e�f���d[{WM6�!b{S˖q42����g�$��jH�Ѵ0���)���C�>Y˫�U��)+��}
o�s��9=�&i�]����wwF7��\�8��8�|Һ��SPo<.X��'�E��"��/V����!)����Eijj��&��)<���ƺ�����Z����Ũ��dU���KV��#��r�	3S���]"��79$�0"_��M$�
���&Y��?���u=i��z�����?�diM� <�@�A� ���q�g�C����P�XY��Q��w��u�b��Z.��	�Sd[���y��!��9��O��\����no�db��ڰ����(%���{pTY? �Ӂ6X�A�?Ϛ���+:��j��%��ٽ��P���s �^ԍ�����?���8�)���a��ЗF�`�|o%ɂ�+�-u�GC&�]_�}�G����w���YXxJ/��0�����am��l3��y���{aJR&=t�#j��Qj�d��J�kE���J,����*��^�5��5��]�]^9pl��/��]U}dU�I�O��(e�N�1�Ȣ�E�d�J��Pp���Ǯ j�7JA�:��������.��O]��["�Z<'z���K���Etj��u�VU7l6�����I*�>[����������4��3�a�	�%�$����4)ʴ�䁥`W��bW�P� )Ǡ5��j@G|�|��T�2a���W��\Q?Q��1?�	�>Q��{Ԫ��sn�MĶ���^�����qH�H�C,�I�u��>��qx� ���6&��^O����֤�ԡ�*�C+�$�w�G�qW��@x �~� Y�]y��ŖB��z9<Zn���+}����Z�>UTߖq�E� ��)��vQG�Bs���mcG�b��P*�uN��2���ȁ~��=��"���s4;�x�"y>�����^N�
���>�{P{��d_��v�f'���NW}��Yb��Y�ϴI����CkTxi% A
�U��b��t;����X�5�/ʎ��w�$�i��dɤ�nX7ڧ.��!�	:4��6G��}+��w�.�W0�ZymZ��_��&c��󿼉iJS�`�#s0��GK�Ed�#������uk5 ��C��̺����oYB��i15�Z�j����� ��r�U2>;�Cإ�*�[���`��*��Qi"e��?/ۦF����� �0�>V�.�]4Gra���9�E�@�cd[�ܞm����Z�tj�a�I�q�0q2�r_�Fd`j .��Aff�*����1o��;������Y���S�8�D����`݂A
B�{4�$G��#�=�d��7yև�f��j ���I�`Uɪ�\�7�"�v�#�Ro�A2x��k(%Ӈb-��0f�XT��T`^<w�p��FOl0����$��!�$E�����V��T�X'`hg\��۸a��(�6�U1�o�T`wRP�Okt`f�l ���{ +���qO]�w%��As�^�	����(̶e�
'.1��xқ�c����C?��lNe*ֲ��<�+�*V�a�P��K@��9&:&"6�J�F2�H��Ba���.mIQi7-��E|��/٢'di�C��+p5�Q�\}g��qٿ|z���},���m�;_nn�N2�o��	xܥdyE�'�i;�L��-�c(�oL�'-���`ѕˎ_�%�"�O>F\`[<���}�� �)�k�M}{�x��^���<m���j����F���������E�0�i�#��΁���ٰ"���>\�{�"��i�N�r5��5x�6C[Hz�I�����}��3��7��J�17y3	��읷Qr|G�ٽ��7D�,�舼`U4��}K>�|�%S�3~^z ;��$R�OZ)��a�����)!J�k�m%�&������}av�ʣ��`,�[0��)<�5/�����
�p�WW�xg�TI�@%�}�A|p�Y	c�����S�\�g�'^���� 
6k����Ȩǽ�-d�t��<�'D�(u��ι=}U�1L����~N�����������ܥ�mT`��������? # ��.�<�w�" �K�� cPn��}��"ni{�?�z�]�@ܑ�V�1�c��x�y�A�(Bmǥ��qk����T�`B�����D��3ن*�V� �X��S���ǥ�i6�����X���n� b�dqY��԰h�� ��+#� ΂�'�*W��^&C�j�J���y�� �jh�{c)����^�)X��]\'�ڗp����`��׳��g���΅�d�o�l��W�&e�����P�T���T���s��e�ױ>�@�lI,ϟa�����!���8���?�g@f��
z8��2ɓ]�V���){4 �w\���%��.�'�yn�TEs�t�bo>�1�щ/�����{
-�;Z���"��� ��5^?�fvl��0�� �t�hH�p�.��p��r�����`��!�th@�t�����e�Ysi%��op1l(�x�XJ����	nZ�/�I�X�^e?{+���*��y~�g�����Q?�^�uF#+%�)��$"�H�'	M���=��O���P�`�����(�'�>�'�b�1�1��i�H�QVl-�9��ۘ��>��p)���ً�i�<S+��o�.�g5toO����IW���C(/�[	ɼ���t�����f�:���6���g�\��1δu�7kzzM��:L�Oq]h�J@����r����I��
9��2v�k<f�/�I��bp��]��Y�p#*��;���[!lK�/��jΎ(c�.����'������&�Eh2T�[��L�ڍv㹺�:��_a���i{WV�7��Ѩ`����[X�k`�,��{R�@j�	�y����:�+f�����?��"G�H��Pn�ˇp=���(U�P� G��cp�o�6���� �:�=��e���O��Y���+@��}�Ը��ժ�����r,�8���Y�U�hŋ�&ÿ6�r�r��,�,)#5�J̷���)!f���J�W�HR��ԕ�:* &uOL�]�{ 77��A��=a�;a�jK5� c��D�l�(�NI�\�N�t��c7��R�IeuC��X�5�k�7wn��#���/�n>��zk��EW��<��W|7FO��棐E��� fF��]���f�z��Zh����`o�8��-BQ��%���c��s-A�-�摝"]ք;a��U��Kc��%�A
gy���]V��큯�x&�)�(8v�_6|qQc�:<V�˗���N�� (ƻ傢�3r�J�'� ��M��"ɧ@n(��$�7��]���c��-�}=���t�T�����Cje:�x�颬8=�}t�5;?f���G^�إ����a�e4��%~�fW�R�������t�?v���+xEp�/�Si��a�@�eW���x>h�Ɉ��A�ŗ�R1� �/��):Ո��ܾ6���u�����g�r�W����pk�nR�ZX7�أ<?00�w��~�\�����\O��:|xO�U�C��R��'�6��ِ�i��:�N�2\u_�9�`�|)������;�w	`l���
�.�&�	�J~�n�e�-��zܯ��d���I>LW�:�|�k�N�
�G���/���*.�J�l���E�G��{��<�HD�
�}�P�Q��qP��i���;Q��~��/��f|}	XZ(!�1��2�A^�\7Xe�o;��r������T���+I��AJ����HI\��b��3r��������vfo���L��b��C�3������Un�)�jߖF��������?���u�sx���0)<���`��O�馹�D�4�i��m���.8F¾`Jn�����y׃�5U��k���#E��Eh��:R�(�._�/��OZU�%�P,�Վ�'6{L�v�)��/1.A��f��N1F��;�},��V��b����,�������\Bm|�&a]	&Stv��LK��~���ԓ50�����E����w��-�sT|�K���C,�0ԭ����$[|�/�� s�;�ZĎ�\i�](�b骷�����_�p�m�:��'��z����4������x�M߶=���������LA
�Ǌ�]�lNH������������v���6����$�{,ELC>]$"��J���瀌Hď<��4�|�\�gR�\Qţ���q�ɫ��n�õ����8��5T��#˒�.~�i%3�v���7O�**
ĸ�[����~MA��l��<�M�A��o��4�d�e�9c��桖�҃�V���o�ݹn(2tR�)������Ҕ8c��m�"`���ڌ7
h�-QZ:q�K�{�G��}�ϋȇ�I��"6z�/uL8�5����u����9Ԛ_��U�j��b�Q��K|䬯��$�8�1�� H� �li�^J�?�W��=�1
�sJti#y��Rtּ��W�H$%=x[��Zc&��ʝ+��.���ّ�:}^�����|��[W`�wDمE�l�"�8	f�%\��B�*�JK �%[�܉0d78�x�j��
��%S�z"����||�݅���+_^[	V�#1r��x�
̭�A��0�c��8R� �ǀ�󍭁���	��8��$P�=��E�v/��C������u��?�*���IYU�P�Ҙi>�D� Oѽ7Y�)c| 8 Ì�
ч}dTE���T���߼����>�GD
���㋀n.s,�6�����*AF�:E]�h�@lUY3A�?���C2�5ʁ[#�qj���RxŞ��E9r�m�:*:n���j��CY���ZW>��0�����DD�#��E��u~IV-��z�bs�jo�X�a���+����y�w���n:��[�Y�C{g���]����L[ap��WD��.�r��/M�܌�iS�1}�OBo	���`�����})��N� _��6��q�5�Sd͚��{c�,7�6��U�⧣�/Ci�^a����rI	Z����%��m&�~B����bO�{�K򀘸ǘ2���I��"|����6r�s^{+�mV��N%�J�eD"��м�v��P��Ѐ"��̟�:�;�*Sl{�J�"�Q��n����|�l����&\���>��/�YŶ*I���[PV�n�N����%T�~Q
ݐ%f��i��QIxc��ƣ5�g%��3�
@k���rD�H��S���>"���>�r��5�>c�s�E֍^$�l�a!��F�M7�����7���>�M@�b��w@��,���h�(���M?1 ��X].�yD<�;��|`E?������W8��U�7�"�x�����C�+��2�}�u�m�Qi/�'`c����yS��-�l���6��c�&�k5h	/Bde�,����2�Fm�����$�֬t�;���Ly�Yz[��n���"�fO ��"3��D����,݈z�N�����aʱ-����K�
Y�&��d��j<w�{�2^*�w�,3�t���B�k��OШ;ǟ�?t!%�b�~��6:Ku��V�Q9!e���d���|��
�m����6�� y�`�uۼ*Mn0Nu�n�S>a|"![1���MA]/7�_[����>�8s-�zȊ���\��0N�P��vL��"$8)-���b�L�>����ɨ��A�@��2$�4db�7e^�F/c}&J�[��d�9=vX��闡�P�j�� ����}*�̕&3��nJ}n}]-��p����I2J�>��ՙ���V����@�E��B�/Gp���#&B!$�
&)f��L���6t)�3���ހ��|��`�R��,����_���|�fV�a�1JCO���'�뉼�2��J��&Cs7]%0&�S�Xa�%���6H�rg���g��"h�A�T����a�T���=�~h��e�	��G��>�=��XF�=�C�����iO�ύ���Bz�*m��>�+�&F�<�ϓ*pH�|�ج2��8�f�h��V����v����v8LB�����G�b~�TO>w*�m�w��p�#��XJ|��/'E�䊸"P�� �����5��QU�>�D��n�
�����N6�@�:���Y;�����k����o����?��pb)�^M_?17���F������nr�Z~��f_(G4(��Ux��RAHIb]]n���݂�.����0^���Ī��Q�9-%���<n�{���J�ۼ��!%�$��\	篧�s4�6���1�<�xQ4mR�!+�(@yt�j�X2��#u����R�;��f�����g�^�d�KæǶ�݊w�4��iB�dЫfp/�!����s�r� ���)�:k�kb�w�FӮ��Q%!������ZIiM9"�F�W� �Q/��C
�w��J����`Rt�<��{��qWi�� ~�\p�ɵ| �L�{E��h�sZd�U��M��P�Hn/sU�3�2PN�li@���3����K�.������R�0:H4�	�������9�g����>(�^��(��tR�KQˣ��p̶U����+�Ց��ъ�-�Ѹ�s���Q��FJ���L�f|��rk��X!�C'�Ι�6X���Z��{��q�X=x�3�:z8�������?5������}��.��A�Q���
3�m`-�G{E�m�^ݦ|�e�>�LYn,c#�ҥ�w���sT��u�{g!���i����=�s�zf�*k��Â ��lg�Sw0|� ��L%:,�쿃~�Eؙ|�<���u^K��$�uߝc���]�;�x�o�WM/���H�Ex��n(�av�DXX�Ơ@����g�Գ�+p�#�d���0c+���`�G;𪌫_~���0Z��7B� �#��Rǋ�u^�C+��*I	#�~�vx���T#�n�9�{d�mM,Ȉ��Ǔ(��%�s,N�%�˘ �����Wb<>v��^(W�D"2"OI��I�~��׀�c_�� a�������Vp`w}�C����Q�ڲ=�Lm*���5��2iZ�+�X �=C�$#��w��ߘ���8�6�{������Q/��,�i=Ԗ|�B�)̷��Ffb��s�(��"NL��/�sL\> ��=��]
�>�0}��M�Jl�n�����gH��5RQ����%RvA�9��s�b�ƺ�Mz��΢^�Q���� �l�IB�g�p�������ڥ�E�/���l�j�R�n)���I|A�xA�`���F�u�/�f$�eð�����6����o�O� A�?�"g9ƑC�d8�2��?�ب6�O3�ݡW<M�ۯ�GL���c���Ѓ�Ҵt�1��=/�m�p��\�ړ��W8��$Wq��^g1�R��Ls���p�&�#ovq��y^���U�f���J�b�d��_��}�ü$WrE1�m��X���%���IH��'#�=E���]n,��m����r�z#��v�i�9�M��b��,[Lx#_��ƙ���i��]��YA ���Q�6FA%'R�-G0詇X��N���f4v�g�iu�R\���͆i���z��L���-1��#�S���7�b@�κtT6�z�چ_s6ȱ�5]-
����=���Ei��� +�vHP�ȍ@( @�0v%� ;:���em��ȉ�Q%�E(�����9]�3+��`L�nb*:|�e��x�`����X��M�p�r =J��xBZ���Q��#n���6,�DyU7g��A
&Ёbb~ ��m<��0�j��8��h��H����}�@]a��Z8a��L��sг�c�Q3߻�*&�;��w1�YJpw� �n6����8/6�7I���[^�p8n����'���X!�M�w��|��(od��R�Ҵ�Q;�Xh@[pޣ��js߰��4z�����Cf_fW_���+���6��Wﾪ��r{��3�m�D��m:#ꈅt�H/�U#��VS�^�uG����{*K2\�� ���NH.�LX��hHv��l��b(�U60��Sw�C�@�ޗl=����۰�����n��ſ9��+kꄺ)/�J:�+?~`@���RD¨Y�T�r�Z`���_*1l����p{:y�
�빏"q_����_��`	�'b��6,�ɔt�T�|�{:�}UV70g>�Rd���=��*�r�+K2���$��)WY�x*r�[����Z�'6�r����K ��v�<Po�g��8r�5�B��X*��1p3��R����������O�b�\'6��Kw��ʨ�$�T��sFXCa�:�uBa�g9c��C>0�2*nŘ������RA�Yɴѣ?,k� ]S(Xp�J17�J��d������m�w����
ʤ���t�C���LeK3VWW=ư["&T���F��k@u� {Q�8����,�G�q�S�i��v̊�K�j�-q�缣0F�I�(_�ߝD�n!�D	x�1�;*
�L^py_v.I��IܮfH�<�g%�k�`U?6~�?���Xh��C��*�/\g�s$��i)���M�4B����o;�D<d,�� ������<<�&�ͅѽ�(I�Iq:8����:M�蕄�5�\W}��� ��'2~6쪅shL%6�ʷ8 5�a/_��~��l�f*6B��~D[��ן�/L�<��0��z�^�H���5w¼$8d��j�����h�	ʳ������>�F�փ�:	�-d|y/Ή��~�	�b�ŻX�ifDk���p#���4�� &q�@�g��k:���z�q�_�hBp�]���tȴ��L����M�v��I���89�c������e:�6�,`Wp`qL]�lu���; M돆��g�ڊR��[����'�~k&���q�:�W�Q�wE0#W�,[7;��H�;;��l�w�Nq�CU�QJV���}��z��d$YN�6Mٍ-'[}xN�+��ZyR�f3򙗈,�Vk����V۷���.��Q��Wp��R?��sC*rԓc˾\�}u�~lΚf ^��y��1t�F��C����f+u"C�p�l�@L��>Ө��"�Ӆ)��M�y��9�n�^�=�����0N+�x�Ƅ e����޶�k� ��+3�?�ӱ�q�ab�9��B|�O�tP��k䀘&��5��ѳ�@��@�&�:�ѱX��*���g����)���O��	�������[8�.��a��<n�����N6a�l�J�6�0�𸤱� ����I�ns*��di�)�����Q*'�(S��wğ� ���x�戗��A�0F_�Cw\����@k�)9L�4@�f��d�o_\���F� �o.� h5��*�����{�7z��>��8jHVǛ�T��#��������ܞRV@s4���8�� !���h��mh�a'�b|@�G�ƅ�k�n�[�)��vT��+j���D.(��]��ؚ�� ��P�ҽX��Z� Sx2l����.#�+�����f���F��Y2�z4��*�L��PoP��'n;��Y��C��Q=`E%K�1���q{�E#MOl��>q�I�"_���y[P��I�	U�S3��ȫ�{���FE�7`��bFi��%��]��#Wuz��ո���}zP�������B�g�����h�a>��F9�7)��v)>f!�r�)V�Ϳ����4���8?7���jE�\v���⒎���2@!-��ЉdSV����(�+�8���!b��V�������~���-Q���g֌ّ�F�Q�)�~p������N3��m�%�(����u4X�[�����C��m;89QY���X�V��S���&��B(���'S���#�,����o�cD���W�����A�����|Ɯê�8L��E:��Ԇu�{i��jF�X�o��7��q�xE���[W�ɛ9�S`'�����_e�ف�\�+	-����߿?�6�+5�a�(�jEwv�����U�{0?L���1t�y�3�O��EK�1���`��7�!���/h�	|����&��À�8>`��l���Ϡ'���A�2\���	$������E�V"X�`�C��d���$a�YS�1���x"��>���'�I�j,dp��rBOQ3�K�g\&q����v���Ϟ�
3��[
#�}uVV}W�:�I���6�\�����Hj۾��y\%�T2@.L}ԙ�!F���]Ўn��������Ю�'���G����jo��r�,�Ճp��5����ʙ�z@%F����ΩsEԩ��]�)Iv�u��^B�[[<.��B���`цR���Q��9�l�m�6�䃄l]��.ߌ�I��.C8�SU���j��B���av���X�2���
�r��M�⠯��?�t��UU�&�G[t�8�.�P��j�����hOH6���)$�CQ�2.׷�;4��坎�a�lŒ��J�᪹��"�ch���ҽ$���k��nm��=�CU�M)�O}�������EI����V�O�fR:?����	vT���ҋR�zGX'��Ms� WݴIl��3P����������WĤJ{�1�y%�l�PK���T��9n�G���X)��KS+�3BRJ��]�}��u��}4(!��-:w1�A�3F�V։"~�ꆣߟ�T\'��OC Vv������	�<0�;�/�e���i$֖b��
��e�/�~���=�]*�ê�m6���轎23�]XK�Y`~���T��"I�XQ~Iq6T�bs�c����KX$��?��ϱ����B���\�j���^�70�8���2�[pv�j�C&�nƓs��n]��f_zF h	O�G��t�+�:T�u��4�^	HF�	�7Q���WҐ�Ke�-+���@��p;�(��cI��E4�y�.f�y���0�
hF�'�����n��O@���(��C�H��s�|ԬB����g� I,��q���de�l��Y� Xt�>C&�0���}��������ʕ�؏y4��	�K5?�1�wK�M����S��<>��?`�߇�It�+y���.,BUs�a��~<t� ͼ���|�`����=Z�1m5$zu�}$\�T��I!{J΢�)YSZ�%�X�M���T����Z�&L5�6��"P6��'	f����ț8��l��bkg��Ooǧ]�:?2U��� !���y�)���Љ0��oE��к�6���L*T���b�NL����h��'��%�|y�B��qn�e�al���k����E5�����N��o�٭�m���ef�5��^�Pd��M�n���0�p��s>�L��>�n~�V����%���b��8�D�ܿ+���9��"Z� ���ثS�B��ۄ �K�3^�sk3P'�s7c�"��v��eC�Fo<Z��+%I�L���!��h���e�7��2��I�>qg�>#���<��}��rp=�ſ���@g<|�@�oAZ��+Yf�i���-��u��"�$T��՜ۿfw�m������g��!x�ٰ>s�7]'D�9	�l2�m��X�>W���޳
��1�u�ɕ��3��N$Υ������B�4���Ǖ_fm.r�xqt�lN ��w險K�Q�La�M��%�����>��Y�d�P��jJj֯G:ڪ�{"�^�I����I�z����	I�o�ݱ���33MR�g��9⬐����̓-�6�3�Ze���"�Qeg�R"o�?E���ܜ(X���q���	�zs�I����1P�W4�%������R!Yy���-O=v�,�:
d"��fH�5`31{oz�`��` 9ly+-�[W����V�e���nV�ϮZJ��t�n��M�v���'���s�_�}­��݋��]�:n�����3�
��E�N�+*�O�"|�Hb�fC��?�I:��X���`r	c{�l���$��'��L#Z��5[�7A���@�cvNI�X=X�q0���]{1%�(��P �|����5j"~͌�MQ��Wd�������	fd��Ix�_�]���	aٯoQ���m�r�>a^ϑ�������3A4�e��X��xI�|��o�o{��yF2P�mj��$����@�b�113�3� ��7����1@[�D�˺~�]������0�f���k;������x�j�W ^~����_�R�$.�������7�YG?
sz"��n_��'6� :�o�������vg4��шb�0�;�W����ʖ�>�������t�V�:��O�N�M "�`���!�A�"�^�A���7�[�� ;�ɧ?���'B�͘ mo�I�p�S�� �z�կl�klKn��<7e�a(������Z�q��ш>�j�y�Yu�A�+]��ql���	��F~`P$$ .����ϐ!�~�.N�lC<�7�(jq�JVf��H;�Lʢ��iR��E�5�W�b���3�o�pm���z&AJ�,�~Q�foP5Q#�;�x[�Я�K�'��	-,���{���X�W=C�W��������%��ٌlA�����	_̥��<�%�WM�`��ߞևʋ�Q�bR�V{�����l��VyC��|Ȏ�	�D�zZP�ʈ���L����&yؐ��){h="�6'���J�)i˙Z�cĩ!�}-m��-��t�'�J>��[�,N�Ճ0�����A��/N�m⼈�O��~�����Zۗ䞠�������
��]R5�,�y��q��_���D�c,����M��s��b�K(j�4��t�2����<�P�A2;0�� �I����ǥyn�NV)h�єt�Y�Te�`��f$cQ���wq��4���G��Q�� �e�u8X�&�QNs�͉�~,�9�5��4�u�k��&�C�AboJ�}S|�Zs*Lҳg����9j;2�[�_�^�b�ֿc�e�|��`��O���4�p\�����Cipl�L>s�Փ�Y��8�[,v�Ry��y�6�n�-�]�ڐlH�,�L��j���x(H�ab:�Ӣ���.Q�"ن}H��gl�ĉtR~U=�p~S�W��K�>IK�N��e�3�����?�� ��|�n�넊�`���vٖ������}C��F���J�"�� �W���-#D0�E$-) ���
tN��=�&��Oi6F��j]o�6	$���+��ڗ���e�oq8�k�6Q��LK(I�N�M���K>R�=
�2�ʯǕ�8��Kީ5��
~�s�oQ"�>>�����%�O�j?�uEK�v��D�2���>�(c�d�䖞��+d �<B#�aM��=8�
G/_�Ju�F~򧸂�h�� Y�Z,[[Q��|?G�H L`�\~���5�3�|�Tu���w����Cm��%C��T�sϥ.5�DC_Xi��B�~@y��y�W���3T���>�JL�L�W[m~���h�YBN_��Oο�Œ/W�1T�Z�7��|Jޟ��0��a!�mfvoh"���pǓ��*X����qP��7,w�*ɺ�zl3+((�h�2ڛt��vԴ��O�1R��6��Cf��%F��F>�f21����it%�E!^P7Y�H��Ʊ��u�ٝ������e�֬Wmg�X���s]B�6�����(l��Z���e99���yMKJ%H>�[�3`��,o�H����I2�A��Ģ���CiYľtv�^t!�+�L�si#�iE�s����߈��,�Fb�U��f·��Y��.T4�}�S�3��;	���S�u��9d�:�ō׼�H�f!qk�j=����� ؎lB�<�[�!E��8��=���\����{r1��R��I㲎�5�`�e�Ԗ�sf�K8�߶��#���>�e�ݾ�"�V�Uk,�Y߈sV�t�HEw���ā f�
v]h9���r�+�o�@_

	\~�1��}�ds�$��\�ʕ׽�S���;����zU�P��I�s˺Z��KƳ������z��W�ʀ0��rlRs&a������$��*RS2�h,�1~�[c
v�*��-=&]�c��So�ؽ`b\6ՙ��9�;.��oܱ�^���3/���)�c9�^��RG����A@�L��4�x;B+m�[_�a�j���|�\7OcZ�.}!�������9&�}�Y`�oc��w������,��eP>�}|}�m��5M)x��/����}�D��c������� �bD/:���ʡrS��(i�+M�cD
��	�c��P^.�p��U��s 'C�ښs�7�b/f2���(l���H��C�O)�y�M�[�q@�}<K"�`A�}ܖ^�vL�0ʓ4.{�u�Rc2�t�'�tK��Б D������|�\nZBD��Z��J%eRX��;�˨��֤ O��B3��O�W_�o��64??<|~!�G���A/#�!�Ī���X�J��J�k�,��Q�͗�2��<�By��d@��p��zF�!E��e`��7M��OI�5A�%���Vd�wj�zq�,kn�
�Qw��wjF=�艛"u�x0������Gk�_�K*b��ǅL�0`IÉ�*y�r:צ�͞�|A���1�/�y�u<E+�SJQ��\g��]������
�*Oi��X�a�̠���am�ڠ��.U5�j&.�_�_�LJ���ѧ�2��S�3���Ҿ4�[���ʡ�(������U�V��h=ݺ������+\�d��� dR�Ƨ�gJ=���;8�.�a7qJ��p����ݖU��"�t�j��m��G}4���)-3�%&Q���-���q�]Y��BW��i���Y��t�y��7�����+r���o㌪�Co1L1Z��̛  =��M�[=�(����ʩ�N>�
	'��J��Z�ܦ84#��`�X�r�b�ُ:n#��vU�����"< ���(z"G�mn�Ɵ���S�s{��`v����W%�4��vO�����#3�BW�I��߿҉"a� 6�^SۋO��ם�#1i��oU�uk9T�cN+M�Dd�ߘ�k:��P����%��v�ɩ���@5����c�e
�ar���J�?�Nt��C@���tA�$1���^���,/��hbe%!W�9~���s7M���K�V��x�[��oI�F	�~�)����C�Ǣ�3�Qw�o���� �͂:#`��p�l���@P��t�	J�{�}���F��V��»G���~�"$S�A @�lygD�ȿ�f�YN�A~@��;Zn���C�4�+;�
 �+�����_�Q����W�	+��������d��U]�� �j�#�#n����ݾ|��Xdl?`�C��f"�R۽�9a�9��l�~�/���4��ϙ��y�+NF�-
� E&�>����D�G?�N���;i��Ʋ�=�#���B�d�54��";ȉW�CH�#�Ƥ��4�����n�h�Y��m �������7�Fs��P��PN�a��Y ��Sm�g��%���\��j����$��"��"@iz����i��VJ7��G55#:���AшP�{��D������g�p�6.$��89��!���w4R��}��݋�4�1tZE�(�w6n]+X�i<Z�y0z8��ٹa��x.o9=Ij@~$A�����%"
�q�3�zZ954n	��mi��Z�๤�@u}��u�e�`���:b�m%�V��{��1�{; \0��Q]�@i�;g��kҡ�j��u��ر�+@e�3�B{M��<��f�u�������J|F
oB�9�_9 p���'atn��-��K�
j��8����Ϙ?ϲ�W��1����l&�ѳ�ȍ!d �����U���g�u���Ƙ��E��;�+�
X��E�A��$�����̳ם{�qE:g������:�X+}�-qS�������3�Q�zLr�,���B�J��yƦ�̌��DH/��[GW2;U6���6�L��l%�z�@�F$�*�m(�I��&+�`&K�M>\{�v~-��M��ei)iG#2A���\�vL�uMh��H6z6���Vر���U�,�Ӥ���UsC&粨J������H/���KES��f��o|���69癑�'�gI:}��::4�r�(����ܿY��#�M
'Cg�R~����Ꙩu�?�k���-Ή#O���pB5����A�r�!��aC��eͩq��x�c�Lr�X�O
�ti����g��ǝ��c�A���n�r������b��`Ƒ�*v�c�!�a*��H!5�95������C���]G�O䞟1�]�3��O����~�yn�f_tg�\�i��,�*-�5�0�Q��z��5����{�i�z��ƍ����)�J�0l�#�W��H�`o�P���Fg�'�</�κ�������\�����A�6�l�'���}N�,L�;��@|md��U���w	W��:�쇎���*�Y�G��c_L��� �hL%h!�rj���Ň��_0Cg�g7�ψ��,Oa�x�]���2���,�j�ί���f���������^Q߽Y�rU�d�S�GWjw6'��J]In졔>� �52�a��T��W�a��@��h��#&�N�M�h9���xbG/����n��/F��|i(l��'�A���1;z�uH, �o��� ����~�k�s��^���5�"$he�˹���٦u$�~�Bu��-I�>��Z�|C'~o\��[�0��/!�;s�M?��$c�M���۞�p\f>\��X�LKd�jY�tL�_|��u[��ޝo�M$�u��>3����C��6���[+~kLԖ8Mb0�Q	���0;&.��� Ȼ)	Q��P0�܋͸������_e[@��r� G*?�,���'��z�p1ǊJ�P`�I��^�
��X��*,��F%s�#�&��gKUn��؇T���О�9���4�ɔr��ԓ�b�s^]�8����j���R�x�M���Ĳ���mvq3j+v�ګ�j��� I�聜|OU�5�d�UR�뻳��A���y�L�eo�V�]  �+�ʱWO2�T���U�Z��꫱�RAn���U5mt6�TV?��(SҨ�=d(��m��*Q3���\Ѷ\�����n��7�H�F)cH�+=�q-��DZ����J��a���m��IL�lѢ�ψ��uR!g�A����W�L���s�Nl�'�F�����,WF5����r�]ƹ�2a
b���P}�2�qѽg]9:k"6:�؉�N#�'
�3D��Ӏ<����hMpy�v��빀�tl&z�i��%�aP�c���$S���L}~�᜾���H�2�P��7�َ.�.M.�D��(F��WA%��4m�l2j<��NH��~@���u�`n-���]�����exO��eS�H �s��yȵ�Q�s���Ed;o���Mbe���AX��AE�s����!�Qơ�9�l�\@�6�(�)��ue[��r5��F�B�������˴�P�"��wτ�-R%n�@7�aU�M ��MI���R�/�6\�'vK`VhÊւ1�@\�RXd�G��GX���=��;�B����tYk�( ��~:��{�����B�ib�=��°V  /&�9�Ԋ�)+�e��>m[`�0Z�ν�B�ds�d�@�U��%^j�<g%�y?Vk���c�*�S�3��۰wtݜԌ/�����k{)�T�x=��{�5u"�WY7?���x/�ۂ~����j�`�	^ß�x���]Pԧ�J *�f�ٰ�an䏧�S��ƣ� .�#��Le<Y�{�#��lm��g���8��6K�D��mQ�� ��dj�oqG�G�8��O3���T�2c����i,rUŀ��J�b�oS�a'���c�CpDL��f�1��#��-���
�.�s��0
�� "���-_YB�{�pb$*�+X@G6'�ˢ��;�;+��[�Ž�����BTQ��y�a�"���G䬃�)԰7�<% �)V�$��1 \"Ut�&��l\�]�3Ve!3��-���)�n2�Yn�gz�P����t{� *�zvs;�������A����֬侲��DI�.��
��H�v8�,M<�t}��!�
ҡ�?#����",Ǟ��H1�k��K��L�7<Rx����"⾥XQ��>)�t�nTA�eźC�$��eaτwC�c�^���l��6j�s�C��>�y,/��G��W�4BBA:u'�+��]e��A�#�#>i9o̬���MU��F-�wj��|�̣"��Bé�i��Q�8*$�Ŝ�l�&ڗ;k<��>OɑP��r�����)5H�Ry�x ��XoJ>�e`��=�� 5�J�;e��\P_}�n�YUi+��L��m�r�`����խ<)�G�� YE�Er3l����V����O]S�Tx޴E�=����n�Jׯ�<��u��bW%XK!�x���|dKQ����k�6~��8l�c�r�Q2�Zउ�c�&}N툷�՟S�\�~H9�}6f����{��o'!H�c5��h�rC'�d&?��p��/)j;m���o�(�2K���
���C]d׀Ci��� ;�@\!YH�!w����o�>TZ� l@�����^�
:Ѳ��
�b�\��68�� ��-Wup�^�D�	0TI���hw2b��Gi@D����BoH�,+I�ׄl�-�J4��o��!��7�*����S�t{b:�i�GB�4�i� �@׬$�S]���j�GD���7�m{��
]f��'��1	��K�����ϡ{�f윪|v��vρ4�?��X�s��Ok����l�|7�}<*`�6�-"��=8�-�f
ެ�ve��H;�v����>HŶ�gŲ_���ۢ�^&��ya���mk��w�WO�Y��5�A��1�K����q����Յ.��h9��v��P����T��)��Un�g�&��3�'��b,p����d��șkT8j�k4t�� ��7/2��|�e>�H�ol��K�|���[��v�	�w���w�G(g{��ڴ�*�(�K���% t���s��u�+fI�E��!{���.�@@�g�Ar�J�M�K���h�<���\�E�ai浏4�k�}Vt"0]�c�)	c��ux����y=B(�W���͗r���|"_�n��8�����~�)Nq�]�����Mv��u����aH )�a��l��U�ISt.��W��Z�S:�]`�Ҟ��~ٞ�H#*�G(��V�e��.{C�_�ff��7�!nZ��5���,��Ѻ�Y�,�?���j����@��~�����8����'��+��ʥ� v��z�� M���PW`�Y|o���Y��Z�qj}�6��T�5옧}_\t|t�Q
�|K)���xBqDhh[T�z�91-��Z�"S�&� H�*�Y��̖|�j�9y�,�����GN��N�cHg�xlAhN�����5�ڨ;�Ԡ͗�qs�z���nE�nF��\ŢsyB�S5#G�-�G�3�o=t7xf�X�\�4��k�A���l}a����S4��^�����\�lN�[<k�^	"�gĉ�R���UJ���Q���`ֿ �/r󋦃�RfD�{��nh�v|^������ۖ#�y�ÈG��\��{"�4-��/�J���/�]#^�f	��Χ���;6B �U����V��ȑe)e\�Q�uO��';��c�'��En*����(�.צ}�M};�1L�64&:���W��|���\I����I.g������<�"Vdun�t�V	z}=���5���2�h0� ���0�Khw)	{��d��V]��+o�C��!�ߡ�Z�ޡ`�$�|���c1��$��+uz���{�'�W��yb��"yW�B��R.7z����J�P���~_�����MN��Rd(B\<���ik��	Y����V(�[�����*��+�U�i�7 3P>�ZO� I��m�R�u��c���f�(;�
S&����_{�{���)��!�����8�=���WD�+���Х�6����2 ���`"�z����f=º�5�:\]5���w�m�_�?ɩ��<�7����m�D�gܺ� �u�s���*�z|�&vK�X1��rU�1kX�n7��I�!�F�i�G�71���_�� �:㻿����XŤp�>ß��o�R���kn�vX}OȒ+�H`�կ̘G=�j��� ���!Si�6�cv���LWZ:.:Y�UǕ���W���rWM2�ZpW9�� Y�&914��+����v���ͣ����o�,���u��ߐ�?0�m�n�f@~��a��}?�8���9W�5y������NK��d��2d��:�*���!�{�w!y��Dឞ�~�g��H��-��Lp=�糵O�0Y�E��pd�+g�zu�iY��K`��~�IC����iU������? �?H*u8��Ö 4��C�)0�pPn2h�B�R[0R�u��0�s��2�o�x�O<�Fh	D�%{��<Z%�Ҷ;I�:H�H���
�<��h�F��	�_Z*z ���շ���?��;2I��SCY�m�ެ������^k4�f�/p�D�n籍��o�@��p~ˢ��W�
�B�x�lԄ>/��y�5W�Nǹ���K��AH��>���ߨM�c�~��i�Q(��He?�c�PYc�8�&��I2�`��ɲ$Z��c�O�|Ly�1�@�	072��]�Vg3����t$���%�|J��I��p!�iڈ+����y�1�>Wxt�k.	�mV����
�5%�E����"��Z6�m�0�Y���@��r����E(���5�Uc-�u��Rx��s)��at��$��du���ﳰGqQ��Lm�'�X� s���,���y+�RևB��J���F6��a˦�R(��H�[��ė7�4��D���7W���K�WHZ�Vf�Ou+���Gl��WO�H:XOV�d2W�Fc1�4f.�G�S!�$O���%)l�d�Ti�}]ƫ7����B�q���Dm�R?��&$��b��3�J2���<ԏ�]�-S���d���ϋT�5j�1�j�y�u鬵���svv��5���������|ȑ�~�������8��^���Q���S���PbQ�̚DZ��$�������{���Ι0߬ ׺���Q�QZ�Jh/O�~1�����g9�
�5�!��g'@������t���h��Gi�X;��+���AL�O�g�j�n�t�'�Y6w�U}Z�Wf���ힶ�0��4_52Å��[vo�%�ER�4%t���7��9J�7!'"��y�E*�5��xb��/��w=9Y88Fu������u�����Mu.==Z�Ω>����K�B0E�F�4uCQ���λu6����GmH�V����LkvL�S�U@�����f�.H�,��$��<gP�W&�o3�9�pYe
�9��&{��9S�l�{��?B�~ ��,M�J��}��bI��(*د��1QI����<�U��!�ޯ�6I�T$vR\y�^�z�@��9؎�$:X�nW�xm="":�*�o��ZqL�X#0B���K�9�L�}�U��r�4����y�JCL�%��ɨu:�V�u>�L6{�Z���o���4Bљ��A���z�'9���;��8P�_��5��:��h������c��ht"d�.{s{�A59J��OA�5��g�o��w_���&r�/Ӗ������j��h_�>}�ᣟ�y�����?�	t��3� ��4x���Y�S��^nC1%�����r����7~�'�c����K��F������|_��K4�^{����V.�sH �o�P�S��q�R#)��8Ʀsӥ-p�{��0F�:1�l	-#���u��cN�"��H���-���.�B��M�=,���w�eOp��zMG�KS-��fa�1��	n�Ji�?/i���������%����4��R�3o��.�'���	_5 ��}hp�es��C���Ԧ���9���NEF=Pm��$E�͓)�U��P:M�u�WJ���ġv��^��(� �D]�I:�v��?p�ܔz[�L��	c�'`:��v�~�Ʃ���������`�ߏ�k��D%Is���q��� ���Ό���$����z��,o1i ���]R˫��J�7���n�#	��|d�*�0�h4�C��3����g_^"�6iئ�npj\�:���k� �ΰ����瑢&j�kl�z�⟮W�qp&�j�$���k�-9�l���d,E	{]Ճ�Ku�~�׼N#�2)��j��g	�c僼�E�z������2v��1%Nh�:6,3��
����ε����KQ~�+�ua�b�jƸ��-�����
����z�;���}}�l�c�L�Kg��5Y��_��`�\�~ҟ�~R�T\��!u%���՟�.�mGl[Gl�^��L�g&a�,�5�v�	H@��dH��'t��>�k{�ٌ#��h����t���h����d|6xW�W���xs/���q͞�&�.|����#�ن�c;?�h�P�t��KZ)>�i�Zm38��\y�t�X��F_@1-�`��%�`���t�=�ڞ���Uh���'����Q�/��2U����K��y�I_�<��-�I�Lt`Q-��85�7g��ڽo9���Ùd��G֦@r����"ĳYrj<�bcs��B����ެ!U�d������E���
�׳\J*�$��h�p8���T�>���)8�j̬� ��n^/)d#qҮ�R/Y��Pە��8^�;���	h~�=d��$ó���]�^��xp��i��m����a��4������O��b%z]��'+�7�5L�G,3c�d�Bsh�)34F�Ρ��,�%\�|�����%�WN�4>׈���\�'VUS�T��$��H���)3۞�<����e\���q�X�(��m�jp���0G�sf����fmy�{�8C^t��;��ϔh�_�/@�x�G\�Tn��z�P�����v_	����� yՙ7������sy�+�C~�ɹ�Zy�܉�5����f����Ķ*L��;5T�s��m�ݲ�c�7Z�]�����U�n
��!��NZ���u�������s��Pu,�n���W�w��&��(ӻ�!��(�!B��kB��~���ϩ)�!@����<�(%7�-{|DZi�5��_)��.�L����]�U%I�V� ��&hY��~-2���D�R�Z��Փ�Y}3�(��@�4��Y~��~>YO4�j%m{D����|��aò�t���~�DM�`�}̝���|D����Y�񩩆�+��h*	!?M)�wTwO�:_�&�uC���+�;a���bKe���8�V��E�x:r�E"�i�5�|�Hc`{M���=���>O�ք���gH�B�Ui�����F�h ��(�u�Q00����9d��ж`�C�ږ�]c4 �h���G��$ R٦�^�6#�{>%BN5�����$�	��=�|����@�xwe�E����I3_L2����!�k���V��� �A?B�g�ӻ�g�����idny�X�_,��6�Ry����āĝXq��T@���п|4-,��� 9T4
b��������c��py�H�թ8?0qqb)�K�t:ݸɑ����靶�R#Q�2N-��\�j�w�=���+z�(4{�o��[Eՙ����s ����]%S��
�����'a�ń�����p^�}A��̡\C{"/T^5��Ȏ������R�s��^9�<J���k𼗖8 ���d��T��n&j5;y�a��C����T<X\ޣ|s�t0�=��GЗ��XG]2 �r�TO�}�s-4�o�w�Cy��i���Yu�����/fΚ�n)-[���v
7
~�	}B�O�P-I0�p��=�q��K�i��zw��c���U�98?��%����b��zܺ���)�)+��;���b�B~�F�o�MNR�)jKF���X���l�tM�s��4)~�JR�%`<!61�A��*�0<�(a�{�rm��D�G��Ii��;�6�#vŵ����VA���T�s���u2w�o���lazB�3���m���۹\����B��~�%�ʬ�yѩ�<�U��� �9�tΟ�L:�Ɩ�/�L��4� ;"Jk�����X�nC�#��b;S�B4��~ޒlgr��8�c��\9@k�:�mv���cO��ٱ荽��ڔ���}'~�Jq���Ǌ`t3��'��`<��	a��l�U^Jg�T�߄>g�X��h�֞:(s��lD`!� �o����9������l��<�̯��4Z"���v�K�>et�61�ܺ^*���`p�X���0�+4Ի{G�����B��geY�����D
?L���9���#)�7$�p{��������9b�<S�=.?,Z w�*�@(������&��a�FהT6�xN{����۫���a��!��^J��O3@�������p�,vm�gW��#Y���9}C>�#��7��u���:�q�}��k)���L�9-H�""�b�P� �,�y�Ršu����Q]���=Lv�{�als�������1dm�{+W�k�7l�p��sI.dq[z��,�=r�����Ø5���{�稿��X���|�(wx �9օ�^vP1������4s���C3U�U��ק@�c���\�G1]1��bg������~��Q<��gz�Τ����h�]fWl�ǿ������
���3v%��GP�@�'�%�8/�c�����׊.����ٴ"�lP�����":z�Um�'�^s%���-�E��\)1$�W�Wa� IB3�u��=���R+���7���#���r�r���RL���G�z0����z��_�a�1ˇ5���p+� ����a��!9�3��ny��2l�������-M���8�wr�Z�����/_�8�q�1k���D��7���o�	6��7�^G �6�غ���͡�����)�/�#05劭���76t��8�r�{�[yK�&���"yL0yL��C˔���Se�����4���q������-�)�p�t>�gT���������%:I�u�7@2�"�+[�:�K,���5�@�?����?�j��_�(�5��4vL/��T*����J�+�Ar�˸��"и^��˼K)c���˼6�m��;�Ŷ1�p�����Y���tsJ���f��jTmj��Y���~��@m����)�a��3 3
��,Q�7K1��V9�8z!"Vb �B9��7��]�|{�r���~H��Ƿp�~}��O�Ͳ.��#�9���	f�wd�F��m���`�l`_(.%0Q �����tX�.ጀ)xep=~��"�������E�8]4�����)<Tޢ黒��,(>�X�W��髧�׷�l���d�/�4G���	����0�W�m'�|�o�7v��/~��5�7	�킡e�u#ֻg������tg��Ԗ���2���&Uq���'��q�&n���P!-]�7�O*��ۍ���V�ԏ�� ��G�|2��� �8�@[��F��7s�ce�&A@��~��L5�;v>;p	~%�C���DR�Sx�v����Pb�U��m�EԿ���^[맲�D8�v��5�y���4A.����
�A��g��X(��M�1�&�"0�s��4x�zN�W��l�>���?���Y���1v���sr�n[Z�N�T�'�nt��ۉ2"ڳݙC��VjѠ��е���wIz\��o��T%�A���I
Ȟ�Te��\o�-���}IH!���)�f(-�I�Yӊ=ޱ��_470�|aX>/��V@#&}��}%fh�ĥ�M{��fF��,�~�a��5����&�*�	bԆN�|�ҟDx���#U�n�����\P�{��Z�q�4�%��>1�B�%y@%�y�s�N� �p�O�e�t�"I��YP��YRP'����0�\磹\��8[d(,QmY`KYe��]L�!���� �1�"��%�����v��]@��իC �`jY����T�;�u�%���E�卤�Bn�Ru�������9%�}J=㬛�9����1���b��H��H�:4r�B��0cОj�KRQy��I�~/^����Rը�Tj����V�(�"V0dZ�UJ�o�5�٩en�>d�ƴ��/x��f8��{�=M?�)���½�NV�ؖ�ryV9�	��X����]�܊>P���˻��w5�~��޶�l&�#5�0�ju:nb�"�U8��#e��	a�ib]��&[�����`�#�c�	�h�{��L��5$Z�qOOߎ�G?V���G����Z $�N���^�g���G�P5�9�+���u.�vO�(#I:.L���:��*u5ھٵ��H��&���9���th������� ��&����_[�efFo��S�>,��?R�E#�>\	�ͭ"F#��W)1�#�!�2���v�C���a��p��������]D����+�1�{ܸ#�}6�kO(�Ʊ��1D�5*J�=�!;���[T�wD�Yh�B_B�2s����������Cwʔ!\��|�km=�Kp�+g�X߭Q���:W��4��L��tN�)o&�ݞ���`3-<��)��&�vd��f��8q����CA����[E�[{<1��M�g2Mu�o��-�`XD��b��ٞqUgh룈M��`|����I�m&^�N��	j����3=1���ؽU�z��;|�E\8,0��&�o0T���F��QpQd~���j�|�h)��a���V���~�~�0���J�Y�K��c��j2h���n�5={dLZ�B�r�0��[�������$Qڶ�pH��Xw0���h��r�D�1B���|���#L�?��&��`s�
�D�B2�KeV����d�I���H)�(u����r��[r�Vb!��ȱ�|���K���N�?����m�w`yQ&+�Q������X0�5S8j]wl���+U���R��W�>�R:�(j��RW�TεfZ���K-.�x�a����qDIs��V�
��.�������53�2����eX��r�u�koo���.{M2���ǻ�2����ȣ�I�'	�����"$0��L�{����c�Th������l����8-Iϯ��m0b2���="��D�'g��GjH;ھ����f�L���A,(nT���Ø��E��_�T���-��^���FLO�4�ҁ�7�����7h��L1�T�RT��u����[��"Fm=Vr����o�{��[#���6=E���F5�B�Y�~g4��r6� �E��Šr~md���?�Aˆ���"���T�g�S�w���m�A�ȱ��WW����A ��N2O5MF���uG����a�F:)���u��]�������.Rać#�C�����^��Cԍ%m��p��ށ㎑��:�o��S�c�G ���92!ly+��~��������.�A��}��ڟ����$�6����������.��^L�s�9�l�x����*�zd5g�\��k�cY���=�s &��fU\>{x��ې�Uձ��^�@X��X)������&�S�9h�t�@�F���lRM��</�p�T[��8�U��,�~O����^M�16�a���['�F�K;��\��`AGZN+^��N�=C��nA��az�&��K�y��to����3�1-�m�-��%�ʥ���`�͏��?���F�ǫ���5���%����Z���?�tfF�UvQ-΍55B��F�tҝ ;�Cw�Ix�Ur�񭗒���'H�:�^v< �-��P�raw�D������G�BX�������M��?`�^f	#�Ib�:d�+�w�
��$(�l�B9��}QF$p�8(�;���������ߩ9-�ǣ�4/ZC�����f������Ae�%qy5\�7�Qp�W��Ml���@	�4�2����M$��nU�!WH��⧋+��g�U��C�y�m�B�_z�C�,è�c;�3���A�vPe�A' ��{�B�q��3>	|Im��c'��r���E�9�Hy�W�]lW�T�%�e�z8�rU���Ԟ��*�n4�S����`�
�Bv�M2r�V�<�Ga��>��}���_Ş����[����1j�"�?�����x��5=E�$8�v������N��1}d�gQ�&���K�&�r�J�b���rGx����C���u��ÞV�ü,��R�(
�D�)����P���L��k�o�����W6�gO�w��x;��K�n\�m��E����X}��K"a�گjT�c�B� u��n-WM�8fg�0���xM����-6�k�ZԮ�p�!���?5����1~���p���%P��9t����uJ$Ii1f&ϣ}��yS�Ƃ������'�Ӣ���!q��{)ʖlu�� �ء�"`�05s),y��`?�L�C�I�����ަ���>d�ah{R�l' `T�`q��,k��g1��0�t(`
J,Ut�	|�\��e�Ե��5_�E{	��d��_�SL{=o:��_��s��������1�P0��t�����R"����;Jf�@R<KHte��fH���(�Kl��ҝ�O�
=�1tl�/����_ù�����%��Z?��M&e7��KH����Ӽj�-g��+`�u�.�Qk_�9��Ԣli�ɡ���uD��VjTaQ�Ʀ�-^���h&Ҧ�1I�	7�e��W��䑖�:�tFn��ب7�yL��*�<G5�� =��h�5�9D�5G�}$2�ƕO�	Q�л_U��Y��K ~1��m݃�}��
MT/]g�� �i:ۅ �{�lT��3dCȸ*~�P�T����%���5��Z��"C�4���Rk���We,���.�� Sa%�A������-��Cs��N~#�n�~#C���+ѝ���4�w>K�>����Ui{_�f�!��)̋'�����(	z�jv��c��Z�v R�TE^�y����ѽ\͔2�E�Dx���|W�v��5ԑ���>�U)Oo��mK�ʀ�ؤ4UI�Q��~"��CA7�^AЀ^�t���!J�|��ij��d*Q\�����w�n�-�J�MV��0�30��&�.��ՒB�v���4�����V4�kdl�|�(RĚ�8b��}CO�<j6s�E����'*�=�'G���z\��h������&�_H��P7D��
��i�id:���ځ����VV��i�9��ךW
3Է�>q�1v��r� �(���=�o�v�N�a����6�a�I��H�2�zP{��\ ���o���LŋN����Auvؾԙ ;���H�ʻv��d��9&��?��r�5I�t���&G?�>��3f��(R���r�Z�1��`+�o)Y5i���D�� ����Tܓ��g��{I���Mٻ�����E���V��_F��.)�xn	D
9s�?�
�
l��2?����^i��3FY>��#�t	y�g���@��G@]?_B�L��X�

C�{��<%<��n���࡜�EZ;�.���@�#(�۳��0V%�_s��W��=2\�
ȭ�|����(�]crZ�[ޮFr���Z�H�b@
.R�[/�� b��T����9֓Ѹ���b�2�uT�+�N��Q����܋S\��Xh�w�'� "���Cը;�&oW�����/�wr��~b���<5�8�PңR�Ӑ���P/��L�Z�����ᕖ��7��jJOS��I�
����%�4����ם��a�:�C��"�g���F�30�!��T�Nr�y��g5jw]�_Wf��Q���Q>�>�*xm�������nV�П���%Vy���
�
�"�_�J(��߬�פ�f����T��9���J�P���!� ^��_[��6���9��}�] ��h��++���N�sj����e]<�I�G�ó7�B�����|�5Q:<O�0E��y�v�%D˲�:ۏ_�Q��{�T�b�{n����X)����&�Ar���)u�U�g��.��H�����Y9�E:��i���:�_挀�SO@��(���v��U �5P7��ػ�1G�y�-��}�}]͢��L�3�XV�
���I�v1����t�� �R�yi$�5�z�����-&O�]e�eycEx���N�T��v��Z)(�&�P�(��Y�h�^�ʷ$��Ќ��i!�����]�Q{�z�*�h�z�f��6u(H�J~��DNt z�2>�7�WW1\�L�g$=%����ۤ��N6�)ծ \/�-���7$�y�"3��]��WNX�(ЈjȎ�f�6�6F�@�ܣ�02G��g�Q�n�C�7R�����#�#��QN
�:;�8Λ�ئ�0��]C�^]rS�Z�푿�2�?����q��v�&v_���u�{L>n��b*5lC�'ϒz�̲���V��x�.���(V<7��~�m���/�Y%�s։�?���l=UA�itO�����4p�n�ٗ�7��Vԇ�\�n�&�M��a����
�G��h�5Č�U:�a��w�/������Y2�5�H�gj�\գ�ףNf���̸��/�4m���������@4��|&�̦x��,�%�Mv�u����P���t�+.�Ȗ�FtZl�򘼤F1l����*-��*�I�t�y�r
����}!�&!N���Q�=���y�]�%|���m���W�s<�bM��m�߲�:�%���K(ߊ���적�Y�t��� G�C��ڟ�n�|�e�$�2.d��c:Xij3��&<a���@L�;7
���P�p	��ȣ���q&�����$�����9p]��27�y4�To�i�풹k%�x�������%2f^�7��+m����FX���G0��>��׹�m��:�ť�^�hx�jV8�9
�F8h&��ӰVf�s߃���k:�-tK�X�6	�0i������nN���`�jb3c�^�AK�Z�Ư�o�f���5�u��ā	��^�_���Zf�Ik憞�Z���?�����������댜�DT�d~������8?��s9z�	r&5A�����&�hg�h����F�<r9W/r�����{b2��6B�G��ݐ���-I뀭˾���'9eb����Zg.����������j�.ߘ����HU [����,�\F��KD�h�a	�-���`�Z�2]_�<�3>������<n��3�]{dsO�Ԑ� ̸�����[W�	!w�(��I�l���m�O���,�ĉ$���;aż5P���zG��I�����]E�e�|l�w*u*��)I��ݯB�����.�|�		�C���]R�쟛�<RXB���Z��R��Rҿ�3R�@|�40�Uҭv�Qn��$�f�p\�a�%G�H�]�h������L��(:0�Z7���X��oF�1a}k��;Y��x���[�v"��|�3�v� Z��0ak��]�E��=,I�W�T�L��4M@sh���zp��@ł%�����ڔ�1�q�r,G2H��`՛DF��RI� ֝d �ް��{ߧ!��ǈ��+	�m������G/T�OC
����J�Cg���E�tʟyЌ@P���������0��.������x6���3u��ȫ�T1<Wx����zǐ&Ǡ�UpQ 2l�eC��։��ܒ�-7�]	/�RN��7�&�>��|攩!)M��XCg����H�֟��B���u��JWv ���bH;��A�uC�z��[��er�Fi�Ր+��F�tZ�4�x����,\��`�z�:-���þ!���/".��{����0�&j-��-��\����	jmS��I#9x���ϼ�'�b�C��;�zg������sf&MS����[�����NeQ{�xg"-��
�ŉ��p&}M��%R0�n	�!����@������!x M�6����9�B	A2ު�3h�ܲ��V=}h�;<��Ziy"-SlWL5}�;���/����8Zg�VE��2!D�1*�B8/��o(_h��M���A� �'��Z������*$��"K4mn��ɣ>x�܃�v�+�b�#?���d�C� �N�B䖓�.�z C��% Յ%�aHD��Q��4�1<Lt��e_v�)�o'�<8�>����~$π!�F�	��î����~�r���4@�,��6h�?�\�N��ͪЗ�?�q.���=�⒩���I5������]+�<�o&q�{S�
,��T��y���u�ȉ�+Ka��|n{���2��UA!��j�#fH��� L-�̴ X��%q�+�w1��r���	�����t�-����ܡ�E8uJ��,���Ly�� :�6#�=*����,!��pS�C!$E����vm�WC$qp��~[����P���3+ŏBZzٮ*�,�c�Vʰwh17��W��8��p�J��n�ʘ�p(W��c!���Q��&.����J�f}�
�%=3�yN�v��4G39x�Qf!��u��%;���u���>���� ��q�3��| %zH�hj2�̝;Kx��VA���gCGHЈF���:t����2�O�������:�iH�/�.5�Eq��3�Y4���'��F�'�>x6�Z��/2	O�]�9���7��p��ځ���s��D�N��5L5)!
6���ɩ�{v���B�^�)0Af��_�B�h�`�r�&T!Ehd�����JL6�"�V�֪ �a'ս����37!�+�tm��&��M9xv�K �K� ?55?CL�9ʶ��/�P���7C���Qg N�=���UU�I���p�<~B��2�V���Y'/��O	���y��(l���B�(7�5����#: -�}*J�s��� \WxzprS3�\�����n�y���X��l]oM$�l�� ���$�O�اdw�u`l˝u�i�A���x�o�-Wdi��L����>�+���$���H�2�7SX�b�_?�c��0�a�}S��"u�,��{�{�����F")B�P���������]�4�����Lx�`� 2�նȧ"6Dm��Z֍K�
u�0%<q}�tt¾���,X[����y�e@����U��4-�c�u�p��	��N���!Q�P����m��n\����b:�l)\�3�@s��'o��O�w��_ ����PoڡP��a�eۨ8���������wʯ�>����r}�����<�]���Yr�+"aMNj��Yzq���ji��g ���"�_f%�)s� �����H�q����?w�:���F���E���T���mB�7��Ck ��z���|9rO��1}D�E9n?S��x9�f&O ٮ0��0�/h�]�Ň�,��<�F1"]�-���|�I��^Q�w^��I��V8͂��%#�yܵ"���"�[�ߕ"bFD\ ��o4�M�g�U3��F�����ҽ���2&{:�%'W�uTJ���>�6���^Ñ�Mk@��Jv:�W�r�����4j9߇*v��<�
oO�B�{,�9����*�y r	�3�Az�@RG��Y�����Yp;��ζX��o�� ��͢����V�_>a6�*��o�k�=D�h�Rt�';��$-~���ib�i'�/�����t��z�>�#o�Y	���O5����D>�Ƭ���5}�������k[!���vv��o��22jys�K�>��?�̸�;N�{�;ͳPH�H\�
K�t ��6L*��":�Mj�nJ�����?t:�׺��4��!��Hr�oʵ�>��$1��I+p��=<�lo��a�9.;�;��z
���}E��X�Kt����QF���ܖ��۶�Hʾ�E�K�y����`ӗ}?�h����q��Ļ��K��˾i*������芒GKy��!?�L)�T�#m��ظ�Ѵ�p ^���p,��P�6���b�q�]�B�iqPqhSi"��0��w��C_'k����q�Y���c
�8o��$�q�^ �hL#-�6_�
�֫�f�$���Tl����+j#i���ji�M��N�Ϭ�O ۟��k�Y�(�&r�iUD*ۑ>��4�Nw(�
��(��OU��1  @n���l��w�Q���(��,�3���K���^a4s��珥w�s��	�,63�C��A5��J���w3���悅S$�P�}���ϗ�AV�ԯ�h�.�[���H��ޔ� ۅgiD%�0�C����1�|�-O$ �N,��6�6�#P5X��Hz�PU��-�	�(\L�U������Ha�|�Oj��lY �%��c�.���H��}�Ӣ����)�y��a���9���.AyF�5��_-��n���T߂�KE������b+r
X��g� �!����l�S�a�N�FK-��iR6��N����j*i�\m��L�e�a?Ze��kϘږ5�b��k�1ZA����S������5�ԑwiE� ����-Rhc�������?b��KudݸU�_���^�@������{��3A�}�2������7E���w��=�X.� n/���w�½�P7w7S۴
�X�aZ�h�g�u�ʓ��IU��U���/LA i���AwB�N群��h`q�T��{�6�§�o}K�BkRnѪ�7��i�T�g"�Z'D�"p&e�}�mG�g�{�P��ҫ�	椌�!sw��	&v= "���/��6�-�w�;��zo9؆�����N� "����ȱ��Av���uF-����܂z�cĦRV�k���j����$�3P|���<���N�f���'��"�<+*{l���_.w����%�]�F�	�f�c.~z�ɚ����]��?,�K���Bn6�Fr6P􍋜Vn/�_�cQ"Z������% �k�J,tj��8���r�'�=���\yčEu#�&)qn�p
��.k���& R�!@�|�J�#d��������8��,�����i'���;���b/ K���;�X>[.4[�N��F
�Z9�ҭ���҃A��U�Z< _���{@�������.���	
��"BE��t�oHb�`��o�{�t�1�ef{]͵�&1f{�.e?'���k�������{0�XW��V˔#��q%LA��R�3����� 4)�(�h"�0��3-u�N5as�+ƀ����h�븥�5
�,EpʱI����P�B8�Ê"L��l1]�����q��Jc�77+_�b_6��?��Y�p�/%ﮑ���uo>y4`Mﰾnt��`�����c-�GS�y;B!-��8��C����X~m�ʟW\�;֔ ��.�	��H������Ƶ��W��ӢV�$�J�g�i	2�	�j�,'��K���*��+��W�aΊb������_���59�t!?�
	�!��F���h�N �٬�<�,,i���܈��b	��wݦ�N�u3;�#��p�֗C���`�	�Z������!����_���a�]o�j�},S�̴����_\*���Z1� 
W�}-�+<����0�Ei��5�}��Q�aK�?�^�|ǣ�;��`|dl+v��V�m��@��;�@U_0�4���$4�zv�E-C�R-��?���hb�,`!IY�N�33�;����܈\����ήi�{��N_n,w0��t
���8��*���ިqN�?�$?P#��+��$+�M���H�1��Y�ߤxwl��2�KOޑ�����O�&�a��b����=B<��G;I$o!���7�D��im]�Pi�U��K��k%޼����t�����{ʕ��/���(���<����4-[��b�X�GV�B�G�W��J�Ay.IՑ����s��ג�U���&i����j�k�h�$az9y�ze���q�~����+��B�69J����������/�,wp$�|�w3u�w^��:W�!�#U�t�`9��)=�R�^�@�Ԯ�h����O������h�PJ�������I�����)s�w|��㟞#NnZ���2�������MS�����9slR��'̠��'�;�ɒ����x]س�7�j�ѧ�O6��|��`6�� Ȑ�}�+ߟx��u1�[�"s��"_l���J��0�Ͳ�v�D�Q�9�_���	���>q%G^[u����њ�Yx�-G��UQ1��"3�
aelԩ]��U�of���Z���D���aUu㭍Ҩ,�fs�SITJ:5�`1sLƞ��8��A�������W܆��i<1�>s�����'��\*�!��/���&�_���Yz�9o&)'����4�� ;�d*���sB�s�5��'Zv{�Xѽ��D�c��<!'}��S����@;>�d�䳥sR�x��-<h�D���q�^�)	p��C��W)ڐU�bO8��m�a�m��W �c�P��-	��a��7��}�M*��=�9�2�a&=F�q�,V{Dߚo@�[��M��	�:캌/|?��}�3*g�UrZ<��)�6�#5�MFw�("ҳ =�����rE)���_dÉ��>�GT������U��'uM8���Π��� q��ú_~�Wl_dE�=�O���n����>�F�3��E�y*|�6��ҹ9�t���O���$�r�שn}X��}���liĵײ�
o���H
��J���Ijh�n��O��mp���J���;���d)��a�#{�L�n���R�-���$���,z�ܿ�*��A)��bi?+��LyPyz��N����v��ǯ6j8�DL}�-a��ɠ1�
���P��Qk�ܙ��?���$U}H鍂�7U��'�Ėi���c$�k� }uz��44�A^���1̐�i�^i/x���(C�2Z���N�_�$b���u���I[V{ƦTc��щІyQC	��oZ���|��J3�7a��~��",���q�Q�O�B�@@%��pl��1�[��Y�Ģ4b\ކ돬6s��>ڳ��Lf7��_�^��-���K��o�\uJj��G�(�T��ᶶ 0�X�����SDZ��욅0[@Ž��27z���oL�Q�|u��� ���y��1�.W˰��=w����IQDE��4jL:�@�k���D��)ȴ��~�9�;Ic��P���w�;��}�tŁnrv�A�P0Mǧ�Q���T6YL�U�G9��gTƑ�#�S@~G��@���g��Ҿ%�z���~��❪	*]i��\˩ �_sw㞹��	E�$�_ب#�HgƋ�\���ޔӴY�=~���p�tLv��-V��ƾ����s��xM��K�rZ�S@�x�-mK9v������'�����h�͔�U����)W�m�b�L��~����K�"��j�=D9A�#-'�*p���.��O��M��acG⡄�ސ���'���-D]��>�&U����8#���{a+H��r/P�J�\��OR����-���Y.y=����>6��=L?�C��p<��V�z�<�b�!O�ߥ���~x{5�|��{/��"��Q=�4�B�(�uzk)j�'MR� �A��>L��$��
��?#q.�,0*���� JJ{�i̼�0��ڝ��Wi+)r��iʶ��c�������i8h�p��ϙ�1������rڐ�)�­�.H#�h��k&d9���9ep�![10E�c,�R�u��(Z��q:v�@\m���;d����H��e�P���k��^Y<D�Ϋv�ږ��La�7���1z�m�,0��I���l��(,��gU4�������Ԅ*r��P���zy�;o�Ft�*�fd��x��3����~�H�-�F��l�C�#"@�_�Ce����ɂ�(1��0����a#�H���t����j���ł3���4��"笼�Q }��/=����3�*�-A��j �J�G�)Y�
'�+�(�P�u�K��*��W�H�:O�}���Y
u|�H�Pt��r`<�y���Ok�r�n�OX���q����A�[_NpЖ�㊢�t��h-Ⱦ����q�>6h��/o�o����-ڏ�}�/*|XM[+�.̱ɭ�u��n}�r�~�$���K�^�4�i�O��x��OUc�e�dݯD���@kI���o4�}"�a�g�&e�҇���7z�xJ0#/?%��u^����C*����&ɍjƚ29��7��}��p��Oe-������=�͎�2�A4Si+�	]�U���ư��e�-]F��E�5Z�#z�� ��z��il�W�*���eD��$<�d/�
C][):���j�=�?�
j�H�E���~+�깾�G���+q{hD?���v4�z=I��x��%�a �Mv�Z�T��ߖ3K���;�8�ր��Hڰ����.W�{�κW�IV����8���Î�RJ���(0z8����x��J�"� 
�ҕ�]��nEO)<���Z��1�+�Z���I���rxC�������&7���^���M<:�}�"Ч��Ǳ���?q�v����ͧ��Ï'X�O���
+��/�L L���Q)%���ǁ���.����#��.y'���}��凜�5ҿ%�S�R9��*���(���`��Àa'$��|=S՜�̶i��Z�����şB��w��1)tԎ�-���Q�l����&L+�_�� 1ݍ�t�iܖ;L�)�{�JEm:� I��#
5����ؚ�%�3�]�?�|�1��Xja1���_8�鰑A� �B�f�=�՟Ġ�$5�ܭ��6���X�$39��g����]ׅ�:� ��gƄ!����)I��I�2ym�j�_��1�^9q�j"�m((�9�JO<7@t���^<mVt_q�DM��x��X?�b.�t�
3rTȞ7��WE��[ی�m���%Q�9��u�A݌P�W�z�]��4!W��$�?��BJ��{޸�2֌9��{т?r�V8�����Z�eXsW�p뷃���(%rś��3'c�F*˓ȭA�����<ye:�/�c�pf�/�N��~JZ� s�݉H������+B\��GB�n�5짧W>tϖ��n�+�v��[ve�/B�$��1�R��i��S�.,�>�0 Q�/v�`<3���m��������q4���9D�w�鶼�Uɉ��"�D��^Xr� Â��|��@pf���{�i�5� Lrz�-� |�*�8Ԇ�ƳX�3$�s�� :G{ˮ1-*��=��_�����k�����>�T��D����k�	��Ի���g�G���439�*b-EQ����{��t]�<I��6U��2�"����G8^&bʛW�n ��'̄���̦�Ƥ.V�),w!����q��`�(���[�%�_���|m���&�a�8��S���P6k�� �z�Mu�Ə�(o���������p%��_�<p"�u�d���W�c.tj�ݜW��N��ɘ�ҫ��i�@<�����|Y�h"�P�H#zL}�B�nm̚D��֞T	��\�U��&,�"v��G���@7�����>�U�/�|oҭ�AM#��Q{��E��%G��U2�H��VJ餣��j� �x'U�Pq�@�9O�
�$%�A���C񥾪c�O�d	�P*�YӸ$.nO@��$��s�ך��~�mw���a�E �y����wTMU���XH#d�V6au`����M���!����pg �F�R,���� ���.��*�GF�0����D����u�	�N^qW�p��	��9,�Ԝ�1�5�g�a�E��=�iZ�wcK�aHI͎j���rBV��0<?�X��?#=X,�� `�� O�l�EUT�����U��w��.��>N6��j�-^�y��[V�1����օ��_/�Es�H��p�
4m��V�J=�޵�3��.%�G�}�F�@G���z$*E�|XZ�Z��2��'nBc�g��7��,���e�,n#��Ss��Q��4a�6�X���-��e��h�5�2ث�8k�>�Z�IGN�݉1��`w+h>x��H�5$�|l�����@��PR�َ�a����I3mWR�h��,f�̞�XRb;�V�6�����ҸИ"M����?��������~���q#�����Bї"T�7�eL�:x�b�oN�H�Ry�/�D��w�;�7�-�n�O�5ZkM�f�c+m8)җR���\��x�Mv��&A���:99Z�����%�.)�'[���վ��k��(���h�'�l�7�>�g�c�א�΃�e,���= Ͼ&��]�P	˹�{�)��銖�t���WԬ�r����Hܾ�#�]+����2Bo�=��p� j�bN��xBj˭j(��f�i}+�S�l����굧��H3�MKA��r�#��5"e�E��;T2�.�n�tP�<p�?R�I���.֚��S��"�Y:ܔ�"%�dD;d���,��I����Cm �o��u����R&�|���ou��`���)��M:?
��d��-hJ�h�}���Q����$��=x��+h��RJ1H���m T�n��3rJ �I��Z�Ը7m��{5�6�W=�9�?^do���qި��﹟S��q+m/v��-��M�Z�G��7Ş�{��^Jj@����f��qD��P�O��r�vt�9<~��k?�p���F���{���2��>&��[��I�%�J�tH�ͲlE~�a,qh�����Z��䰁�v]�o��7܌�����M���������ebF�D�ܛ\��G���]��W�d쵮��c�������j5p���."_�I�N�Թ#�d���gd�	,�oO��:מ CHy� f��佅n0���ۣ�z���"S�u��<�b�	v��mt���11�e�(��۸�FQ�����/v�`�/`s�	�����/#:���8�Q�r��q ���l���z� ��&�����p���E''f�=գ�g�������Z�Hy�D9v��ݽ��V��d6p��l-�
�rA�s��ʮU	*;�&�S���NҊ�jخBӏT;�w��4��B�J�'WdO+�k�MB�w�.���6��A��ɛ,`H�\#�8����J��ȝ=f5��;��3٢f���]�� @�O�����.9�R�H�ӭ ��ߵ�x�R��9xsj�9���"DI6���1Hc����\���Laj����1�k�*����>ic�~$@o��y���z�=��ƈ��,K`�/�ǹ�A)���I�}N����69ő�j;(��~ �������U4�י<RQ,��7˓�C6ظj����������ҝ�s��D���bb{�x_����*���=yK/5l����$���)�[�����F���)>o��În���[�ȞT���e��N4��+��Hr�rK ㏐���4��S'���R���A���_�u�vB|2Hm�`@����"�&�ͭ�S0�x�38�x���텷��|�LO����z+y��gmNx9�j1^L�u�.��T|�n��az�"t*r6�o��'u� !�V�kv�NEń�6AW�Y�	$�K���]�8�[H~I��"��~�1�R';�-;󴊜VAԬ��	H�w���6)J,�s��2!���bǭhьB	U��[�9H*��������irh`��`c1�	�����B��>����;([Q��5�wϨ���LߖN��0y��$�̔a����u'Ф��X�b�EM���~S�nE�F(��L�ҍ�vY`��iI<�玈;�����l���e��B�،	y�c�|�>������k7��JWs�㛐���&��mzM�U ��w ���1E�=�VV�Z�C��H/������ٛ��ԯu��R�f�DJ��ӍLY�Ԯ�4�:L��i:13	z����S�\�DVpՍ]}�q!���ad˨��m8�e��5g�j	d�Z[���{��۷���kv��b�U�mp�A՛�q*$_��"e�Ec���A��������أ3_�*���� r���Og
_�<�Шfb�d�3E���VP����B����g_�k����j��|ز��S԰B�&\�t�O|�Q4�vc�P���%�h!]�ө�Y�Bf+����6�=��g� I���# ,z���T��&ھ
���G�����ܭ8�Q!0:0Ē�n�8�{�s '����"��?���v���B��j��~�X��d�!�^o7�=�sUw/�0���>E$�Va_~�p�NeFL�O��e�C�)\y�������M�rn�CJF�F���;�6�����/��o��&Z �P�+���#���(���7�8w<nME���c"�cOܹ44��S�5[�t"(�MM�$��Im�Z�������p��t�:L��'�	Lt�^)�����(�)��zlzi�������YЉ6_���G��E̫�@�؆HT�_ �b��6��y�R:�}�%O+���,C���u{}���$�4-H���v <�v���IZ�	i��������ϥ���e����'Z�����5������WU��<!�CyQ sH,�cݷ����q��#D"� %�U�W�1�l�*(M�MaXZί�"�yG�ϙ.I|�����S:��5�{5.-́�s%��v��"���cJ��$�j�_�6�3Rd�gU�$Xyͨp�r\�!��%30bZ3�ڋ��}�[���K;����g��!��=�x�Z��Ĳ�"Q�G$�KFe�ޏ��)*t�����K�P&n ��֫���Ea\1��\
�(nb��:6ޘ����p�RC�YH���v�&�&<h��o	h։W.8�Q�
��	IT*�W�68�:8"#ȀjJH����ЛX)�L�#��-m̟�x�,�t 2����%��#�m�?���ۑz��G���6 ��taa����ݳ-��&OTH���[��S8_�ӕ�K�^��UQ���'��#��X�8�׀�0�;]v "��#���|�����Ü �DTQ�8�9u=k��ľ��E�.�#�Ѡ�Wm]n,�M���xv�^���B'K��c��YV~%�1R�P?���g�P-7V���u�J�ѳ��΢�����s�G���;�����x��Y��x�� ��r��kRn;C!��ރ��د��:ے�Xp���E9e�l�p%��>���ߊh��}%Re�d�X`��D���<�.Ȕh����J�z�Doy��l�LY��<J�\�|������5nbk�$���v��(o�L�QRnO�}cd����Cܤ����:ˤ��C���E7����:�&A�R>πE|[�m��M?��/n�&P�����eo&+cR�mFJ�����Aݹ�6���K�!B��B��D#�����Kh]ض�ɯ\v��)y_ac�����dU�}c+b��]���M�R !֩����;z�(
�*���ư�
���w����d.P(�*v�ТY<ZW�.��ɠ�:��q4����S�����1U[����,	�U�"��^����W@�+��S9���$�H���.44*M�C�8������ z�Ɗ����ǁv$?5DS���_�H`"�30UU֝�ȼ
R���Ѵ��-�dR��tw�A������@,B�q,9[�aF���g).�ǌ�#�;�����O��|v`{ZM5����L�.ZN��iǚ�]�0�����rÇl2.�KWW�UqO��A�!��8�p<���K�y��A��<b�|Jf	��(����"5��=E��~0�<"v~�OUu�F���L&¨���O }꒪��6�N鋹C���X`՚섿vs3��s7X��I�Z�C�mm'T�5��A�S}�b�nb����K}[7:(����ύ8c��e]�&��q�O�$�I�et=Hl�,o�B�g�AmGuт'��M���# hD^^�Qx2�+V��F\X���۱��ﻐ/u�(H:)̕�J8ѓ*ɕӮ�.jR������������B��Z��t��Y�:�ZX,�,���L-tBYf�%����nN@@�`�Aޅ�	x
�c��J`�+{�t���DZ*m��}D�zS瀚���9`UC9�ߎK����$l�u���ܥl�p�G�I��yI�ǒY�l����
�ż"����j;qdR�yI��wŹ��a�r��`�#� ���օ�}&�2�1�6�80dә���\���4�s,�k�����9��*^���/��Bs�A>*٠e{�\���V���[�Û���J'�,�5s�g~��������(1�i��+�
f���lCpX��;�-�?�+�7/�1å3��[�|�p���t\���#���a�r�DTH�G���MM�ba>�@�*o
|��"~��+}KĀ'lƫ�y��훿�/���<|���H�2�E���.�c����U�s>�P'��R�rB�
�DVޓu�����������!�ĜNtL.US����n�3a2���w��9B�o�X������):�=m{Y��g�_��`�;���:��k)E�\��e�e�eĞ*�lP��qW����4V�;ޠ[<�Q�K�K��G�YCC�2���qSt��N�"�t��u��kG��)���"��y�z
��u�������BĽ0��v�_w�����e�e��DC�'E�8��C��X{�) ��y��_@�n��ʝ9o5#Q`[�8k��g7��u5! ~~Я�� ��/�+C��)ڋO���(�2�K.(��15�J�ſ��C�:j�+>�bW�!�u��K$l��,�t=��:�)��;��߈����|	�Dz�ꃨxk*֝1�4��\d�#�Es�Mw3�o�\�wpR-��gR�Ħ㪠Ta�_�)������I4�-�ٹ��B��x�	5�?���f�:�+Z���j�#uQ/{ҥ��@p,?��=�2�@��7�����7F�Gh0\Z5)^�֕�$:��+K�Ţ��?����͊�q�U�Mr���;��8���������I�G#�0�uJ��9dͩ���=�O�&��"fZ񿚷�_�ō
fW�gk�R�-�,�||���Jy't��5��S׼�uK\/~k	�|rIt�i��,�An��'?�n�ٺ5�_�s�"�v �b��M*>	i���p�jN���ts��ǵ*��u)�l�L i�|����ڌn���"�+���6� ̙٥`�Dk��9�ډ;�����"��`t��U�J!�Ak��h4\�N�3��#�t��kyq9bOU�ޱ�7�L���W��*�m�D��z3'�F�����GD�(]��r������Jp\ܾ�!u\�'^H ���F�a�uW).9���	#��)A�Y��.!
A�xE[h���6�����yq���l=�V�d!Kj����7��	Oô��x�'��u�2_�]�l�h�a�W�q��T�2�4O�a<��u�M��ywd�@���x�ԏ��s���q�����(=�vN�H/��נ%�G�b���2��i���/�C�)J~�g�R@F�cD4=C���l��d�/I�$@X�Q�"s�w|uDKxV��{�Am�U<�P��1י�=�<�x���ȡ�� ����(�a��
���%�P	��0O�-#��w�O�$"}�{�6�v;�U@=�T��kc��%�ڣ�� O�_2�r�x�,q���)�����أȠ��T�/�\#��G^�T�~����r��U�n�PrA�S��2c�����Y����MU��x"%���Q1��-E^v�N�z&��l�)�#��=݅U�\����2���t�C�Ǩ�L`�?��+<���#/�(T���z���L�Wf��V%>�!�vv�T�ڒ�(o���g<j�������[d�J+�tZs$�'梓t����~���q��++jY�4����U�>9V�13���<1��)�p2�@4�*ۦ�@#��O�� ��u_�;\��2Q�	��ַR��C�H��@�])`|��n��\������Ē�L<X��W�u�� �	s���j�A���d���%t  0�
X-�xQ=W�)�e���D��3>I�@r�l�΅'��K�h��&��>\T�ǒ`�V�%��I��N8��ѢZ}��	Cӹ'ћ!(�����I��0��ۉ����(���4YX
8괂��Y�(D ��	;����8��������[���_�+�и���xT'r��u�dk��,��w�(`�-���B�o����^�N���?�g�d$@c�d���B�vN�[���K)�⵴U�����oݾ��Q5���2�p|�{��)�Z��4���t�0��(	�k��&� ��,�i�s�dΩ-��5������o蔿x��fq��\����{�o�����m�E�C����n~�R����$��-$�k�����KZ%k� �NbN��@�0��Iы-�������p|t������:#ͣ���73��5�ݼ��-C��Q���oY[U��-ɓ̥��d�5��G�4�"�=��)��z4jJa5�5�+���U�V�G�C���o�'kE,i����ex\,�	=u/�ń4��ǳ����yv-� �-�A�Jh��] (:�F�@.�u�v�gu�b����P�lx(�g'|�)����{vѐ��K
QT����O5��(�ߵ�C+[�\���g�� gE�	�b�lV&���0���8�|�,o��\3���Gw�DI���f3�������mm�Wњfgm
U��)ǭv-�?�Ds�~��f�Rh��C��y��8�l��	����jϯ)��!G�bSG��^N�v��%$�~�=�O(��d���bz'���ص�(O��
1G^�m�Z�����[�u��W������R	}8+�q�:|n
��.�|D!X���Ý�vA�5Pn=�4C݅���p�7��m��5���\��x�k1�-�[�c
&���g�p!�nŞ$o��.��-�[��1����X{�a�Bp�,��Z���� �ɠ|�@~Y���0�m��X8�V%�(�t֗>�<�ܯN6��M:�������9r�BT/�<J&ioo*Ŏ��ˋj���3�����'�0a
�Ϧ|���)?eV+A����q�������C��{�ƪc��fM�ǂ�OzXD�ci?c�&PD9 �V�TMǿ�5�����`�t�������$�M�J���HNe�0C�u��.�5z�V)=B�?�G�����7/���3��\���y��a��M2�_Q�i�g��sm	Ϣ�
���K�@O�����[\`�����9?�Lݔ�؄@4{Iˠ":�]���%vL�&�f��fHf���1�8Xj5ei��F�T�7�Z�#�mA5�tqn�=�g�Tƫ�u�i͉9�']�>>�^ ��x��1��*����?�њxI��i )LF�@_ ��o"�5�\�D�T|�)�b��u!V=���cQv���D#�HZ�I߱�/ �*��Rk�����Fč �C����t�I��:N�����#h3�ڃ~΂�����{�gmI��2�p�*-5�gD�{��8����Ol��QH.ߞB����,K��=�-�#1�M�޳f��@���Or��I9)�H1��Շ�i�T��ئMV�HB�u�?,Ƹ�s������*�vj�,������2�C4$����8r}�`N��f��Ɲ` q�-�j�@c��*�!�/o�>T�����w�ECinG05 �89I H���D���X�[��8����RA��YZm�|�D�$EE�I4΍�dǾ{�0�^�PSՓ��n>,EM��)�_)[=���=&L�3C�o�0Ӥ��k��Dïg ҫݮk��(���M�	���~��/:"�O/:3#���݂p�F.Z���^W���hEJ���#���>�M��jJ�5�.�DQ��<t������O^t����O�t�!�ss���`V賂"��=;�q��,���p��m��h@́���4����<a�*���~\�x�D��X@Fr8�_-H�x��i� (I�4��J�Vw�cC�����K��"V<P������.ʌ��=��l�"o�'��un��z)B�	�B�3>Q�q��h��o^K�+�1$%��<���*.̲��H!�����L�vB:C��f��1�h��5?���=���I�g�Uf�m(��(��겛P!���~�E���;�M���#���dgɽ��#9g��Ǩ�c���

7s8OP^���bO�[�8mN9B`�������(�n�@�H�� ��E`�iΪc@0p�s�)}��'�C���D8kKZj.������9�Jj��]@��m��x\�N�(�Y<�������k���	����G3f����6Yv1̻��G��4���4=4��ę�5WSN��F6v�eӭ2�� ���8���c8� r�m5��1��v�!�E2L�����z��YFLF�*%�W��Ao����vͥ/]��!���HX�"`�?���Svϛ���]ސ�<R����$^1b��}�S���Ʉa���[AA����-��h�; |��*L���M�'�K_��8	B4�e$7C�c&����5�\8>L;�j�!F�HlQਦ� E�W\��@�����ìa��e��2��"��#[�5;g$%S�^�#�)�*Y�}��|&�޾�����X;t���'�km�>�P��Ҙ�IVGn3����@�
�P��3�x�`�y�����)]��:�����B���,�R�1,D��]���<cf���F��gX��
����8}۷��c��v�e�w-1h�`��&q�#p�8V��6�*��Ճ�g���=N��z��
��ݷ��H��9x�T�&f��Q�͙ �}��E���O���!ѷ�/Z��X��ˡ��{���O�>P%�I:�\wn�
��I�,�q����(b̈́g�k)���w-�:��ꃊ;Iz�᭞E�/B=M�ַqcY��SJ@��9_���OG���a`�"�J&Mp/��xŝ
]�?2�M��l;ga6��k
��׶�GyW�rc7t0��N��P=��[��b�)vQ�Ȇ<Yԫ�+zm�B���7��:�y`��*(m�����NJ+�@ ���h+��g|�h0�[�����`/����K�)$>�{��;�P�oS�YaoZ�,&=DV��*��aA:�Kd^�������3�ǡI@�\M��c�GF�p��{����/�}���g]y�����>�����>��R�hҥ%:YKi���&�����YmF��*�K��%�V�
���jƢ@�UD�z �%�i���&R�����Z�}a ��Կ�c-���6Z�����ܵ��8Ƥ��_�	�^_��B��N<{�UT�wT�9){���@v��g��}�%�z�#�@�:fbu���X�ܓr��A}�U�� �2�p��Ԛ�)9�����Vc9`_���
&�fI�  "l�	�b� �׿��1�8ي3Tο@�,@��f��r�U���Q�ք�%�.	�!lu=�0ޤ($�y��.�nqs�әr���Gd�.S/F�L�Q�%Q�:�G����y�	5EYI��%�J�f��t ��gƟ���� ��,Im����wH��>��j����g`I|{z������\0�"
<�M8�WHX���)dS�+H��j�+�=��Șݘ��߄�H�2������2/f��hN�r��<w"��BR��u0�b�!� �l���S�AD�"R�#���Ƀ舮�	�������O�����Not��.a�5Z�K�/����z?���!���l3��v�[*|�ȽM4�����{���6�&���~o!�t�G�ga܌#K�������T&�� �:�iO{x`�Q�X E�*�*��3FQ��#ٰ�j����+�n�nUe�pe�ؿ���p��S���Q<:�u
�Et��������wBv��Vsu�`,�
��z��Z���������4h9+.�&߫?�ԍ:������a��_�̅pn��c.�2>v7����	ۤ�寨��Z�)��8c�X�f"�&���2̀dљD^��;4v��A'Q{��G�H~L%R��!�Ә^�����gK$�C�Na(=,��0�/�si�M��嗀���|`9�ӥ�K�g��9ם =�x%{
�U��gI2(�eM"��+勺9t����������u�n3c��6Ka��0'N|��C����c:tY��b��ᄽ��DMʅ#_R�:�f���7j��'�,SI�O&�Q��L�-�cۭ�E�%��K	�.��ݧ�,�K�q�Y���6����;����儏�Bo��Hy��+��k�AH��BQ��s2�2����[\��5h�۟�q�`��G�������/����-%� �v��wĄ��������ľ=�c�6LDF����`�e�l�H�$Ӗ{����������Qć4�<1����ߐT��XU$���Z����"�vA���G�B������S� �q&s��ԯ�3cf¬����^�^F��s�#�W��Pv�sw�|���Rg�Ys�q�8˵����6U4�Vi�6��8�H�^�lF&8H9�	�mY�@ s��J��hH`��Z'�W��s���T�`2�e=<��k����]��C�5�⽵� ��aur��S�c�����ovM:6}���4&��pV�^���1SIS������W{���Ѳo�%��K���fS�#	�@�.<��3F4�N�9�;��ʟ;\���}<|`���w1�^��:�]�̈~/5��&�ZqQ��C�k_�5c�2u Vձ�"����F����Cn6�F�YE��1d���&Jg�(0�t��Tqܹ?7�ݪ������N���a'WgD�T|GR��U���!v��^lNXt;��M�I �O�$������ ��2nd·]�+bҨ�̧Y{g���n~W�� �N�b��f_@+v�;����ٓ�m��?}nq72y7�=�;
\�o�/�6���u�C��k6�6�������X���D�S�����%l){�*�O���ِKձD��?wG���#�-uU�_��Z�\��{�K`u)���с���z\L�75!�K�.ʶ����y��s���8U��ž�Čt��%�ˋ�B'����T��1A�/X�~�Ku7�0�xޖF�����ɔy���Ù���LF �i�=]�ǃ�-�ά��+K��ͬaH=�ئ�+�r|H����?�=�*�x�@�*M��\��ś$��Vk�)r܂P.c�o&�OL�͕zɧE�Fcf-��y�����+���m��.��k��Z}�!�$��Tޚ�Ñf�p�*C$)�{��T�SHT��gY����H��4��dg(Wo��_���q��\w�!�mx �ۀ�ώ�{�aH���J��#��^|�� ��/fN�#[��O�M�Vz}OA�n���������w�A4����	��CL(i����rC�:C��).Ej�Jo	^yL��\T����V�D�����+�����P_lO�_���k�uR���Q��D�W�B�<e�1��wfX���`u�>�=oRa�>�\-�F��ΜH�yS%)�U{$X3�$��|��{�V����������Yalu{7(���S�F�$�� �-��d�߷��O�-/��~�v�Z�d7��R�G2�9��cie� �S�p��]���#(qE�$�I�l���1n7/+Z�o���*�%gߺ�C�Qx�h�c�j
�w�MDL7�0�+��A�ک��E~��C��'�g�Q.�WJyJ'3A��!T��ƻIO ��h��2��@[��m0o��,m�;��B��\�36����Sa����Gk�l��m�Z{{1��R�+=Y��� �L���mˠ�@�Aj��{�������C��L6�-�%���Q�'�;{Q��%�4֍�w����2f�~�`�"sAL<�g�r�#B��O�j���*M��@�XD8�]��������1�?9��Ԑ���x�������'�@,����pX7`�m�Z�a�YK��Cu�2Xx����i�8�󔷎0i{<:���Ց!A?�^f՘�]&�o����d�m��~�^�{6	D߁��o�[�H<�A6x	���Ot��ĕ���_(��I@o�!�U3KK�(��'+�d_�;�����51X#oˣ�;���]��nWl�1ƫ�3Nb���"�5�{����~u�l'��lA ^�}&%]]<���}8��ɡ�t$2�cK��l��w$O,�����O����� ;���?L�+����U�T|ү�J�z����/���;�� E~�=�N���M�j&7R��vM���_�A
����Ry�����H�1�:̭�� �dE4D���oP�SEL{����#Xu��0� |�=�+J�R"�V{��7h���:�����-ʧT�-v��Bys��Ot�?lj���j�]Bn�EEx�#�x�~x]v�5����2\���]�0�;*>�E�z۴�+�V����]�羾c嚅�3��t�����
��-(��f���m�9�g���`����i�P��,x:[�'�=5m����6�H.Oh����k�2��Cg}��*���B���k��xd[2b��/�Z}ߋG�-��"�f@��Ěq����*�Q������W7<��2��ڊF�����͂9,�"���_���ԑ�5��̠�_(�\��	}��� sc�Ip<�;��%�">:ts�9qt��"�N�k�F3�]�ɾ����� ��a���(��g˰�� -�e>(��"
Q��I)/�V%�����=	Be�˽*��V�WB�w�����sstW�f���^2�2x��E�H9c�)灕���V�+ޘ�e�v�f�ge��!dl_���p�����.@b��6��`R�Da��~��?8���a��[����|��<�#M�eѰ��%<#󎽐�F=��:~r�9��pt'���(o&�$عO�}�N� ���0���n1:� N���C͉�s��\ϸHR�:��q�ͦ�öH)���,�E��� �_.��Ǣ����<�k�$�ײ�XD�^��y��h��J��|����z.�ݹ��I�\s���FN
�XE��qf����<k̆0���I��xj8�Xj�EJ��T|�e�Ɗ�Q���؎�;n�on=:R���|$:(Ƹ�*�26*��Pوr�O�3�uޥl��������ǘ+�@e��� �+�o�˶���ϺH<�sꪜ��2������W�q���)��@C���Є~��?����z�"�2V7���b��D�� ���Jvg�UƱ�h)5GӎA�6�0i�5�G���ѴW:���8-
��}8�'��k~(��jW��R�X���̴�ܶ(+ԠC�ך^dA*���9��3�l�J�w9�.�R�x��ɩ"�n���V��s�������l�"r):�wdn�0����Շ٩�QPY���[��lL)�����i��2��[�܏�-e0�?"��`��a�:�f(�|Z�#�<�gc�V�H��!�>; c��KWD�HKփ�M���m�x�#-.Z��!@]���N������&���s��g�]�Zf� �w��	��U��}z�pc�X�Ce�v�j�FЛ��v<����(�5�<��M���
�SƇ]��d�\�O�+S.��j���8���&&�}yM(��wÀ���N�M�g�<�V�ܘa��ٍ�?�A� �0��i�H��d>^�N[������jj���Q�'�n_V�;GA�����n	~8���-8�,��w����q)u��q����������C��?�@s����;Ò��BU�u8��x�����_���;V���6Qg�l����������$���~�E�|��t}4	H=?�A����f��}�FKB�s���1H��.>ʔ��PJ��	t�����i9�X(��G�-����7��n���sffk�IQٰ�{���y;�!c����A��,FB�h�޽�F+��<�8L���4�`�˖>^�ŘM��m8��ܖ ���`��ط,�Y�BZZ���ƅߦl2�X�p��)�޶��D���ryX�;�m�/��v^�a�R����-k�)�m�rֲ��N�ۑ�����ш��M���,Z���蹟��L���3�Oϭ���s��Q~�s�		f>�(<	np&����X+�Jȱ��z}Z�����:t5eA*�c!�Wl�iۊ�Ժ|�#�%�Z�+�@��ǌC!�Yd��w�k�5�hL��c���fj���m�5CT��I/#x)o� ����r8�}o٣�h�d�kͰ���?�1��	\�Kc�]B���/�C���x�gڭ�k���X�W�$+���
`(��5�)Ԩ�ւ�Ud>��_�C<��?��"{���?�4_}���y���
��Z��;���k�.�K��9׈ѳXH�P3���pżh
j�3�#5l,n���Ý+J�M֓�!?]9L�����r���sQsCV3�X�PMd�B)LK�����*��ज़n$�sV�0AC��7��)��~�쉑9�E����j��:hE]%9wJ�9C�|�/D��J�
w�#5ATɒizĈ[�VG�%��� �쉷�[\1����_Oo��L��h����p����Kh����ӂ�D���n�Ͽ�ʣr�8��=��3���I؍5�Z�R�+Haԛs ��Z@�a�1\����1��^9�^j/TzW���U���(�D���/�d�y�{�Q�7J�m7�?�F�n��E��#�^�t�Gg^����Mڌ8���`v(c�8��m�'D��> z����4q"!��Kdx�!Ġ���'3�Us��
&�C�L̃F��F=��[9�81)�-�Ni��Ii ��2��f��y�h��M�x�8OJ��o�fJ5�H�Ľ�Ȣ��-�����
��;4S�S���R.A�_	>���M.�KQ��>8��[�H��I"$�u�1��h���5��?(e�2����le�^��2��Oo8Ehj ��?��z���WAWOb*q�~�_����T�����=���3�Y�
�T�"%��#����	�21�yq�u�Z+B�2Íl.��ϵ�!�M�c7+���^�^[���B�bB���q���q�2������E�����YX��d,=_�z�HYt6���bP/G9��}�ڌwΊ��5��g���F��>������:��_�4ǂ��m��6މ����i*Srk�k\���iz`�ބڤ��t���I�������O�j�A��N�D�!V���1�����F�c�f�%73"9��������N��uNs�{�����P�&p<N;PqM^!�L�!��n�2��L�F��~oMAY�����T�O����Q�C��M�y�������F���Ω����q���u�������Xq�����l2�!+���Z��.���궴��� ��R�uɿ,ì�A���r(X׺܊���>���Q���s!��������-�.��h}��Jx"�.�ft���!��S�(�y�$�f{Ӻ���2�Hl@̈+�>?]��_?����j= ��X�]�t�ՠ�*�~��^��5"f�P��ɤ��NT���~.�/��@��d�A�#|1�������B9��rCN�i��cЋ1�)EFO�,�5����i9����I>.�<Uv���ԭ�-Խ脿��m�7���g1�Ϳ�w�O��![���P(�7u�"��'o�X��S��}�u�oR/mn��Y��>1�ܶ��[L\3� g<�^���zuh`��dx:>~�8���6�I�͗�E�'e�>f�u�n�'���c�,3&?
�E�W�D���ꨯa��[�>gy�a�{r�:v�� ��� �X�z�(���9D��IK�o�2��h&����X���Y��^?2�h�zȻ��D�w��s�L�|��k��O�2����f���i!0������}_��0J��Kѻ�]v5~����"�1�vf���~6[\8�Y��B��۸G82(ʺ�@z����$^�_;�$�ǈq�-���0j���L7r�Ux��[lz},O������
�����F�Y�ƌ��W�u�L�6��;�������Ϟ��S���9q��I��$d���jo�	��)����`M7l�_��cd�m�:�C[a�����5S �Zyx@C�Vp��<?b�@���j���7s,��Z����y.5l�ɥY-�֬:�΍P0J�H����X{��^J��*�!�I����W��%w7��QR�*���Yx�J�����8�?�j�N�;i���F��#0���q��`�J���dB�	�˿w#0����5¨���a�Q�!�Y�ذ��ovU���%�0{��/B,�\�$ሑ�6V8���AS��m6��}֖�1���|D��󿦎f6���ٍ�����xE���+�l�I��
���o������	+F8���3�����7f�̻R����Lʮ�dZ��6�`湎b�)�˦�Z��ڝ����+9����Ɂ(�c
<�!͌+����5��@;x�R�T���,�ه��#K)�u6��2��}^݉��4��;������
G��XHV�p2ȭ2-����3���4��n�K��m#�{�w?��+kb�j�%�ZU� V�tQ4���Ɔ�!�ݑ��^����&�1�WK!-$�3�D˔�*�7�L�n��-������6��S�vt�X0!�~���gqƻ��a��W�D�P��
��ᯩb�n"��P�Y�`��Z:Q`��̹؏�d��S�标��r�D�W�;*�o4Y�!���{Q([��E�X�8R���z
�}1�\�{���iCDGk�?�e,�EĊ�Mݺu^��Em��D	�		��׶+�tA��`�O�!&�^�YF̦�î��Tk���Ĩs�e�߈�Y��*�*��^��,���0/G���Q��f�N����si�:�W@XF�j�SK�][�:B*)h��>���ҧ�0:[[>/.��Q��51X�������!�&,C��̳694�㈻�"+Z���$�G��Q^�+^��Y��+�E�9���s���q��>���j�`;"���(bR�m������q�<����ڲ
�7ﯠ�#7.I{ n�ǨG�e@.�#m�
�w���[4�w,�(�|�W>U��9_�><��������2��
QΈ���R�f>�{1���c$�Y�4���
���\��W��o�z��O2����s7̷-�R� ��B��wϹ�������,Y���^�K�)F�}��%v2�ș.��WH��<4}���:�x7�Ȣ�cu1���u����/*�i ���*1�Ş��Yg��H���ijI���^7����Ze"W��²��7��H�[��uRC�߲I�P�2�e=l��W�A����3i��c
�T���T~kV�㫉�/�����:`��q
�zG�a��#���|<I��r}���X�;�ۀA9&h]8V~���b��vo��2"�{9H��K~.�Vi�T�'E:-]3���bi�k���zL�c�󖓔N�yɥk�u&ů�5a�^ںz�φ�N$7����1�V���xՅa%���5�6�A��p�Ar����Nՙ֎!;�7`^�O�n[���E\p��,�~�ޓT������V9k��F��Ī�^MV�6Y�x�k�,���݈ў�|�K-��u\��G��_Y]��~o��Zm�MN��>˅K�Xhae(��C�z[n��^�e�"��.�u�7Sn�o�fu����=MD�
>j����b������~e�Z�kgLF�D_"���e9G���t�������I�0T���s
��Ac�+���f*���� �VJ1����@���#��Șiyqg+yG�5�=�,n�	�lج)G�$���)3�F��W�an��߃�c	�P��ح�`�勠̴W��>;�NK�|�����+#ϷJ�>���H�:vSfb�*����� ��)l��*��N�ȇceH��0�RK&��2���m"��*Z5�:��˫�_�~/^�*&��а�V��9�`�J����Yb�����oi*�0��d5��!s�!v��-�F]KD�sE�-�U	�X�]�	1c�
؜,��*hK��v����2�7$�~��5
|YG��0�ט
�d�]�p����"����ס�mY�ε4ig�t���������(�XJ�`����h��e+.���8wQ�YDu��VuM-u�_U��Xb1u��Z=dXٰ�>���#���<ӷ��l�\���lj�k	D_n=�����vLtN5�mU��YWv��B�,�C("%�-X.�4
�D�H�C���ҥ�����}>,;qa�����fڴ��	:�U�[�p�{��#"�Q�#����Ǿ��j�Y���3N%� ��:W}�x������w����=W���I���<J.z�e;��V||�kp4h�\��,�����񮕈N�k��!��{�ukY*����2�&�`N�M6����=ag�U��r���wh�{�- 'g����농�r�/�Ճ5��.����lv���`�F�b�w=�n	�VS�XbW3�o���	*H0A�n�U4���od�	�횷W���Ph�?�v<�I�#�A�~LB�����;�C��e��t|�x��s���	"٦+:׼�1_ѐ�;�Ƹ�/���*�,���,���^~S��Fm����W<�~��@|j޻;���$ENft)���wޮ��S?	��}D�{(>��QXMĕp�ZG�Ct���$?�,d����W��Y2�v�o�\]�	��?+5°�h�7騦7P�"��̇j�uyOO&�w�1����9�����x$�#�`��H�$6���=*��j�Uq_�ٶ��e��G��R3i��@�	ۤјSi��5��,*�kަ�ŋ����2r٩Th,���~V���y���J�m�q�{J�R*���@�S\����)̠�\��KSGѾ�~���W{��5����͈�D��(Z�ީF�����_@m����sGƕ������BnfX 4
��a�������̳�\�qz�ܤ'�)�$�_8��{��o�'��)5�R�5���������O�.^q�9"J>.<����|F��G�I=J%U'1�X���eO��$ԀLv�
{7���]�&а�E��z�;���_˾g������`�%F�\���3�	��u���T�@���;����[&Ͻ���~�ѥ���(0�m*��W���)6`�.�4��gl5�$�뢶ۂ^�|�)��Y(�j�fN�Rh"��/r������f=��hެ;�C�0K���Gtຘ�ǩI{�y��ͷب�����e`�a�E��4n{O�B3͠Ŭ�f�l��,m�t��i�bP|m����t�j����{�Й@�^����d�(�[4�[��G� %44���,�R���;J`TI_{q���pNd\���y���o���|c��ؒD:�l�>WPDi<�;b��:>����h��[�i��+i�H�g�J��C�E���A���q���چy�F��<�c�-È�ao#��"u?��m6�l�ˤ<ȷ{�'�n�� �	�(:���=���`�/B�^�	��<A�I��?p�e%������Ċ�e	�+�YU ��"d!Ӎ�}�`��s�|��5�|�/p���n���ҞTލd5h	hI @���ݹ�������љߌ���ʼ������;����@�����x�Od���C�q�﹤�K�����{��*�����=��0P�W+�������z��!4nk%=�U�M%�H�9��(�8��U5 tA<d&���C���,6u_ �}����o�"�1^X�T�'�2��.�2��$��'��E{��H�}���;
�Z���(�2����I��#��{1��5��`i���5P�,��)d�Kkb�4�M&~�;׽�q��ʶ�@]h<us�s���QP�"ey� ��������h/�|/���V�<0��ϐ�ca���J�&��Ⱥ��Cu���[�����FX5s�\�fN͓���D Ɯ̐|X�x�P"�hiT�n�Ҽ[͊�9�d���KL����5��9Umj��5��qjW9̡�Dgm�V[���.����$�ueQ�n�Ez�^�H5�����1���J������6�@���PF�43#H3�K~�n�p�7����'�YV=s3��}���p�����4dU��*3���hS��aR4�w�+H���"�F�
ì����uE9m��:�!��L;��Gy�iE`w"�?q�$½K�1H��)���Z�`7G�S	:���G�(���H��#g�ZE��7����1����u�)ɧF������	ϙ��ܠ��'�y�T���qa6H�B.k?+�S�����kE�4����*���s�WCLg���o�%��'a�<�����w*��˖F4�����D[��^��L�P�Is�R� ��P��l�E� �8�pF|�>tn�ȅ�!�;e�*��C�=di�DS���ID{L(-���ٝ�7:�f���*��� �FY����-����������!S��RO���1�j5[C�aaֿ� O&�v�]`F�,�Z���F���V�o rԵ���|�
(���w3:�N�i ������Ej��	z����/��Z����s3
��
a$*9JA?���HRWk��9J�� �a��)��^=�Qkי�+�ˮ�P�]�Tk��癠,�4��2�pv��{�#��~DM�fޫ[�l�'Ļ�l�}�ǀ0K"�B��w��V�2?��\=�>����n���G�}�/�Ę���P�;�ۺ��8�G�C6.�J�q�'��Ҙ�	�W�����PFcR����$fB��Dܪ/H��c��:q���8�3� ����a>V��ݙ��T�w��o�����M�Y�I�$�aٝ��pI��`(�Y�uЎ$�TQ��~�Y#���ȼ�.��ʟ=ǃ2�����d P�xM
xlG��7��	j/I��8���2>M_��~��E����#�@5�F�x��t�H�$td�����%;z�ų����L��s)�����PF�_��Y�aZ�+�����y7�s>��Ѹ;U��!_��F$%{A�{/AH=d�G�)C�G�N�F�3{K
,uN|�ϵES��|`s��t���[�(l��D�u�����\,"���Ā�}B���o^01�J�(�B�d�P���P]��ƾ׆���cZ1���re�܈�pq�o�H����`~��= ��� q����`�_Jh�q���6팏�f,=�2�d�Y"�)5��dg	���>WD������lP,���z�/���޸E�t򌳨��~a��-,�G�!*�N�U��ub��!ԅ�F��mGG�N�����mڣ�Æձ@�I@�V%�H�b�>O{@;��YE];\@'=-^�W���)]��oH�� �l�A�+��<Ǹ�"�{��I���S|�D���a�; ���Nz�;�������a���;��r	�����kԢ�~{���$�Nމ�Єq�a�F���2�I�)S��Ұ��Ȯ�v�ǲ��J�e2}���b��<�:.�/�	W9f�T����)ہ���'����c�A#��퀫X��7�ap�Ȫ���V\h=���iF8z�����w��#ib�n;��D��?�P��23s�3���Tֻ�6�6��8�A��s�� t:���Y(���S<�9���p���*p�i�ؑ?�`���4�x�,�B!��cT&��M�<���x3�K�Z|�AN-:��h��?<$W�����0)�ݒ��x�RH%u�w�'��]uH����ъ�6-����U��4��ɎTpr�g��__�U��j��LUN��z����8U�9�d/}hy���Q .����#p������S���,"��a�s��Y��V~W�|3>։�_�e���ɩ��D��ky(��TB�.8;��HŴX�Wч�j�sG����l�ߊ�~5N����j��h+"��Ǽ�K^�|AEMۭ1� K�M̺��_��X1���������k0(�^�F�����{�,#��)`���W�^���T��z6ײ�n^�$��08����5�u_i���q��+�PIY4�}��!��<��ua)r,�]�J�H\�'�~<FqcS�)?�uGѽ�5�Y#��员�k�d�I#O�"�/��
Hg"$���R<��C�e��
��^�,����TZ�h��	���՗����=sn3��s=���r��Rѻ�'�F?��S�D__�[e�52yr�x:p���٬Փ��Կ���<H*A�CV�z��-�`߀�F^��O*r��qXX���'vl��/FT�O᩹��L��Za���0Ɔ������4$�iglE�f���� �˱�C�iY��^�:`��̶L��O����u)Cjt�D؜�hgD���PϿ)A:,�`xY��<�	�T�|7���\�.8Iy����y9�U�D�OC7����[�_��Xc�|&
�%7r)�Xa�ۿS��&����� ��b�t賛�C	Խ�3�E���;կ��I�fEd��.�6X��Ѻ?�C���9�7�?���?���.�C�wM$+g�ه�)o�9ʔ�M�u����ޥ*������\0=�R(i�%�k~/�Ԍ6x��8�׫it�u�,�\�iZ�WX����i2���G��7e��U0% ��:?ΰ�b:��GZa_��:����+��4�'9O V�:8��PT���T�/ ��,�e^9��^�7��H��E��-PN�/3�k	��4 �ٞo�q)i�Ȳ�^o�< u�����@Q�v��G�1�h0d���69Bq�-Ou�c�5t�����s�F�*\�9h'��Y�p=P��R)�t��w���~-�K�Iz�),��6�����'�-��7Vn<W;�MD�.s@�5�W
��#�9`w %����X#x�tA���7?����D��t�?�l����4I����1+��+��F�_�5 jL6k5��;&!�ɰ�6��/*T�(8�6 M���I�y��V�\�FϷw�L�Q���0�ߪ���BQ��}?��Y^�4IR@��2MB���
66mX��jL�y�
+�_����:\V���玶�"{��#��ǝl�����eӊ��8|v���6�(��n��׸�2���up�����>ys���ڽބ̧���K�`�V^�D����=��'\��vk�)p�1!!�m�'9��^�UNF"�����+p<Q���.4.r�{��N�0� �S:���h�"Y]o�*����b�bQ��[��L�w?�5S90�(�fD(BMQ��QN��3��$_�#)ڑ&�=�<�4�P+vP�]lPB���"˂��41����g#k'_.�y$���>�lIqD�3�T��h�R�;�Z#��`u���|�
�}R���Q��`,���k!k�d���R��N�h�hwa�0��:��E�re��i�!GMb� ��{��W݅�M?�I;P�a�K�m���)[fp��7�V���\�kB�)OsI^�h!�X�:�
<N��K�s�{;	e�H��;���F���pI����UR*(�'62SŃ7CEJ<�z�lz����~�fi���e~������N��_���R�V���t��BG ��s�^˨GCI&�"`E^���X���Ɔ]���7�:�k�
f��2"�z�U��N���6O�����^[n� ���+ߊ^�Y0f����f"�r�5ez�ܴ�����ѻМϚKÖ�6�/j��:�j��
�T��f�pt�L#w�QEs*\0c�2Aw������;/`�����?�0.tD���C��P���mBVkL~�\̖�����G?��.����#�r~mL���6��իfj�2
_�W9��)�(��r�z�t~���������o���)�w��W�se���;�rB8�:��j���������B�m+!ע���$����+=9���)���O{�W�7P�	]0I�����U�'���Q�,&K6����9c�i��b�I�oj����V�^0��/<l�
M�����h®�=?�ѩ0�o�S��+Ln� i��`6F�F��M�IG��X!�:��9�?جZ~�׋����bk���n~X��3����z=w:�b��H��cw6���t�4Sbd6FA@�w���ݜ�x'Qf�cɅk�n�$�=�v��墍y>�[J��9��%Z���;|�mk��� 1v+Q�H.���F7:8�Ƥ�w��c�;:?{	�2�L�G|��|'>���� � �Y������c�P�pȪ��g����T�t�v�2s������s;=c��PC�o�PvI,,}�_�� �T���G�p��!�!,Wa��3W`o2�&�c%=qe�9��1 nT�킇)��� W��� �+m��%��yH������:t�=��>-����M�=�0�x�� W�|&�˚چ0��z�a���`E]�b>=�|��ִU���f*"��Uy�#!��`�ʶ#5�a?D<�qnL���?�a��DK��|�=�#�T�X��T�M���@�L9�M�y�̜!hR���&�_Ⱦ��:ɡ2�3���ɔ��~ŭ���Flv�O,X���{�ǀ��M|�_�릒HY޵y�3�#�%�T�GaV%��y�愇QoR�8�����`����i�s�w·O��F�0D݆�5��C�e/߆��.�Bu��K� ~O<�L�`�&?�5��=;��"п-�ç���+'�_Z�qd]����J$�M,���x�Lu��
z��b��	u��;�;~��$-}݉��_HQ�z�$&�X2��~��h��?��J����k����ɗ����0<��dϱ��H/�$!��P��mdx �>u���ƿ�Mø=��ӝ�0
��I1FQ{w6TP~���a� ��ټ�N�<?np���.��h�ɂ�����x|��u�%�.�+�/K�c��
�!*�}�+84�J^���j�ݛ��T� "F��ى�Xo��0������da���ՕTG�mF���@��/R�_�̆�ۿ���ʈ�D��u &�.s��f�'�Bt_��ͮ~]���l��SSoO�80�|�kL%�T�oڹzT�Hȁ���ǏO�5��gq��.�;-p��?��f@����c!?l�@�,Kt�qdB�H��t��S�z��0mA��sc�m�������zJ�&s�԰��v[K(�ѽx�j�C��噠����7�������YdO�f"��?�:����'��p]4��lŕZ|Q�\3<������x~�`÷����ɴ:8���I�����������%�Vj)v���A~F�SL�ܱv����Enbn�q(��mG{�
������[��wFd?-7=�K����ˤ7҃
���Ά�y7`�K$�!�'���M[�d�n5O	)����N�j/��t�joU��|�w@\'�͛4Y��FsI܅��ǯ'��GO���+��Ʌ&J���T��Xs`��Ch�l�^͐nF��Uh���]��Ǌ	�K�ͱ	��e�_��.�$x*Q=���7,TA�+�� �A��~��aMQ�Mx+��P&�� oS�	b�/��!��9f��Ξe�z�l�JgR�'ӭD��S�%%f~���ԠDv
���]㊸sE>1�u�a��R=�>tM�`�ō Z�k�_����9<��#<����`UqI:x��}�.^=�����DЂܾ�n5~�Ժ��\��� ����k%� �`�wZ�)&�z��m�L�v��ik+�-m��^��l��]�3`��%2�QRa�Hsۍ��-+���K���I��U!��.�_�Ͼ�Y�?<<B-�Ku�c�_i%7�7�8�N�r�����"�k�H~�xѵ�(p0/Y����sۃ�z6�2K�V��˩��o:[I82u�؃�Y�:����⵼�ɰ��r&��_�G/5��nN�ڨ�eH���yQ��.�����~9!}p��{�B9����,�'�/7�$rM��C��k�sC���q�����=��6���C,!�0�l�I3p>/��q�܅1����W�����D.����2��:��`�0�no�u�������p2�w���)���\��0=�";H1Hě���������_SY��G�S�QDe��m��mH�.�T���
kU���
"ĤMj]g���a]�0.�L�$���s�Jρ.��8�����U5��Zۋ�Y���'.wx�<�юu��f6cLv�y����0��olB�����+󧿈j�{��w�KϓcD�$�N࿻/�т��y��K����{"�U�DQ��E\+Ln�A���dқΌ�Dϻ'L��4�<���ts�4����5�#*][���Ey���(jm�r����x�z
B`�x
��@��i��9(q��bB�iϓM��u�L�P�Y*�<T�W���?�i���� ��G�ъJ�'O��#|(2%"��U!8��Л��d宜eY*�x#P�Q\�ۓ�x֒J�	�$=CtZNX�i����+�_�q"=��8hCݹ�I��'�ף�H���8�EN�{�]%�:t^��0i��t!�B�~̒�#��P�ꍅDcd!�>F�/�l�ck�_�ɐhI(�U6�|�M�E�xk���p�����yf���,�b��
����lh�\�;�q��x���yRE9�Ο��'�1�8��E؊ޞ-���ƀl�*�+/� �������W }�z��&�,��Hk߬l��:�A���i�*Q��v^�|��#I��.Ӛ���6���g�����D�6����A\�E��f>� Ba2w(�zp�V��jG�G<��7p�K�����v���h$D�$��|\f���L��1瀄X'� ���5R���STI�
N�8����h�,�Z��{FPw�"�ތ��6rp{Y��v�#�5�I����,�w}�{��8ޝ ����ؤ? �kNRó� ���g)�;XC ���`�/�(𝆦1	R��&.J`Db���z��[�vT��*e�+ E4�[ϘH6 �$��
4JU�d!��`�}���	/hL؋�SZ�b�#�" :��xG���a���'ޑ˭����4�a�:.��[�Э���e~��z[E����>���ÒA9�3�a���P�y-�r��db�L�h�Q�}#۸l�kw����"8U�^�Ew��k�pV��,:rŰA4q˼�*,�����ߣĽ�������	C#0	F�t[����RN�����Ns���5��h�m��yMUh]�v;�,�1S^=�I&�Ͻ�`�A�/Δ�S|����qQ;N┇Jw�<x�}R��sHY��mp�v���Uθ&��o�vX�Η��)�a�F�� ?�|�7�Ŵ�Z�Շ�Q�?�[�����Ō��]���j�V�G����d���a��~�+)(��a��}7j3�<k�]x	�N\�j�@�Guަ�t� ��z�L�f��~��ȈSa�v`�*�ޘoXuX	Ue5�������q��{���'�vP��'�;v\	1�Y�ق�J���ԡ"�[�6��=�)�\cRq��4w�p��!����"X���|���@�|������� 2W�o������U��헐�k��*~qF&����n|'%��H��=N�� IL��&:g#�~�S�>�K�� s�K��2մ����(ӵ�X^�~iyYh�`�A����'�ee%:Oh��5��,� sס1����ʇ�d�y�Z�! 5����B�C�H��*�"�^�k�0mpl��DKniY��ڐ�U�H/�,-nr}�z�y.Vh>&`�o��v\�w�[A"9|~��T���%��s�ml����J��0��{[�ũ���-�Yz��Jۇ��N-��F���e�����t��y.#���~S�W'�e�5~@��4iD9��Ѷ�V=�[WbUC����͋�߯34�Z��om6�����D�%��́��u�pU �B�L/��u\� �6�ŷ�O�O� �S��}�ϸpF~$ۮ	�s�r>$��I%��&�-�*��5�˫�'Z�e�67�N욢P./?��;��F�t���~����Ն��ꀝΘ�r���J��Z'2��N"keK2�6�?07�?W�Bi�/�n!kp�N]+��[ub���	���W���2�hA��<��9.P�d�/�^�^��|2�R�1�Et2�	[����ߡѺO;x��k���~�Φs���g��i2���bl]R.�ξ>[�g"��G�X8\"W�M��Rm����Ӆ�nr��t�cII����ç�P�J��xH#海��E�a�S".^��xut�0�?�\M/�ş�u��<�Q�]���<�8��8�:�V��v���_�^s��ƻ��9n��k�y�P;�`I�(:��98��5���:E��x��
��E�!�<B��0�=�#���c�e� ��,<�Ս���~Cu�	R'��uL������5���4I�ϊ(I����.�0b�����Kj}���xu�����M棩�&ߘe(
�p@i�$�VT�ǡBعZ�av��}��5���x���1�qH��7�..[��橊�N��=��񀽞}�c>��O/P���'��'��ɛ�@�3�	9У8R�=ݓ�*�$:��-K7�\���(Un��<��pR"����˨�^�i��벋([ꂁ�������J]��k?�?�ݾw"<NV�Sz�9�*5��� WX�2]�΋dIņ}n՜܋�݁�\1�K����������8�b�v�;qj9X�a׍�Jv�U2%���t��1�h���[�-λ-���T!�Y���h,��Rp�³|�+�Ω����W�	@�2� �ͬ�" �՞:-�q�e�0v^M ����
��L���{���VBZ���`�F\�8�،5�N�*(�����7d�y���h���B�i|���I��2�y��?%y�x���:FrB>j}Ame4 |��>�[I�I���.	�8oC�7�V\�������[�(�?���2������σ2��@�2����Zł�;�������i`�w���dE��,=7S�W���J.���)Q����Wl����N�߭�"��p�}o�Gw�{}�5��x�M�<� �q2D��l*Z���t�$��*��2{�%���pZ�����kؽ�BV�}%�n��~RB�
Dd9 �!���,��IS�C~i�3.�4�!�����$�,��c���SͦV���s춰���caF���	Q!*�t�91i��޺�;j�Aٜ��M��W7�;pLOP����҄�$U���N,ٴU�x��3lj+l��[SX]�q�������\��8�i�d> x��W�r��:��8�f�O$+������&�*V�,�DP��w�ѤL"&��	����?/�ł�-����,�u܋�LW��v@=�(g[y�f5��N��
�G�������#,���Pf���Ա��1��	;E��L��*-ק�[-�"�X�(�V(��քsIC.3�8���C�9@j���5&����+�x���ϦM��1�vd�yk����#��k����c�3:����I�,�c�#�}�Z�j�q3�.��W܀&uN�t8 |�/�bXy �r�>;Z ��Y�gfm/��5A�#�R0�:ԓ�&�0�C�|�Ň�8꼳r�-�������%[Nzy� �d�|Oք.c�)�l?��i9�@ڣ!�0H�+ ޛEB,ވ$���Dޘ�2TH�L��'���ڀX�З��[�2M{d2W�\�4x�(�="���\�'�{*�Eջ��.��5h���gd���f7��?{J��Z-?��a�?��.M���� ���yϝ�\�u-�1QE����u��]ϟ��Vj(k�{��X�yHy	��*�o���BE���e��c�o��X����h���+&���K:T�<5��V�ɇS����Lw
)I�}S5��;G����G@&�ƈ��9}th��%{U��O#�n1�A�/.�ft�):ш�����O&Ip�ٞ;0���鳺�����*5z�������6�mnې�l�C��
}R�Y?|J�8��VP�*$�����3?*$C�zH&�_o<��;>E�`���K����"q߷T�B�cZ�#�d_q�Ǖ�%��T;S��^)Y+��Ԋ�V�Z�k#����p����|4���9�EXW����}�	8���L�d��M\�pt�hT�7���U�ZA,���e��n�^�aѓ>��ht��
(�CAxM�� �eM��Z �>�ߠ��b����j×���B�^^�!�ݣ��!�p��^f���W� J�{�_�Č�`�_\���J�ן�\���9 �挲��Ka�&A�V�&/Ũ�*�&��Gd3���=`!+�s�J#�}@�UI��V�3��u6f:��Mjzs.Q�wĪ����oB�Ű�����&v�z�S���0ן8�Q����ÛA�ytգ5������w⬖"�s���Ɇ��q��P�䚝x��%�R�Ou�Xϱ%�zO��^�
R{��U�럜n�}��Q�L+�y�M����Ӕ΍D��:q��G����^}���2���#p�_e����l��Ι.V�����}0C��Z��6�HIv(a���%M�e|̟��h���x�!�߼�z����]���������%,}j���8�!�^O�Q;3�
�R���e��W[�����d0]k�J�����G����Y�*��
�:6�O��pQ��^�E��m�F�:�Lu���~���`��r��B�02q,�>?̿*WBYCK�*�1[k+>+�h&p
��\�R�U��S�UB�0�Ft�{o�Y���;���w�
�"L���H�̼�O�&>����]?�ep�Ҝz�]�W���9� N�Fg����~ �^ H���&���Iz��j#��s1{37n���-�d�G�_��a)����CHت���S@>��H8q8y�l}�-2"Ѩp7i���eP�D����	�����_�9ۏ6WM}�|($`��a�l������/Y8kfc�w?$�`H�l��|$�J	c����ǻ�+��1>회��(�U3�'�&����%5��_�+���E�������nƙ/��R�O��$��E�p}�\���i�eٗif�`5���1���p���9Ӑf����%8�'<�፰o)I}
�&v�cF�P��_D�S_�AʿZ�d'�k@�	�D��X�����[�[M���Kb���c��A�9�P���,�._Z��}��&S���p���4���-qS=)/D;!C*Hz�0�j�vDN�}/���Ō�-����x�p�1,Ih�������:6X�9zq��o���b
Sg ���(���}8�+\�S��� i��͌�	�C���&Q���@0�3w>�=�pye��c���)X]�D��aH���pϜ~m�i\��E��B��#�>��9���= ��u�a�w�E�!u�G,�I��dzt~Y�v��`Vdh(�,^��-�1e�t��WM�L�95 "�0Y��-lժ��`>��''*�(�J*��i�g�)�Z'��2ԏo�j/�h��$�/�<�LЈ�&����v�������C�JΕ�o�D2�:=�'H�&�-O}1�Y@��m[\�I:���-�=�g�]!�#�c��?X$��G.�����6��Nm�
�^;0���&�Ҿ��͙�9�Qt ��o3�]\k6���9��_^4V�������-��|h� �#�ϟ#} ���*���،t�M\q�i������%U*N�QHL��Tx�5���V�����Ny��G���O�ч�2�}ha��X<J���%W��'��?��T�s�>�k�[^-"�5$Wn�Q;���L~9���Ua֪�'_3&���.��L3�ѰM�p�"��צ����R_4�Ro�IHx��
�o�@�M�;'��]��3!3z�)�}a�|����8p�e]�o8\�AqեP.�{���-�F��:�E�La>��1�����E������գߐ��:j P�B��M�
4xdw�/s�lO�m~���ԁ`b^$>�1Su��&n�2Z��%�s-$�2�_-i��	��r&rk���+U Z�+e�&�5��&T�_ty�s�߹۫��m�����ڸ�`�t葚9G�bĸOL���cQ�k���WܿXt[� 卢V��AźHą��\��?�|s#�� ~���ݥ�/PS� �G��/���hc�=���4hv9&ƹ�)!��7ca�	���׻�9Ƈ�W#ln9�s��� �7[^z���$0��
��r7l�C�LE�Z�a �k}W-���쪺e�e�I<�����EG�@1��{3N-&lҕWʉ�(C�X�(�W�KkC�bB0ﺑg+��y�M��d%EX���Nv��NS��h�A��9�tۂ����2N&���+}h�Ʀ����%�'�Y�Υk��C_\>V�2������I\w4��d�o��l.`��ڱ%o���
Oi �ȷ��+|ei��$��r�/��&�H���_�dY3[�(���x�=��7��Es�-�W��m$�Ly2�<&:���bɍL]k+~��5~��ea�4"3V�Ώw���򱖅�3���߰�"j��B<u��v0�����G�[7�O]�&���Si�[-
p�st^�s��X4��r�kݸV���"�AQ��R�S1,�(s�_�DN�c�z͢ך��5��e\7��@�!������ �h���L��"�d�j���8D�b���)�˖�'0�y�W^��V5R���j�cQ �:'��H��S��ӱRLܮ�2ȤG�Vl�T�iǓ|�f�\Ѣ���X�Z�؇�rs�h�$Y��2��4��\��x�?A��nI>�/���Δ4`�0��67ӥ��G($�~-)Q�}D�4��͔�Jٟ݌zƶ�G��h�V� �;lfdBI,|y�a���T!�y�
�����O|�IJ���!��QN��l&6y[�D�_�-���\�A�ދ��1�d���6�$�����"i��[#�}#���'҃G��8U�@3ɂ	&'`��pLQC���悆eI�if��߾�R��Yע���k����}�L������/3��V<qW��u}@X	���Ŷ�=�?����	l�%��b0D-1_w�a~�2(��q��%w�J����V�1.�n(�I�
�OXh�G�2r�(�I��	���LK7��\Z/�J��葌K�!������f�K]SB�n��W���]���\��"���)h�`�s�+Qo7���e7��|��0�Ϛ�R݀����<�͢-׮U��A�ӿ��1S�8�o�G����WR�
1��D�ډ��x1 �3��	Q��mqT����m�V�?1��-Q�7�]��g�<�m�����h{�:���^��E�=`}��1L���·D�Έ�x��_ˏ_=Z�E���%���M/����~�r���6G*A���ϳ���MR��V��&��\� Ю���']"��/hgoQҶ�$�U,�ə�\o����ϕ+���>:*}��Iw�nW��v8�ȗ�!����7�V�1�����ԓ�r��rb�ÙȬ2�tba������g�Z ����t�� ��[�G�E�7��:��;��j��-Gn�%i�j	S?-�ì���N�b�hor�4�����KN%��;����Y\����B��:	�f��=�,�]1��@�z�}�]p���0ڏm~0Qړ�� ��J>�cT�K���~���\py�uw7裇���;���m�	;����R��lA��Q�V���\	��2�*[uʦn	5{�᤼)qo}h;����SxWiz4�[JI�#+F���O�{����=�����1������6��[Ѣ6�(t�E�p��t����cd�j��'��YrN�����!��^�8%�|r�H��6ǖY����릷����H��~&��0��J�'_Wl�Z[�묐aŬ)0#R�M��˦1��U�G��Yy�䯕[m��2\����0䓦?������rz9�&�E�/m�H`@/��&�5̓�m4�䛩����E�׌���z��!�<	�dl�l�~ӛ���44U.�)ˬ9H߰LTv z	$P��hl�oS�J��R}�2���\��W��t�a��� �]\Q��~M78�M��%p���m��ypԤaW���k����?>�hv��TND�c��<��}0���#)�(G�5���L�'�o�J�R��=�]1�4��5̽����
(Uf}sqB*
�Ȁ��iXȹ�b��;��M���(��.��T�ձ�w=L_(�y��p���V��ų������$��X?��j�p�VWN=l}������y�����]P�p����To�|�f�ڬ�J��t��r�ܽܡD_�h�t<��i�nt�I]y��Z�9Y��QTg�����)��8�"�`�>�AY�5�G���(2�쀙P��R�z�Yw�"G.��_5�)�\�.A�<��R�F޿gS-��k_6�K�7��A;��!�@-s��-�1���5�>�FgY�	� �7:0eƧ��m��^��Ru���Y�W� >�<7�Yi�۩�wW�̔�����,�T�Xf�`�(،�u2��Le�h+�]"� ���Ԏ�z93�}jO�09^`*����@�sT�HK�Ĳ���v�^��]
ՠ~�`�N <�T������MD��[�˫5�8E;���b2e�(��8?���-����� �B��O�q�,��:�%����D&�ze�m�l@gN+��r@H3�K͖xS�l��D[��_	EI��Mr�Mv��WZ3�G��]�f�Vk���N 1���v���:�N/F9���5��˺0�0�]X@���~�����]TK�6�/�M��L?!�\+�\�fA�"	��+�_B�~�T��ewOk�e��(��*ם�W��&�H���q�*��o��U�`�|l|ݖAA�56IT%�����c;�ŭ#?�zW�:�T.K��L�U��b���D<�T�"q�E����>`ևrnT����7�S�O"kN��m4�[`����=��Y�X�>\st�mjx�M0U�wL������uI!Ȝ��cH��+k�x�Qj�YK�dA��./{>r�akh\h�	�>O<�eӇ#X��h��W0~�N�x��K�QTg<=�>��r������Z�ض��@)�%U����ƨ
<��M^�GB��:���C�6'Q$���:%	��0���;�p ��v�F�#��cg�m������2"����ݗ_���B#̞XM��]iO\�H]�h���^�P��s'M�ex����@_}�ӣ�q�HB�����-�*�$��!���]3�*5�D�0�U�Nh�h$�7Mjϑ{�n��R��GU�J�������7��a��K�1Uu�Nk�SB���kŊ�J/�>��~��@�<q���R��(;����m�*�Z l��I��vf���Mf�c���9T�V����h��E�A���x?����%:D�oL<ۋΌ�t9?���?�KmH�$qt���ɟ�ŕ�.��*����;���yϊ�r]��[ӽ+�� ��	���i��悔�kL��'���y`C�@6��9��ApC��}O�{�M-���� ��Tj��P߿�r}-����Dԙ��4�rB�P���i���+��pUF��w�&}��TS$�a+>D���Q�����p�ઐ-,׹#�3�[��=<TҦ��y���iIl�~�
0��Q�}̪7!�(%�Wn�)y���� ��1�\���ر��}�B{�8����v8˽�TsM���1S���ko��z�V�҉j��G�k>{p$�����^`��(��_>|~}�?��:a�B��_��Zr�k�V�?y�u=�J�[$<5���s!��W���ډX36� �M�f�PS��TE�O� x�x7�$߿��!H���B>��@�>d����q���w�ԣS����|��B'mP�3u���#O��4þ�R�Э����YI�ca=G�Q�4��]��2(����,��'��;��XLm��B<�N�ǁ�8���.��8��5w���ֹ�����a�N���3�o�c�4l�c���iId���b�U��M&吩�6��\�i�Յ=5D�/��G�݁ɪ=��~v�;��<295R�q\y��
Ϡ������W�<x���?ƴRȹA��@�6�,{?�J�m!|tÏ���(�����\����ڍ��0��aT�����)f��gN����)y�1 ���B��(��t���/x�I��ޱ1��q���L�2�"`��މ�ռ��/D��CE��W,��r �J�|<��4(Ւ�Wt��&=����&��}\�0�8�A�b�r���K$ �	�6(
�`���uw	=r8xIՕԟ���?Y��?s��t�%yz�t��Oц0���i���Nh�0�P㮕&�q�Oƛ�><zk<��Q$�.�c*�V��N�=�dZ/y��n�8x�f|��F�z������T>17���63
*��$�К��,�ۼ�w��c��vN�!J%��v��A|�ۦ>"?!;��	�U�N%�=�"�*�r�Σ>���<w�-]��M���$��fjI� �	&��ٰ�v=���;�9zx"Y�'��5�:�][�s�S���x~���#JB��aq�s�r�+�^b'�ڎ��:E���Ϗ�/��/�-ןdb����{a@N�,%�N�Ҋ�du܇ׅ=���.��
���DP״Y�_�V�K�}SF�^޷.�|��G_#�N�_ʓwRr�j'�oՑ9���䧤~��$��A� <>��5^Ǵ,g��
	Wa��f�oCR�SUa`B����+r%g](6a��O�>��G+�	_&;�.Rvd��郐�=c<��5��f�q�����5��61e�i�f�xW+awAe�y��̥�m���ゾ)�'��o�4`9q��No!0���U�!�1��@�{_rr@O��P�і��.�.����ޅ��l�+q�\�
�kQQa��� ?�5=����FL]��WY�R��޳�j`F�[�{z�_>Ly��d3C���6N*�U��h!�*�<����9��u�9$}�j�>���9��T�~磛>\��a(h�����f���0������}h3��4]�UE��o*p�P��JV�R4���	���~���:�Q�K��2�ib����|r�ԥ�֦5Vb���ï*BB1���nL�C���w�T���tK�`�X��|w�=�h��4��^���T�]�=��!��)9�O
WQ�WC!���y�	[�1��+��U�r�kY�ϼ`ŝ���4��0/�~�K��ݗ�x��T���2�!���z�JԱ]�Q�Cݑ�t�K�a�#�%8�3҈7�
naM��8ZO
�e�+k"�u-�hY��S^�8z�7$	)�	�#7�P��м�yu'�
�:`޷�q�Ad�����f�Վ����Qǰ}��<��:k�����S�����P<T���ʂ�B��4,)@��a��ϚQq��6%gE�6�έ��f�1(�޷L�I@�F5֔�Ͱ��u����<�DD��l�uKEV�?�$ʐ⮕Ӊ`�<���:[�r�a��w3iLӱHTW��(d����
��SFA��j�̥���`QR��@�|P�G�|��c��s뚙e�ZIIUj����S���'$#����IH~I��%�ɭ��[dj�yz=o�f�t9o|�~8����4fY����{��R��%�����Z��~��j�9�zu�G�B�9Y�~�`Q�A<�H��5%[�5�9���'z�� $�y�<��0��X����� ����}2��F�����jf���c�K�3X�t�GO�����R��$:z^S�Y���d_�y���'Mm�ȓ^jཞ�����}��5?W��>n5+ȿ7/y���A����y���S��$��of�ȡHe&8�Lp���j�A���5�2`#��p��g�L�Ӯ8�X o���Kt��}���0���nU�l�W�Jy�����{��l�Q��~z��{���'z8Q�o�/�B.�h��1��sG��(pȡ��5]�Z�۪���5BZ�P}Ç�D�6���]b4��4s�1��Ëaf��� -3=M�ˀҴ�ZDgY$º�hmW��Skxh	G���|�~��9�rqbv5��ٍ�pT��vY�9}(�qs~�чB�b�~\��$���֖���nD<К[����q'EI@�;��ӄ�<H笛,D�5�����?9�0V+�Q��
ϰ7k`��8�o��e�t܏�.ByB�X� ��d8)�;f�b�T��(B�<�H%г�-݊��ޚ�򲣓�=���[�=��(�?������M��8��]���v�J�JJM_��l3���;?�-NxU��tC+q	�'�W��r<{���m�Z�1��U5�������ޛ�P� �Ș����� ~O�Fx����f��鞷	�}�L�M�Q|9�!���D�Q��\��}���u�Pc_���
k?�7¶��єm k��Q%��a0�9@�LtIC]�M^�x�?��i�g��>�G�+0��\��<I�P�# �7u��q�|��~��B�U����L��[O\�)��qD��;F��� �V�@�_	ڠ�`��~��eW�AT��K�&�#oV<K���7:�H�7����q����{P�;8Հ��ܨ�R�~�H:?\��R��m�
�������o]Ǆp4}&O����P�S�h��9B��u�D P��u��K&�@�x(������-K^1��v�8�~�����T!�j9WP�:{��r�Lq�.E��Q�7c�{Y
��Y�b��Y�S��7����1[�wX��Z���&E�<��/<h���Gˬ�Ҵr�^�����W`Ae�	|���i$)���Oăd�?�b�P�L8�th%�ras�c���y|PiW^���M�ȋ,�q��l�u*r�OR��+��q�>EB2h�������x��Y��8� ����R�~f�VG���f'���M�C�"}��^��+�槀j�'�����8w`�nQ��&�b�K�P���oC�a�����Y�dc�T�;�0,NB�Bp���u�2�#	oC���s��� ��:�}�i��f����5�wQ�E��D�vf��ν�Z�tR�>pu7����h�m�XD�A�C�04Y�/�^RKRkw���ҙsȬ����Y�^wq+�%-ύ�󛴒D����0�J�FI�c��-f|�X�R�\�7�iM7�2��͑I�z�=�K�/����п(�ε��|�&����!�ؾ�)IB��\��&1"��U�hS�E�ڿ��m;z�Sn��|���w�/^*8n�T��(�,�MIw�}���.�_�����Ƀ"�}���V�Y��8F1_P�6a�e#t�J~��$u�K��� ���`����P��;f���^�D_�&3V�*o'�k��7����3�U��[�Z�{�~;�m?��%�\���ן.�7���x�D$��:+\F�q���|�����Y��^T�wT[�~|�p&M@͹3���{T;*�H����m�!��S�#��L"U�c�C����PAtw1nuT-ws�(I��!�
j�&f���qJ<��7�TD�3�%%N���E^%�zWZC ���l��{i=��^@��f4��-�9S.h��}�9���4�����kP��3��D�ͥK��R��vw�Ux��F5�왊�k�����C~��P�!S7fj-p�w�7I]�#�;=νD��ܭn���?%zP�g�h�	 �>���˗��k��f�$e
Z��ʄ�è���VO� ��������tpſ"U�B���V��F�U�����������/[IX�D�����\�J���PI~L�We����{�-HCDԤ�n�����v����G%�:�Mu?�mG�.�?�fx(�7M.(��@��[���2!??�x�FiȲ���!-��q����vӘlP(̠�P����fb)#w�|'��/�p�1&��̛�JD���F՛B��4�s('�X��;�Q$a������|e5�7�7M���fL("RM#/��[3���P��>.q�P��*���H�����m��[������;O�בּ)�<Ȍ0�����=�`���x��&XT���o�������0���c��as���R�i�Q�ME�Ej�ɡ$�*�j�PjIdy�	��ɰZ�����=��\w���6�lŧ�P��U�����C/�}��lx俜�r��1{3&���5Y�9�|�|���7MN)MӸx� mB���d4��iR���Aw���ZG���E�~�P?ǃw�w����0��+ �"�j~��3H;jLI�7A�����]Ͷ�ǚV�Ӡ���ͬ)��6]
R�8#%�h�Jr�p�	 ���d
�_�U�%=�]>~9����YS�7�!8gy���;S�4J,S��:��3q/��l�,�HB���0����o���d���F���'��/ɒb����X�	$����@e='d@��$�>a!{�� ��5-��\�!��XC.��S�e�j��&~���VB�/�?>��c�i�e/���oqwR�*Mx�?z? �ք�2y91�z�.�Ѯ��ۂ^|~�)�*Q� ����2�`˓�Rc#{�:\�vd�Z�y�X�	3�8�����c��]I4���۝}�@{��q=�h��e�S�S`nB(��_�����=>@�&:��G2 #��?���z�y�?��V,���'l���\%�����Jř9��+NgJ�=^a�E�(
�P�������ovo"D8�E��g�i1$)��<��DC�U�#]��Q�e�U��ރӪ�}�kNL"E����t
Ս�dW�U��|PQ��헹�S�W�J��_2��`�t%)�9��DCl߽ą�U��[����՚����xP"������Rf�����1��7%p���sJ�2�� ��*ITӄ����H�LV�5�= ��R!�2Aqk�=�X��5J� �~��S��2A��� r�{J}x���|/ѮuX����
�M�Y��G{��v��,A%�������S��\�iLKA�;V��c6�Z0y�Fk��A���\⌺s2;�KvL�-W�!�i"��W��vj��$�3�
�l���K�${��Ib��\�+e	��Ϙ��m�Y�!��*xV�GV&)�D��*�A^�f��֤��3�G�V��"J26-�`bq֖�؏�~a<Y�[��*����U�8����|�Ԭ%E�$��t4h(����\���P_k�PQ�	�=�r��+j��2g	\� e�/s���)�Nǅ��`岜z*���N����^��эǸ.J?��L�x�l�HkP���$���'o�V��d�]s(*��kG�>%V26)�6պ�zo���F�������\����÷O�d@��O7 % g�5]&?rꁽ=���ӓ��[$#�zߓ���_w܅��fcm��6��!�ZMqFK�ő��ZϢ�L�0����{!��4����N+�c9�nH�8���M�g��K�A�?���8�^�guwV;�(�?�ʖ�zXXIWH"SU�8�U*P� �� ���B��&������}�Ὓ ��7y�^iJ_s��cZ�29�k�ܵm��+���?l7E<$�U�-��Iq��.��2t���<�O�0x�u��}��`[Fl��XF��������|S��5�2t�-V��4�vȊӔ�@���,��n��Q�w�C���͘��S*{uo������w�m�j�!=�G�����{�G�	:m3�;�)ww��Ƚ��(-D��[�u�`��s�I}�����:�����C����o�D�"kv�D��)Ӓ��Uf4��r�� 5��t�VA_-��I�To�I#��hm��3�ډ��DZ��"�@���'��m�*z�� ������CI�_/��1;Ra�^��YR�H�*�t�UH�r/
�6�����`�0�LC�d�"M��}m�ғ�B�c!tF-B��#O_�C�W���*>5�����1��rW'@��1�3m�f ���!"�"?4��7D��,�p2#��"�������*?�Et)S���w���]H		���z�Q�GByؠV�rd`�U�+���NU��W�,�Л`�*zI��� �2��>_u�=�.�i�W2�l歖�fT�R��x�{J$Bᴱh�q;^ֲ�[�!"����Y~%��Q�����v��,X\��4�/ڭ?F�5X��^����B,E���Bm�E7`r�܎�l9�a��;N*��S�Ց�΢ 
��|�@>�K �����LHt�E��|�M�Ģ��^�oKm�
�k�g����?E�͡ ��WO�VX3#\�9J�#8���R���9�Rm�,�U������1	P����XH��Mw�#��䵨 �9;�x���>��e]�C��&���%�����b]�ua: sFȚ�V-�בw��'[���I�Y�*7��j6eE�/�}�,k�ϲ�����D���u{s�F����F�W�n�����-� �6�E.��ym��F"]`|�0�v|�ܩ~�}����nC}1�S�%�S]��C��
�i#�*/O��%�#�}����t�����wff0�8���;�V�,{���C^�X蟫�|����ȶcԖ:�����r|^D5����y'�S��t��'n�lA�C�14�Ѻ���`�RG�fBw�n�u=��nK���+�ȭ�!�&�����]��-�zhGVDEK�3�+d�Ȇ;z,�bL_:,��$j�]uI?6�R��c�E�xn�1���wQ�p\�x[a�<�&�L@V����sv��\�x�<�V�:�İ����q�=��l��n�x��#D~52'$�x,��36L�!�DI��V�3����<@���K�͈K����[��ӷ���\*��/X��!%�ڒ�Ӷx9���[��(��vɛ��g�4���.�$]�#�©�qp5���U-�fscN��Z��TMv$<č	]bz����Ύ�g��}Qj�<򐨯���;�z���6˩�p�K�01H^�P�D��rf.�RX�8&W��~
[x��ȖF�8(�.��x����D[�t�W�,t��9e���?%MSU+�w��y|pZ�ҋ�LE*�l�T��� ��|����t�	_(~C�|G��\+�Ф�^�Y�H��e!�M }s%�������a�h�(}V�5"�"�᪑���G �nl� Z(�.����L��z�Ӎ��깤�ؙj��7������0����b�$�U���������By�(L�W���R���[���5��Z�bl�.C��s*�TQ{0(Xܠ�)��&[��9�lf��E���B�>/�S�V�T�v5���rR���k!*��R-.�%��PH2�<�:�����Yz^} �e�z��c*Ա(ܼ<RE1p�>��l�(%��$�dَ���/��O�����+'G:O�V}�mգ7n]#�G�:��Z&�&�o;S����(�Y%٣(�b?�E8a�P��]��q�?�X��������p�(�E�9B�i�መ��FW�B�dh��>,�����M�L���!҉�t@N�,(D�پߍމ�����Ȍ�������c��V���A����#<E�@8AU9�nO���-"]sS|q'/hy�	n�����D��K�m<�*�@J�.�=�q|f#�yw?�6�]8��FVe�@��h�~�l��z��KKT:�>~���w�z
�	-�,��>t��t��L22G��"(�����f�����1���M���>���揈 Aҫ9��Ŋ&���=���G˧h��g5��4r�}5$�<�$�~�_}��Qԍٛ��(�`NfLȜ���K�W���b��~�l�>L�IlY&?KnW��W�zk[��Z��Y��G�wq�I�%�u����L5d{�;�;�$�.Yh"��+�m\��9������Wz��)0=��'y�h��O�Eg��'�+��~|ڒ���P���av{���>�ҖW�T�
�6W����y��HPm�IgRi�x~�\E�����;��A�n��� �տU��V>�{6<����Dfi1mo������q�������0��o�%U��ުf!�a0����$YL�@����eWڶ��#� ������/�E'I�F�C�� ��\��5Z��t^s�j�z�n�)�k:)�j֦6.I�C����,�r���[Q�����0�T�L�X[�筡l��Yg��`���	}���(68���?��L*Si�&��1�z! K�6��8��-�"��kG�D�gbn:��z'�{(*I�p_b5�v�]|��KE�k&�U�鸈�K�9mM��_;)Γ���(�l���P�˙�����*�٬�m�`���"�o+b~5��U
e��*��dT����OE�Zr�?� mM�F���r��/R~�,R��.�DɃrą�]����gǙ�ޝck�F�������?�N�m	�ȝI��{��	��:�r%j5Q�)3b1�>�_��{��s�m�rb�|���@�����4k�UW��z�{}�dUK��u��?��Oq?������jX�6�̽l�&6V��Uޑ{eԜ�w#B	6�|ā�U��re�t�yW�"�YԜ��%��lˌ�jCW�tjN�\j�����"�<��@�@�̃�xD�Zѧ�p6�͆
Tw��]�X��k�l i���H�ʳmN�xyRU׈	@��������6�]��y�=,����-��A��$;�T?�l�L��������j��?[��Ԏv*�D
��A:\�g;et'c�c�uf�V�䄈ONTl1;No��n��*-H��3�����ގ�Xd��0�=��p�6b�V{�	���$�{=x��Z�����6Wg�_Ba��$�����+���'����V��%�X7H"va��%L7;O3m��f�?o�I�=�'��P��v�@�^3�b��m b#��ˊS�wmM��0�v�8D��6� Ү�}}%�J+��m+��%�r�91�V!h�+`hQ�/{�`,�9�R���>��F��fg^1�nbߝ�\f�+.�i.��ݐmʈu�Oj3Ѵ!�U� �¹V;�2G�Ba�7�Nt� /��I`h���LC�gO���q'4iD��\�k���d�3|w�t�VȔj�!�X�*�,C͋��G,K�Wa��>�-��$1Hi�0{�Pr���Z�BB�)G)4�%�����	�J+�K�(�/���Ȫ��������Y�(��₡ʧ��L��Id��������#�:�ѭ��Ss�u�L5�Fq�_�v�8f�P��3s]w7����	��7	^�����k`ga��OW~�c�R��!����h�w�;
^�j-�j�}��W���J{���F_�kL�D�:D��'Q�.$�^v$<+����^c_1��Qc��tF��I���L�МX��8�#�s��F 
���qO����6��5)I!�!Ig�PY�"�o[��'���՗��I��z�[�i �Z�2���n����hT\1N(jg~q��U .����|| ��'Fz�
�Y"j��ȁ�`� ��MN7�y� �N��tW[���6�2��N�3�-�a�Y�9�[`]+HDئ����Y���7mŹz������a���

�6�����^q/��%��䫪���EɌ�H�dD!A�U��a�����V{�☒�Qc�UE�V�a�>2W��� h��m�Rl�M�K|��yx�����T��$��e�q��Y�ն�BT��b�I�e�ժ�9����[�>Ǐ�g�8�~,.�9.�S�5��;1���^Q�L	�ILk;Ѣӽ����' S�E-�0����x�ˑ=v��qB�9�)	���2�׹���t����������.�϶ �&t�C��}�,ǀ^��X��ꁣ;�k��zzY��z�3��޾I� �)S��ñ(�9
�(� Z�74	�7�l������,gf����ӽ%��
��r��ƉŁ냝�~��e:$mYG���"+���e"�����^Q��_�ĸ|!cF���fQ'�4�P(<�ܵ|"0C)L���7k-=����I_�dGH����h��O�n/=��D�H lՆ-z]�%��/ǋ�i��6�^ DG�џ�灍��7���p����5v��!Q��g1�|<Q������:K�w��J@��N���wz�v��a� (��:c�̀�
a��>_���"P>3�e���g�q�*�փX�M��U�Be��7��!�'u.gcXj�.6�!"ik��錛gP�>�U��C9V=W30H�U]�C{$QfF�"���=Z���J�eyP����D\�H�P���5?ģ����d�FA4����6<y=>�N�~Z�V�3�m:~���v��>�}?I��xuS�yO�'����6�*�D
����]��%�x#�;6Y���Y�q{��V=��03��8�&�������|�wEW�(�0.�m/K�ĳR�@�܊���[d���g�� ���hf��L�ީ���R��h����:y��CJ�o��x���hc�@��3@J�{��������H8�ߍiq-[���P��o���K�.�z0L<��c��Z[hS8�LT)�`'8���ɝ:\z�p���]6~Pq�b����7:D*��h%H�kn�7�|?@!Ĭ��������22��z����º��	�����[����@x��
���n8�o�.���i���ߟUZ��!�`)$ă�C�CP&�\�Ȃ<4�&X����|�Z��0 ���6	� L��@5�cM��C)���ͥ�,Q��5��4#N�0��`ř��UΞ߅gW[>\B���;�`�ٹn5�'�8EX�<�ʬ��,$��A�B@{�yc��4"��4ҙ�G;�#�S,B.����pmE��;li�)D���
G�����]��e���vMq1Y���:�Fo
C�_����&��b��>�Eo�]'��ad�~�9y��~�gz���'�`|�yj�9�;s4��^�������Ղ�O^��iɺ�a�0́`\�PT���^���~;CVDX���	�2{׏�Lվ;�M�j-��ծ���S�����F:Ob{�Wv,��l�����&�$�<����%0�Q���s�ʦ�m'K�
+@[�����%�d�rݽ��69�=B��1�����e��En!�M������٪��R�Z�� ݤ��� ����U�uq,-R=���8J�oYۢ��5iC��P�^8���E Y�aŪ�ѯB�ңA|߰t*��=[���;�J���H����~c��x�լHJ-]���߅g3��7�nL��,���!o�}���Irm`ɐ8wi���懾O����:�T��[��Ǵ��'�H�
?�B]L����`��8�JM�>��k$���}�ATI�nȿ�+�;�����.�}}���&�Џ�T��EH�%������%��ҙ-�ZW�_�������]����T�w)��l}F0�^�R	�����'Nm�E��P[3pS1h��];tK�j���o���pA��3U5�e\ L+�}2�|8!h�sc�B���=�K�L̻$��V-ޫ�B��4V�ը.C�y=5�"S�q���ʦ��!�������x��0]���c^�X�v��G�pJ���[1t�%Φ�{P�� qe�&z7�����E5��!G{gN���Ў[B+�V2��a�^���Ĩ�)JI��?���Oe���}����Qw��Y�!f�I]�e3���y���NLq� �^�-퐥onJY:hA�K}���H����$R��A�s����['��X-١֟y6]�!��A�O
7�[�
�˺��hq`]�*J_1��|��/f[����sJ��Xޅyd:d���sx����^���̱�֗���b��N=�z�W�b��K��I�g�Y����^��Ї_�W�j���y�r�pv��\ϴ�vg�x��LkXn����J�R>x,�`H�f� VТ^�XH"�$rfu����G�:w��>����M�.fy�8��L��9\����!�C'��j����S򚅣��S�Ҝ-Y� �8&�
���#_��?t[߸I��G����Q���>�z�vOJ~����w�n�x�-���t%����ca`ͥ��4pW�K]�����>��6nIV&O_>X��[mR�h~��?iJ3$��0x�<\�!,|��)Y�[6ej���ކ֫�X���#��8r��VŢe9����#�X褙A�J�~"L���Da;��B\���[�ˎ��M�M�����)?Nsj���l����j�p�}eU�>�"�)�v�Ř��U���7�E�؂�ur�~�O(���z[F�n�X��p�(�8�샖R�[�U<�tt/m��e����_|W Q`m��P6�`�����e|HsQ�� ^zQ- b�1�8G��j*t}�'gCX~��C��A�٪Bگ�"_�n4n�N�"␋��qbx=U�?�M��ꃜ���]�^J-�:^Z^M���l�v{�����s�b�l��p�u~Z�po
�#0?��DP�A(����NLJ�k�Hɇz6?�G�w��WoC߇3�7Y1�4G{b�(=�}q�
Vv(�N��Ԓ��f��ԧh?�j����G,^(�D�TK����N�ܚ�����e@X#�������rO��$J��
Lr�6�~23�iNa-�NoIh�b5�7�0V�z㙇���yFF�	y�̥�i5�f~�|d�aë�C�>�x�k���K���3>�mܛ�ă���2��@L�]�0C�V�^(�Lq1�uk��:��:�֚�IG��B��쁡��p�4�3<gރ`�����]�_���ߺad���:��z�����S� {�I�+������\�����6�!Q�h)YҴ=2��9F�mɒ�(��焠{��)̮ٵႳ�d��0�k0d����lĈeu���gi�>�j�c��ͮy
}u��VkZ������������I��U����ұyeW8:!�1�ٓ�����D��%��7��(&y
Zc^vqo8��h��x�����_�7����[�yq�A,H������K�䵋�2�3'���'fe`�Z^�
�z
�fArdnFp�n��,�$���$9!l���VP�{�H�򗘕?����x�M�Z�I	;�$�dMw�Y9?�xv���:�eԽ"B�ʶ�^�0ow|�v�$a��3�|_�ZRQ86�V'�r|�����C�bO��X�G����W����fh/��)�!�5
�Qv�7%@J�����/6��{�|K
�6(�e�i�muEj�|ډ�'��U:�JXV����WA�猇/_#Y#IZ
��G��"o�-�<0$��%�F������6���"[���6Է:3aj���ӺMBx{IR�M?͹��m�@X\�%z,�c�9G��X�_щb��k�R�K�̟תs�T4˭��?Z,�ً`�d���
!>����}Ӽ��@�4��?�i_!��B]����mI&��i��r;����7��j�Y-��HmҏB���Q�y�gK���Tk	�4��2e^9C�c$X��ۺ�R��@&�Vo]m���p-f�"+�)1�1��ӌƫȔǎ� \���sS��c_Ω��6S����2�Kʛ|���ya�K�x�T컎���{�	f��I�����$�G�!�.p��>PA�ǻ�W!�yFvmwؘ�t$�j A�gPa�xG��p���rc�y��R�<^@p�-���L'��7^�Y��v� 0�1��- _0�v�_�;���)&+��� ���mT˂E4���s`��,&lKr��(��k�W�"�~�}=�֏���ڒ���c����b0�V%�Ɛ������@d����:sO/g���GQ!1B�?]/}@K��jܘ��Лa�8L�<�+�?��!�iH���1X��W�sU�J �dat�'��#��mq&����INO��, \!q���2*����1���,)�&|����	E�<ߊ���tH��=��{_����\cZ��X�F^���Fj]�YH:�yzVJ d��q�@w���w6����Oowc�P,~+��z��RV�\������u������������ں��-O�;�`�V���ɛL��t�j��c^�YKvy�A���dV=D���)dA��jP46A�҆ͻʤzݥS��!�ӌ�'�X�A4�P�Z31I%��O%��=�q�g��ɺ2f��N���fvZ�S˩)G"f�$�� *��!�������Y@?�#�*Uwi�C���h��a[�b�{J�� ��S��
�đͪ�#���\�E�^���gz;dK��o�|Y�8�LV�{���
ʗ"�lB�]��g��/x
&�x�lϊ���3ȾNl�./���.t�*��SO��F��@n��5v�gO�=�q��;ڈL�{Q�t g��1ݕT�aD
�[3%r ܬ���p<q��\�~&��U�Z��01بz�z���ʛ����B�� �B+�ȉ<774����-	c���}�a4�)�/�j�"W��G���}���%�H7��s�� =�{)�.�a��U���� Es.|JR��!t����{nn�Gƫ�Ve��WiR���]�]���1b���_�:E�ߞ�0'
�e����\m{$�G]�㰌X<�<�k�:{���>X)�ҁ�a��bqj�5�����7|���*��r�^}A��|y]�i�Q�f	J�N�-4
���"��P��+%�!.���I� Ԯp&z
�m��`�>��NR��puڱ7��(��4���c��y�k�(d�s�j�$�\��]�X�?6���+�zw۽�c��0�B)�똆�4�ީg^�\�Hخ��Y!.��ښ@�^//d����"P�����L}�6!��i����~�����n���ߵ���溾e�	�'���rl�#餭�5�	����_7�W���`�u�!�g�����ȡp
�`"��)Ѝ׼ߛ)	�H��I��<��*��~+���F:����������r}��PW?V��=�#�EZ�e�������)p{o��Y��:��]J� H�an��)�W�Ȧ�U^_��� #|H��7I�;3�0�&�3`k���H���O�3�Ae���� �a7����AV�ɇ�!�5��6�x�/�Z�z!�hHdD�ІE��ʍ�K@�@vGޅ�{]��J�Ix䈢 �����DݎP�s��Yïp\˞��-j�c_�`P��Y �8��*��vdf z�b����R��<[�����t�}�z��7dO-iF#�g�מ��5�f��.����.�y�U�_�=�^^�����S�ż����-���!�
{�\ V3�MপEY�����Eξ�.�c���?25�~�0��r��gi��%4�i�莢'�9���!�9!tT]C4������Ld}�}@p�x�e�5fݐ:*��x�Y�S����P�!ʬ��Or]ȓ}k�iG��պk,͜��n&ٍ�'�@h󇳮KV�}�=�Y��|�*mjT�.����JmG~
(�v��7Ć3w������f�{���? �ME�*~a�X��.*h"s췙 ��p��<m����a��3�%����7��j��|�t���@��/tl~h��qZb��pV�������6��,�J�:��m"��SaXթ�h�������� j1 ���Õ�6,X�|��.P�5��}}U�g?V�cM; xN�̐�i�+VcY���j���m��s&2�f��+I����%n,{��
C����S���S�%f)�n��������|�Da���C��Qʬ�:.��pG��v�Xc��0,7:9~R��Ri�����q�%]��)��)� �j��5��A��+!��U�:�>���!>r ��AsE�rʦ�Xz��ބt�[�S�6i:s���Qf�P��z�3�,�b�5X�c�6��BH ��^��T.�X9���B�
@�y�\�y���&BG������vYt0^t�,w��%9�W<S��J��q3�P�R�a��N�G�S~���z��t��R׈w�6�{A�\�1�i_����1 T�*�}���շ�_���4i{˘�C�@`Ɩ��27�������]��׏}d���FcB,�H��s�q.C�֋��}��������u��~��ז@�"]���o(�3��rm������
m� �߷�Q��1�:-M+cF	��C�]K�g�E
h(�S�'�h����G}���;� �ϣ=Wc;��8ؼ����ɕGi���Ik$���{��V8�垆I-n�#��.d�S��vu��Mƅ�g��<��*�dD�������(*ò���$�5%������=��}(�
?%����.��׶���ܷ,��>�Vǳ{m}�����"�di���xDqP�u�\usn,�0��\w�zT�gԒZ���#˟��/��J�(�vTE��ɹ��.+�|��	��D`�p���	�{0��e�'3�Od_))�L��������i����en2�h�nn}��կ��Ȧ�����k�#Clv$?�M�g��n��>0���4[R��fsk���{f��.��$3��K�#ַ�g���$С/GvSs{(�����ɯ*D��Iө��Ia�ޭ=�L~�X�*�n!�ޞd	�WN_����V��J��8���Q���'s���ɶ��*=�T��7�"��7�����O���M?�-y�'�[R	���fP����~#��3הV�i$���t��n�-���v|t�ܛ��|ycR�*����
o�Y銅)44j	s���+K�	�B��9&���CE����|�F�ȻT���.�M�r�N�)o�G�=ZB3ߌ ı���z�_?h��g��pt��&�Kη�\����dm���ۣ�%cG��b��1��T�Zj�|�-l�� �_-� ?5|�7�kٍ���+���K3�hT��A)��not�^]i]�[��u}l�HV�[�Ilx
Ә�y�T��0�ڲ�C.Q^
���A���m�L�@6��c��P�gT���oY�q:K�;�)��(4~�F�0D��i�S�06��{bG���4���6��9������l����Q���̉p��r{�����'١�jz�C�aM��-(<�����v����Q�آ�J���>���~o;)�Q�:����� Gj f�@����i?F�XC�} k\����^l�[�;�a����>��N#E��M��8�����䎄���o�v�Z�*+�aRu��T2�>-?M*���*�軳)���WG�t��!֛�+�˔;0�`��"�w�E���;+�,6�4yw���z��z�u�N���p����H���i�w+Ó�`	�MbBD2��H^?#�w x�h�L*�08Kx8�&!8����ks�3�9X�/�#����H���:�g��X0QԱs�%���K���� �9����M��%J�:����oK�cB��K'	a$T�zƩ��J�S��bl]wI��WG�We�- C@e?ǻ�7v�9�������V�F��˵�����(���_�IgX�X��0\Z8�^Ђ��.�ɹ�.��M{ 9��	�(�\��8p��B{��K޼D�y�����$�!H�qAz����K��/]�[�2+�Oo�ޢL�XB4��	a���*��r�g��.�%ԇc ��A���>	�
��I��72Lh�C��#�h5 ����R�jЊ<	_��1T��[���́�G`���Hn�1�B+ɱ�\���; 7�?�ۋs��LD3������	V����~�>��U���=�&)wr���t���8Y�Ӂ[o�Nhח�����U/t��'oF����,�=�+�m9J�w��纣���5���
4P�l���*�g�|6�]�hr�_�~/�\S|��O����m��H��I٭e�����oP��l��EC֓#�g�f���І�,��� �i�_ڱ�+�t�Ԟ�%7Hm�_N�p�.���EpZe�(.�n�)�l~��
�S�Q�=n��b���wmJ�9��.��`�5�V�˄�J��S*��$�l%��E�; �:�u6 7٘2� �C�)7g+���W��[b��q�[=�u [��š�����7��]��ţ�w1�?4���P����[��h6�1we���z���
���;s�4�Z�7�y��A%W�<�4C�;f��:�o�7�����/����C[���Mۢ��s.�]*,��R*>S4��	Tz��z#�=<E�/�o��T��'��k�]�Y�%�0<�̩���;P�X� ]͏�G�?����s)T���,1�Q�R�ے3BQ:�Gwbd�<���х�x䘧����k������2�/�<W�"�� �7tq��"�Q~=�QZ9�T�XŴ�;��XW�d�U��F:љ+�tX0��5����ҳU4�U���a������Y$!���6����6E�S��k �wۻM�C�y����Ӌ�j�:ft�
J�h!ڷ��PQ_Vɠ�HrUক�_��}���LP|�C�R��H(��	y�v�Q��9�#<�Z��2�\�"��5<�J�\lpT�`<�-���Vτ�\�l|�8ߥ ��V�!s��D�ؖ�T�]Y��/� ���u��F�I^?έǌ)�����*;|J�R�u��UP}�~�v�=!\>���^��Kū״ ��zf]{��큓d�
oZw&�L/�Q�+Y �w�I:C5T&`K��r�8C2��?<o(���U�6;_���=95��c&`+q7����˴}��We2c�9n�o��rW�&���=���qD�J�l�?����~��;q���>#G�1f�̥&Т(���O<�̩0��{#��"���H�/%>N8P�n��u�Q[4�l7\�{�Y������������	���vH���^�9Nb�Ĥ�Q�����E�WJ���m>�~�B_����v��TȺ�L�}'f�T�X��))�<�mO���]j�B&�PD���]|
N�$�B4l�^XRnSs=�D|��M�3~�<�"�ͬ�P��#ᶊ��=Ƈ��9^GmH�Z�� <>�X;.^���܀��ǤN���5}h�5(��	��]���ŏ:}n��]e�Ӿa@xCkNAGF�f�`<�Q̀;�G�'#��?���ET��%�? �����U���@&A��w䡰]E;W�[�M7PM�p���,�� ������_�m��֒���Q	�W�(��_�ʵz~���b��Vy���?��n��-��n��Ҭ�X���m�5DK���Ջ���Q*�#�@��<��s���(�-���m���N@QO~�j%v*�}["\qh���Y� 4��6�4�(�Jp����5�千��Y�s�e S]�n�@=�������B0��ꢸ8��R��^%c���=9�̢�GԼ�Lߧd�Ū?Qg�d�W4W���Q�Zj�Q���6M���D�}g�I�X9�R�%���)b�*�]E߯�1业��=�/w��~k�C��!�)���|��~�[b2
,�_s쒈��ԗ�X.���1WN�:������ �i�8�!%n��P_]_9�6�^3"�y��xQp�D2w�gF�2ϭN�J��(��}��B��П�u@>�����I�2
�m>s`�y�C�8�L��ӊ�,��>�- J��!wE� Ռ��m�y��6r`C��0�u�#�t:�sA)�)��:��V�.8!�Elp���t���[��n8�����(�n�� zT_�A`<�V�y��;��������z���ҁd�~��p$p�'��b��de�z1�v��Q�w:3�t�r�&�6��y�.��i{�3lV�u���"Q�<Ӟ�����=5P*���L��D���oe!0�^jZg����~���5(ٸw��F��[A�I�z�`�Dg.���
n�Ne�r��*����_����b@pLo��Ce��4�y�����$�yK�㼦&ƌWm�5�u1���]bi���O:��:FD~פ
�4��l�~�,�U�0&��f��G�ఊ}�)�*�����R�MJ���d��_������Z{�ok$�ly� $8V%���/��ON�-QH�./kTm��L#eF�����p�~Η�v�����\fhB�*�;x��n�u|�掛`�l
(�4��\:Eճ����[muq|�����,�rH&�B�;�OY���q���u�y��#��w���r��e���7rxp%�(��>��#
M*���Վ��I��8|zx�Q���w�}o
���)�7GE	$�@+T����Z�P;ƾ寭R�c�M��G��F�v�Oy��ץQp?Ot�>�x��-qg�����J����ʗ"]�+/_9�F�ڬܐڅa����9�Y$_�;r"ZݤNqq�6=�2�L�j:��Ms��z}!6g1A3V�l�_���ƾJ�f���QE��V�6���UĊ�Y��/����ۿ��9���? E.�<ſ�Ѥ���@,�O��	
�jKQ�s<��w�Bl���3��䕇_i��xD�Q#n��`l�_�z^1*�QХ��~ms�����Y\T,���'[<j>�I�f	��
L�|D��K@IvWӄN�
��D�
�Hd��of!+��$}(+|m��,�]/����<�F���7!9���b"�T�5r�I�~:"��;������R�	��Cg���*B�S�4v���]1�_46�t��!�W�/�(ΐ�A��-���)Y��,F��P�������K�`�m���=c c�B��ʹ4������DG���A�o�k�_�ސ�]62�[����m(��vz���s�̫wd��Ww5��c\��O�E�.z~Q�cV��d|7����]��|�5�d�SB�E��������F�ui}�g�=�%��c	)�KI�����<[�"��Ӳ�Y��m�����k�K
��D�]�t��ǀ$������SN��c�KR8ֿ�ݿ+mv��:�y��ؚv�?L��iVťD
bG��#�l�������8�LE}΁b@6�μ!Yp�u�cs�P&��M�R��{lku
ҿ̑�+=K�*�����8v��)��F4����1M�*#ޔR�E*������QW�x' ������ұ&8H"d�E˞vҚ>�r�����\�1o7};��IӤۑ�Z�W��ъIJ`Z/������0ڱ�,�[7�B �<#@Gu)g���G?V���7E��M�?0��F�X��~R�煫�9-�	�՞](]'��5�ܕ����j��y�'�J~�Pع������N����5�\8ۅ'�v��	�OQ�^� ��y���a{��.�K$l�}�X^g#�pXu�7
�6�A H��^�-I:����:��P���Dw��� 
J�۪o1��ݩ��%�}�djD���T8ӝ�� ��z�aCU���-ւ͎0��=�Õ�;���P������ɬ̦�z�?�r1�%<�)R9��X���1�?]]|�C���6~��� ����.�>�l�--�����]d~hA0?�`�>D�bڜ��'�ܙ�T
�>jERc#<Q.�G������mj"�~i�{�U4u42�^�T�&�P��b�.Zי��p�)�ǒc$P��f�*[�����Y�Y��)�T,$k��:C��w-�\Cг&w��J��H���	�ce�L�x�b���r�̔� ?�R���~��� r+">�9�� �~69���[����p�ϲ>���+ζj��uE��ki{U�_vJ���3&6�xߊ�-�V�]��wAy��ﷻ��:}�C[E�:$�Mt��1V���L뱯6�u�f�c^��^_2�Eѯ"�]��e��á[�zԂeX�aRh�a��oW�x���i6����4�q?� �	az�Ø��5[�-��^����|���p
W�lD�}�'�� �ء!,�^{u$��ů�$�m. :��
���56���fe�H���}H*��prAi���zy�?��."�b��%����t3�K��\�O�̿3 ?)�)��ģF����!�#�f�����>�/K�r嬞������)R�'�Q	�򷂚�^9I$K?7H�$�У5�NZ1r:=\;�b�)��UeJ���.�u�ss�So��,�O9g��
���-��#�P�%����Ȟ��6�҈	�H�����G��v�-��+�z��F�f�c��w@�\�X�x�g�����Z�G77���a�:�h�Q�i`�隀Hp��Fp�h�D��a���[��b�b^��Dn��X5�lKJ��1�}�GG�:a��������a�������d�PN���u�\��}�@���(?ͲB�k�6�k���!Va��;�7� �b{AL�����1�S�m�	�/9���_��LdTU�	aM?�P����7U�$(����];}���f���t������%�#3|��x3�*|���L���[O}럚9%�7f�E2�,o3*$�n�x�R���>E�'
�w#Ċ���9O�����P�F�-٥LoQ��RS]<�`����uws�I��DS|�C��wʩ�,	�3�lpw"��)/�#T5���(�,Fgc�S�Yl��_Q�Ӂ
�˩�O���^��ƿ�"����`��B^g"�Ff�������'ø��T��|�"�p�؇����!�}W����[1/b݌+� (�A�J��j��%�P+ҡ�iôz�\=U$ˍ��T}�p��h���K����[f{�X�kSIJ"�FѰ}P1�3��?��ؿ��P��s�؋?�I��M�������j�x�������u��V�Q��k�앆�Cܡ��I���-㺯��>��䒎y �ܾk\�O�f��"���R��>Oen�d]�m;X@#��r�/�L5|�̄:AM椞���y�{7��BG���x|R��0+p/����VA"SU��4�+q8���v�D֍|�Ԗ�i���m�Q���в���e���faz�I���J}\
f�J|� KڌS��^d�sen�"��f�O�;6��:�7]1��.;�SԺ�^t�i�,�����kՈu�D��sN���� ���#G��F~2�s;�RT=)�R���F}�>� ���YR��G��1�z�Y��B��N@�W�!�]��1.�K��#��M��N {��� � ��i�J��a5�r$;�n\�}n"q(���G�@�QN[����ޞW)�܇Լ:�.5��Ȣ�����G#}���s�z������6�H�h��+>.�<�%m
���Mh0�-(��Y��̑��Rr��L��4�+*������_P���`u��$7��%����@E�@�;d�9����&���Uq0ud$m�2�D1]?I���@���{���gc��4$��l�%!f��w����1��11g7/�t���+�Ǉ^��+?�2|�h�k5|�2/͋a�ש~���^�|�öU-4���90z�..�=v�4��K3�[I��a��ž�J4�x,U�ݸU��a��N0%��[����+`�����h\����6Y[qBJ�w���Xh t�KЖV���|�n#S�t�s�
��>|�E<Ϣ��9.sxm�kB�r4�y-�J@,ez�CD�c��c�0��x��!�@@-�uӝ"�糸}[.!ª_�	�۵_i����A/;d�J.X��'��͔�(�|`0�k�R-G�� �$���S"!
y����`ȎF�c��6��S(g��8��Qx�1SZ�E�"� �D�h�!3��@&:��v��ַI�#� r��3����(�^�_�M͊a0�GI�����!A�0�O���7�����ﭻ��L'zA�1M���o��o[Y����%��F�l�����]�����"���¤�,�xY{0f�M4�р��F�tN��k�<�����Z�\����@��W�7�M��f�Q*���s^݂��冤
�>�n����cF~��=\��C_��u����tn�זMsrQ���W[F����7� ꑼ���^�i�E�1t�����Jm'R��Q-nJ�U�ə�֩���J�<PT�@Y� 5R�38Pf�rJ��1k���u��%&�E_%�0���p����� ��r�L��F��eh	,A����!�}�,��o���6r`:<4�$�����6ش�U���2L�����H�XZ��e�}�����w��T�+�A289�\��TbIL�5�N8�9=@��I��G�O8�z7��l�"6	{��#{�3���s� +2��3z����7�5�]�����S�?T\��-L���G�h}1�1c�ܗ3'O��钠u���w�^SXQ	�C���+Ϋ95��!����bΤ#�) LIF*�ZB���k��i�l(��ބv�����t�"\>����;�B��i{FX
B���Y\zX��\(WB2��s�lnO����VMR?d�,黠���ֱܳ��%r�!����y_B<�Q�bo"B�=XѸ�q/�(QB��(�g����1j{�����9 �G�rx[{H{�10����rQ�%Fץ�Ͻ>G8fU�g�fT;���D�"����Dϛ��sGu"ـ�(��.r-�$e1��''C��T�Db���;�fb�]�pրq�*jhs�CP�������h�<��q��j5.z(zݎP�9X,u��~N'�%Q�G�/2W�Ɖ�gtk�_+N?��`Zµ��`7p(�{���ހ�|	-��м5η�䏝�R�#O��T�Ia�1�F�E_4���3��rOX�����2H���b�"�4j��Y XZȁ��S븟�e�m�m�����k�Sĺq}���g���uhd�c����^Fg�G@3 ������b����,�=���퀸�ҵ�D_���Ù��N��;?'����T�,��Fă�v�}�۲�OB��=zώ�=L����'�+|۬��E
 �b!B���>����Ʋ�y��?�Xuc�D}ן�,��j�Ut��o�)S����q�Mݒ^o��k#M�s���x�#�����lx�� ��'��"��\��>�м���6�����i�����>��!��y{Z���*��$A'�U�&���Ma2��H޲%VZ$a$*z>z{�5<*Dv;���.څJ����ƥ��=%�L����éI�&��&���@���L�j
��I!�s������=>rؾ]�AU@�U�a+wYJ �3t^�*\��W���2+!�.�9�X�97�`囡��D�;��B��Jm�ɴޮ�-ԩ�A���{����7'��Rn�hL�%�ןQ�;�Ќ\q�E�����y���Z&����Dªo�P��e�I���N7������݁0d��y����sc���؝g�#�Tkw�LR�VY�b�Ӓł���#�r��gE��䳛�4�#1��?��ݾ����=N���E�����c%>a�3�u����!��t!���HY�h�<�J�?�̅'St_��	�3!ku�#�J���ņC�:�w@�lpP�#{��p`�4j�+wr͂�{3+\m��Ǐ M7p��a�ӵ2�Ell}y�]BR�D~����	��a˽��\�p_Y����=��>HК4ϰe�"��gw����4p�F��p�B���Y}�%��Ir�������2$��h���B7q����bkh�H@=&�+�BLt飱jyrv�v��Ǳ�V �
����~L���;���篃�ِq�\���,�8�Y|�5>]�Z�s�_�E��~f�q���;<��O���6�䢷�4��J4��0�����?�(��o]�js�x��d�m�c��#�F0_d�������s��b����P1(����g�,m?�bݟ�I��l$��v�U5��1��؆�����>ނ1v�2EH�>^���٘Q�y��@�5��ؚ~2�T�9��5�>�iK�\sz��(g��l�ûs������iN�?��J�^+�^2�~�:޵�Ʈ9�Z��_P��I�(c����:{`��n�+�3Н��Ì�U�12��e�W(%����C���Aۑ��j�+�|�8L��N��$��Z|�U��O�%�b����"/�Wd��N��qua��̉���V.e��?��K���-��hB��ȣ�:�
���e�	�*~n� ��I5DY���E'��W���bȾ4g��Q/u�Lg�¯���ǌ�����܀b��1��df�*;��Y6������k�(�˘gi�� � d[m9`G�R�f2�2��]Y��N�.,��]	�S��ɼT$4:�"*!���JJ�W]~$>�\8ȓB�o�=Ү��=�$��ȩǓ�J�;���3#6
���0��τڭ�3�#�\��?!=�k�"�K�fE�tm�K�r����T���>Wp&���#�ϯГu*�9Z�8b�#~�3��[�w��T$z��Z�s�3MY�!��I$���f��%��`�µ��;c���I0�Zb(V�DgY=٘�N�x��A�-2<��s_�4th��e��A����-'��(���3~����D,O��]���(���!��dF�o6m�PI{>�$����z��U
l�KY���vۊ��E|�5���d�$vj����g�)�ۡ`0&f#�m���B2��DQ�l �����B�:
��u'��sT� ��U�R|�i9��_
���%�1��'�A8��K����kG:Ȱn�l��>h��i~���t�Ѥ+x��N)�W�I�8f�K_��Q��{�о|(�G�6&�?[�YU_�q��xhqZGar���-V-䤿c���{I|�-�l� ^ԜFc6Q'���ėL�cL��	�t���8�o�J���PB[���>r8@f����[1�Hq)5��Y8=/�-� ����[8j�����3�IW'��
�"��� �,�9
l�)�W�7������qo��A�����Rd�g�O��jW�4�O����跷��6nÐ�S^hsr�Jr�������%���S����*>�C��j �v%�,��6��ݹ_|;pXH��$Z}���:5^��cמ�i �0������b�����;��	�	�{�x���4��q	��K����z��l��d���}����n��Tρꮶ�DLw�d8����M]�'Lt���|q���O���}b��r|��6��ו`hy��ǍGa<Fʯ&$()����q�K���x��P�O�]����"�+�"r��N�>x��:#z&3wX�P�4g��Nc��k���i�f�[��\dH����3XȻ���tEi.lB��W=1�,�<GJ�b�up�KF�K��	�G^C��G�[?��{�C/�0������ìh&E��v�Pk����~+
(�ٻ��.��g�.RQ͎��P'�`3V�<�[qi}:E��/���GOqi1��n�U}�=����~�0RBdM7���3A�z��*�`.i�J�)�s��)��%D�Q}bs�O����Cϛ�w�k�W�1�z�"���Χ��F��dg��w?H��Y��Ց�5yܑ���q�k�p���������: ��<t�4�	MU�|`u�(1��ZZ:j9��2�T ��b�b�}�+�bܩX6�\���	a��{�ǟB�k��|�?u�*��<��b;yW��Y���t5<��������wq�4w�{_��`������] b�U9��r� ����O����ڧ֡�
2��a��&�X	�����"
�d�ڼ��\+Ӄ!z��=zk�_f��}P
VL3.��g�>�X5��>��3>lKRy�+��<��Y��@kJn�Ǟ���`�pHao#���ꀿ�A�`� N�BIǱ���X��Yo�!�
\��:�y�����uqv�$�>P������i�(�|�z��t�.T�?���zJ��5�q��W��;�/��λܧ�:�z�-��l���*�dD��Y秭���v&�Z.���\�����'��]9)0�a���c���vR;����H���"�~
�[��6�6�-8d��FO�{�8���W�|�2^����L6�	$��](2g½�!Z�= =�"Sl����k����p�c"���RPQ[`�f�N
k,�� �ñ/'Ҟ9
t���̕y�6`�wڸ�SM���L�!`���_ Fv�B�!O�����:���Z�����Ea��v�d����"A�6Vh��E�I�K(9|̈�U (?�|��͟yث$8������zj����{DoxE$��d�n֛��SN��o�q��0%�}h�s������ ���:���j�k�ܲ�̾��?L3��]��C&��Z���p�O���k��0��_L��4	m9�OJ��'�=�pyzPb��cj����.�қ_*�yVEX4G�U}��A!Bb��g̶��s^� e9��P؟������f����/��9��)��yq�𳱱�"3,RT�0�Ԏ��*Q���L���AE�	ș$^%y�����Ĳ��wT����V-1tU=o�lvį�1�3��s�b����:�����.�[�U���~d;+,�EL�Ї#������RZ��7�s����ڧ ���R�غ}�,�=���㷵�8�E:c! lK�nQE@�ӄ-���=t����P�$�8\_�x̀?�����j=���'9H�Of�)�]i90ޅ����b�6i�E�|Ex�3�&ٕ��E�AL�/�Q�HlGX���3�*�q�jԎ������f�y^Q"���Z��A����@��O.���T*iG:2@��7�,���ee&M�zMg��ln��n?e����2�@��z�b����|��W�/\ ������Y�ͥ�@��Q�Z���J;gڡy�XX�ұ�R�;@�^	���РO�����4n �
%��P7��û�U�^��)����)cb��vX�΃�q�n߭el��T?�
���qA�_����+�=���B�9[�k1%ƫ��1��n��3�{|�]�ʜ�ؾRw�.[�9�%�ߙ˔�X���Dl#���]����bt��,��D0(�_��YEU�&hWN8Y^���/�T�o4#pDŌ�B��������2"��!$��l���snwg���Dv�����BJ����KE`���%�bӽk�G�O6����`�V}��ЅԿ=3j�� �D*�l�����sMw�&޴AAn4߱�w#�D��#Bp��)��Py/�pɻ��G�W��Ʃ�v|I�DU.�G�Z�a��;Z}�Am��@��@������<[��N�`���r���z;��ӞY�і�J��#��d�zt� �F�*�#��;R"_g>b��~.:V�˙�aA.V w���D�ƛ4o�Y5�Sw�,T������dZn���]�o�j )?A[��q��H�����S�.�&�vM��F���C�)Y�X�a�L�ua���9+�����ԅ\έȉ4�fdn;r���(�>|2Sd�F ȯ�#�*DJ�ǥ��zM,�^�J/Z�kC�torxs�#�G�}�b��3��j��j�v.�/�CS\�싙�6�tf�������:�����3~Z���:t4�j��K� ��*����^�q��ȫaQ�½��atS���ō���Ơ8����b&�i�9�̒�t�yQ-�?�"Nr1��sX��DDt�|c_D�E�-�5i87PQ~j;S@[C(S�1^S��B������A.����N�ncס��<:o[],�PzJY'0�P8"���3R�-�g��L+�v3���R6B�	ON��W�tF��X1�������Vb���^�!������V�c[�ö*�+v'M�6�`�h�L���k���S�sY�;�Ͱe�E�0"WV<}��*� ^�
awr6��Yol��L;�m?k{
���߬��(����b,iqÉ�<dW�q�t.�UW~!�T����K�� e;Cw�)�n������|���/P�z�D��ݱ�@yU�dĹ��ʈ���D!�������b �
����q$1<C��F�g9�[q���z:/�3N{��	#���$uXK1{�yn��J�Ρ��_Y\Ǡ=q���|��P���+�y5-��ӫ3��bt��m�{>�O��Hu����+�1�gRE8�y�e��v �W����s�]r�Wn���F�%�κ0�1#J0R�U����X?��~�󯖨��Y-�v"�D<�9�Y3�h6r+Q)�X����	����ب��W@�1/л�\"[����$�@����;��>�ȗ��B������xD��Q6҈��PKMw�T�(�&����X�Z����.GG�G�|R)�Sq��m�b�')�
�]� G�I�B0p�D-�����*��{�ElS��m�85����8�N�b`�h"�q����5!�W��L���{���b[.br��k�i��G���F��&��A�Z�~�x�$qb�d}ξ���׎�����LO����M�a@��r�*��[���C�� �]	�߼����O�ٵ�^9yu��[@ڿ5��\i�-���K���Y
������g6�����8���\{������h5�Ri��+voS��2fZa����=�B�B	A�E�&�;d�����8�X�/�o�Q�vZ�����ѥT�̼�1���n�>4չL�k�L�O�}��i|`��;���wI#R������UEd�����Sп�ZH+x�KR�EG{7��e��L��7���*n֊�ԝݕ1A�����W.n*��*I'�1�3zG�`[~4��%��S�kWc?���T��@��C��<�kIB�Ew�}Ziz�!��^O��(�;B�j
����.ݝ$"��a�CM�CK��v��N&]ŗFa[����$0���`!�����f�(���ɐ�`!����}y�b��˺�'�7�,��$Z�Y��%.���S���I6Ű�3��VDk�����n�{������W����=^�U���I�rw�~Fp)	u��g}��}8�#��������ݟHg�ӌ��iv ��1��]`v����[�����(�n�d����l��<|e�Z�ME������pj	RvaԊ�/w�4����h�y�4[�Dh@="�����%�4��K�ZAZ%�o^.px�䕃p�V��������6�\�b7�x��\qv3:\��,��t�̼&�NY�J������@;pj��C0x���n%����bSV�K�����ڀ�Ee��E�Dw^B�ff�ϓ�b�Y����Լ�7��Y�q'���񯕿�H�������tM񿋋��pז�8�K񄌇Cq�}R4�txhC���ݖ�J�������U��O���,�0KRW��u'瞛�����*�NL��|�O�8[(H�u� ��dLA�bs�?q�s��/ \ˏ��~s��̽���X\րyU��S������S��y�&��fއk�9yhӃ�v�mP�Y#O����Xv�q�>�I�0�7�:D�}�>]��"�Bb�1�<H�� �Q���)�Y�5�	���e��tF�֭���|es�%-b�lR	���Z,*C#ؤ�����R��c�j�W
����M���x�\��d 3t��n_�:�/�D��Q�2�y�cQ�HE`�Az@�)SmT�(BqY�:���˜�]�q�"J��[.�ρ�)��`H���>��W��-=j��2aD�W��`p��=���mi�����K����|�2r�C*�[Bb&0G��'��꒬D�
e+��'�s��s'Ν>M%�%�&M��!��#@g���5�/dv��p���o䀒��B���;d�5`�Rқ-����U�ƫ�4ʊ��?�@h(_)૬*5In\[�N�5d��~����5��R>���h�ר�lxddF����� �aJ]���U��gne�_`r"x�8d���Rzߑr���1<U;�e�=_�ZQMCY)e �7� �*��Pg�D�q�mf�&��C���h�B���(;/5<��\�=�Xy���N��2S���"�@���cpz	�V���;�5ɑ�8R���ڛZ��v*��S���!�k �V��Mv�&}�{7�
���U,S�Ȃ���>��c�'�_[�v\�F.�-���b~�g�P����
��%t�3`���ei�|�f^��Q���_:�=@��.�`���5�{M8B�>�3�2�0�!����r�Z�9�ˆ�mY������d��s���'��# �ZW5xm��.�c�XL#Hי� @�fcx%^�{�]g�`2uV�x�5���X�0����DdUJt��ɢ�*��S{=D�y�&b{ڢ���`�}�VF/
-n�a,�A�����%CK��0�y,׀����}���
�0�UJ�vFb�����E���	��e�	ސ���G<zpFjv�k�.��scG%������Zxp����N/�u�ie�R�Z,�����s�2H��4�-�w`��\6؏�ZOS�Nlސ�с���R�R���>K�E%2�~t�������ʁm,��Bx�Tg�g{��c\���\����o�m֨6Կ����kQ*��5+_��+;�[X�4H˜1�\� {����T9�>P��� ���z]�+����^�O���dF�7�����(�(�P悺�c��;��W���'�V��~�0��ۈ
N�hI�l���t��=��E�zn�i]u녥�B*O(}B�j���R���#!��[vص�Vp��aa[Q�갭`��R�֊��o�,ފq���T��ؗ�t�b�f$���X�y�T�[�9~���Ft��Uۤ��t0����{wnF�� 1%Q˚�E���~��j?l�]�M����g�!ۗ��6���+�M�v�c���*b�-��3�Z,:�6��;c�tx��'�Z�xiq�-�a����d�S���k����'�T�>i}�j���^Ӂ�]�cړ�O�؝WC��E�h�	�e��u�QC��߇��g��3�d��x��V�e��9[�#�'ߗ�ɽ���/(�]!�7E��@M��v�-js�aB�w��q�c�\�"7p��Y��Lq��}!r�Bz%�6�>[���s�`g��Iq�Z.L��bC�ڱX����v��'2,����$�$�+8a�S� =���'z8"��A����Cg�M���5W�bUk�#Ԥ��Y>��¹`�gV7S� �<�æJt
�y�BO6		H�~{���l�S�w����"{0>����� Ѡ���0�*@0��RT��P�Z=�	74h<�24͸}�%��� �)���"���h/�gY=+�K���=�>r��u^C�á�	ȹ��*�L����g\�9-Ǉ�f�G�^��>���/���mT�����a#�e���',��R]pIh6�h�] �ʏ�`0ӻC�yL6����`���v\kD v�l+�e���u�A�D0��6�C�8��5�2(�{ە(2]�1O�^l��e�ऀ�=�����k�B:���<�r�2�ݔ�Q�R5�#����;�q��ٝC-q��v���ժ�g��i<:lҍk�'�g� 9�Ϝh')��5����T�~c�BP�]�
�LM�	���U*dP!�L�D.��v�ʡ��b�sF�*��]2�e��qk�spHb�A%kV���#s㐗u��XX�(x�=�{�G.+�}�3�H�>଄e-y��d�l�B:�W�VA➌6Z������8��PҐ,a��w�f��1����}��h�{���"fbT��Qq?�~z�fba2ޠ����[�L��1���w���"�l�m�~���W�IX0��Gc�QUU?MB�v.�������3��HCSȮS��C��i*�q�� b�;���a�_ju�>2���w��&&;C����2Pp�rL�!�;�J���?	G�ݥ��	!��-����j��-T�?ԝ��вԌ���E�RW�-v0�� 2�;�?��u��4�4Բ�t$co���0bRJ�/�	W�kW�̛�����bԼ^q�߈���z-�mv�4�#��jE�?��r	o�r�~$�|��[ ���?�>�b�V�	Ñ��
υ��㐍�O�:c��A��8I���D$��h�@�늚��ƶ��o�*��?��s�c��3,f���8�R:�o��
|��#����&L8,PX/�x�� �1,Ԡ�1��2��4�4��黏�>��*�3!٨շm���W�2c�yiL��K�S���۷���ԇ�E�k���S��a�\B��
��
'���B;X��AF�K�����A�YR�S�ꫧ��H�[�{����7@ �
�OF�\# ��Ճ.k�u/d6y�b�۝�mhe49���V�34�k҈��gS������@"X�^�@��þ��?h^Ӭ(����C�/�d�r�x���B ��hrռ`�x%�<�t2\M)���Q
N�x�};C�-���7��o����+�@N�h�&�t(�O����W�H&�틐����d�������P�܀�?�O�"7rX=1\Nq}ӦߕpI����D�h��j����}&0tѪ!�Q�Cm%f�j2S��q*��٩��R�����棆��>#�)��Zx����޼^�`gR}�e�GA�iM
5��{����1�V��/�y���c(��N$���%8�/� _^��G/UQ�(��x�Z#x&}�j���� ��� }�Y�"�y���9?�k�2�	���579�v��fl�f1���DGH�"W�\vN"B��wQ�)����x̅��0�-����]�^̗^��ؕ�;N����c7����~���tb����x.t^�y.�9�|}��R�Y�<�z���Ǒ����V�?�@¨����H�2A����F����!hq�؊�"[gv�X=�U{��g4�a!�wҶw۶����F@�u.�������(�s�Yf�/%ϲ��W8s������f�0��T�nQZb�W~o��;�ϛGmz'\7�({����p���8AbƭΜ���HȐ}bjȚEy�vwE��O�����%%v��0��-���_V����(�4{ٜMU��`�rU6�h�h��9m���������v�&�ԁW	Kz�2���^��Q�t���B�v�UA����X�d�nU���U��I�|���I?2��	l�W�;q(D7�����S��Q�qȘ����C���ck��AO�f�u�������w����-d��<:Y埾!;f��������?���\@F傤��s���a�4�cA��ݚ����')|4/Z�*5�d�Y1W�VO#D����$c��B-�P����"��gj�W���5�W����3��k��DSk��!T�
〢c�dτ
�_F�)��]�͆��+�%�#'TpC��>��)ˢ� ��)'l7�,��-Wq2�Xw~'i|M�h��&O�x�3 	��!tf�����1n���������������P>��,	�b�9QjJ�g�hk�{V�����D��\ɣ�riy�b@��*���h��+�3�EWi<'u�K��ZѦ`/X��2|=�'L� Y�J�6;w��4�Ld���S�Vc}�i�C/�Ϝ��(	_�X����\����I_�쩗�tc�x�$կ�V���h����F%˲��7H8@Y���x���Vy�uy\2'����'�9͊��,S�c��[,�n��-\';����SC�o]�=$sSr[1]�%3D�p݌���É��J�~���F�;��FI�`���y��)����p��yPn��p�t�gQ��܇��Q�;n`������Cl�"���]���27�ly)W'Oayeyۀ]^S2u�x2��'18����`��)3E�,fc�U˷�ǯgO

�g�@ܧr !�v�"1�mJ>�ږ�~��+�����^Ȟ8�D��V���t#gwdg~\�Q����z������ס����V��x��ϧ��3�a�
�c��Ύ��$�*���>_���ғ��;��]�b輺�_Ϟ<B��ނE,��m��4!���+CO��Lӎ���4��t�4��!^D�9@��kUB}��Wڊ���^Hާ��L|}fR���{&�3W���f�*V�$�ytڀI�*�5'��p�
V34�:@�[��KՏ�KFAi��Q!EtӱF��6��+�d��O/Oi�N*ҬꢞdC��sy����$᧤�l��3Q�"|����:�)B�g�L�_��So��%��[��
+�K^�ʇ�����2©�� �f��JMK�hR4��$��0K��dF�	���:ț{���]�x�k`�*3���:�F��u�c��۟��ӈ,��o�Yq-,\��Q!�iCH�V_#+\������찵9\�/��P_��$��]bCEsH�	j}<ڝ��<�a� 2���R�u0DFmߍލ@����TL{��J��?,���"gc����cj���J���Ч3�M3e��=�Z��Y������	��n���\*@ςo��/��n�tɧ��.9�;�QLF:����Z��C���֘Y�&����ﭓ\�w�nrŲW��mSb.�O{hr�c5S#����y|\�'Q"�Y����K|��s���\��9���4TM�~�n��؄{f���U �A-�M���lf��O&PW��?+�זK0�t��In�-4�8�L!�~#H��`���{4�X<ʣu�T"J����,;66�33=�j��};�&a�^z�2^}ρ�P�|�}rX�r���!���Xt�n.=v�pV�~ 1�wP���a N����F�TL$��:m#�D����Z�\�QƏGIw��)����q���T�h�d�@zv�v�A:4�������Gׅ��
�Y��/�+���*�9ůІ��h������G_C@���~ց���v����ZI�����S73Oِ�L伿�����,�qm���3%
�wξ�M��X0u/X}#(E.�@̑��y�v�B�h�Oڈ����57�p�tN��J��pɸ��ǔ��<�k'(����[Y�~�{��Q�M�z���[l�����F��r�K`�}Bv0����5�H<��[�[H疔<5�ޭ�'<?q�"��%'���#�~n�e/�? ����
�bk�� �q��qA�Rc�S�[�+�X`� H�$�l�Bkl(ԕ��S%Dq����]���q�˖d��χz�1Q��X*��]j�I	v������G���ҹqq�_cU��XA�K�U���ǲ������o���7�ߑXP�'&��.xjǱ/��->�l��64�8�rU�iU��*���2n���������³rQ�A���'�6�e/�4K�³!rp�qv�z�]W����献��V6��>�K�,�$�����L�`mo��Rw�.�@����G��L��y�Wr��_6d����b�iU�`zM�#`�O�6���H6�2D����`��2�F�L!�C���@OZ�����{�&�{I/orMѾ1�:ƥ��	Z�]�y�M�c%2�3@��PQ������h ����;��WW�i���9�����窰X;������P�a�~H��ʐ���0��|��@�"�V������"�i���-\�t?ڐR������Ȥ(-�|� �5i����V=�Vw�3svE^���۳Q��î���ID=[�<�h���E��ii���0�DHB�0'#@쿅	eŽm\��f�uV��l}�o��O*�uN2�I#�$c���8k*����k�m���͓�� 30���p��fHYΕ�Na�)d��Ϛt�d�h5���B��L���S���(|'�U�����>��vs�N�l'�Ǟ���L>��ax�Ȩ��VF���Ѽ�����"D��h�2N� �:��V����F>�(�}�S�i�5天^��˩��4��"��iG�9�įNe^j<�Q��+���k9���Ʒ�*���j�L$��V�Zs8�R�K�lg,��rI0��%l"r&-x&ߎ�=QH����@��sT{s�����R��yYY���D�Kԑ���o�k�}�����+v�TYǉ|j�5��x(�*Z'R�%���\ݩ��C�:q��Be�^�y����R�:׻��Z�f��c��7�%щ�Kfp#Aӓv#
�H��"5�����o���@5�܇h����?��M�|9c�ʀ���39��w�N,
��<���sL��Y�4�@.��F�g�Τ�t]?L��eO���8� ��l��<�{����q����5�U*-�^����"?(y$y����o�y��Y�S����X
n�ν�� ��;�@wt�r�b;'�1��p�ю�/�Goh ���~^�X�h������jƥ�B-�m��KD�V}5P��Os�B�[����a��������,-Gřu},�\�}������z�S���&���㿋:to��{��z�)��9-(GD�>d��,C[ţn�<eJ
�\�UO�#�g_U���F�����l>���0����&�E@�8U��`g^R`�`�ƭ@Ekd�Ҽ�+��y
�^��F�Xt�OxG|܆�����Di 0�%�9y�-�b�>z� �E���� #7��[��45~ej��_{�ވ��@�Rz����ʍnA����'W�a`2�_�R��{�h��K�w^����Rn#zr*=�o/p�,{�"x�l��iָ(���� ��cCQ4D��� �_�i6�i7Uʈk�'�W�0�"@�1V�H��]��(�:����	@�t�O�:������|/��O�~e��ҝ Q��W5�����y@z�x���̆�%�|ԓ��q�{�MpN��w��:,%>?�<��/)wn3��F��ֆ�..�*�§ʻ=c��G+�렯��7	��QKn��y�dWőm�U�(��Q�<K�^��<[j�~mj�����9l&(��/O.�>����D.aD;RGܝ����w3$�:tF���E��c����0���A{�I�{�R��Ģ��!Ҷ��gȱ���%��#�.��DD���p�<���I5_{8:].�A�BX�zM��ѹܠݭ�VKE7\���o���R���l�Y��H�>1g� }�4�[7���8oY�ٛ��� ��9Q�Q��zcfX������>O�ڇ/TOc?��wn6.K��3�k=_W&.AR8p&��mAEUw	�F�o<�R ��j��3Z�ꐨ��t��ދ �K�����f�Ն�v#K4���k�>V�ߤ*G�ئ{o۵=�'[&#v?�R��+[�'�oF������k�̽ɻM>���rؤ�NUj%,DfÖ{s�AS�22�d�"����Lw��Bp9����"���^�4�F~�.2Lzn���Y���H�g;��n�2��M����l��0"Gd��uU5�\sܛ=j������XG��A�t�f!?r!n��)ct����9�z�
�/9��ۡ�"ѭ�H���b���NL0�(��}9����*��¹�d����yخ��R8-�̅5�30��z�{	��kSN�p�	dǱ�Fٚ�AG�:�mb����18�o ��v�8��ď��9��6w-y��W���:�E�9D.c����V�"ZS��j�9H%� ��|�9����Cdő��N��19r����UOq�X�I�^�׿�i	�)�44�8���t�]������d�%ͅ-��m���,�`�ƙ>4v.	8�!�˯
�!�҃T ��8eJ!�'J��\R��Y�������{r�-2��= #G�mM�2y���*Ǚ\/����%�aJ�~�7����,~�B�6ܭ�󴺕����͖ঀ~Im�P��e��3��7>�Z-3��v9��\���M|)k��Ǉ`�a���8�lk_C�=��ʺ"��ʹ�#�q�����r}�@�h@�7U�
'=���#��A�ޥ�]	��Y�r�J��B����V�/)�d��=W �=7�����U��`͉�'xeO\(��-i*KX�~H�� �f�� �!F��2�cO:r�X9uZ޼@��ev�(�w�g���-�
���ɜ����W��t�|O��)J�RQ�Kj��^��vAI���i*3��� �����-��»ퟳ��ّ���x>{OC�7Ofc��ǥS�2������r�"7<��V|d� ��!Er��Ɩzl:�
�2H�Չ#��ܷY��kv���hJ����窩�8u.w�kf��T6�u� g��`����^����OK��dޭ��(#H̝�yJ9<����+�6�:{S��0��*�����䪎qP@IZD> n���� 2��L��e��ݘ�I�Ϗ���Ϫ��w�{��ЖpZ��'�V�qv	N�~ �\��l6�-���iX�b�k���Y��pϙ��)�r?橭"�𵗺�7�P2�J���y�
�9$�HM��IǴtK/z�-J�ҟx[�H�E�K�ChH�IR���@A^�L�Cy�#�/�?)t��h
�D1��0@�<AaSj^,(ꐨe<����NZPuF�h��F"������T_j�g�b6��tL��?�zbΌ��������Yc�Ȭ�����s{lO�#��*��2Z��Щ�On�_�fIG�v��u�H1�����?mo���fj����-�H�����ٮ��=�|�����ڡ����+Ƶ�Ƹ����Qs�K��=3���td�ٸd%=\�2��"�ㆅ��M?L� ��d@M�w��{�@x<#J}��Y#�QYA�V��Z�UrV�缽��t�7̷����u�$�5G�ш�P'�Dx��s/��������.�Qa$���BV�;�Wj�J�M�#;��������F#(����H�α��ۀޅN�(!�*IglAڧ��۟��[$`�D�J�/5��r%�ȑ��
칎�w�Q>)c�3X6�l�=��	��[Ryga^-})����ģ��R�翦��}��OX(����.�������$�w斁�cFy#���jr[����SW�I4IS�ݼ��b�@j[\p�1���]�f_-�`��m�C�{zؽ����q_Qi젘ZFn.�!�Y�|���>aeV�������0��7j�P����i(�i�r��M��)�?&���t&bkB/�MVWP`����#����)_6��b`s���\��hB�q��ا��Yx�}��o%?Q)n2���P6������k�M���$fb����Ǵ�ﶌ�X|��_��ퟌE*Mt(���W�,���;rP���L|xhYA�E�����5�.��L��(=��H��]K����u�1Vy��\��K��H���e�U��Zf�Z���Z�H �d7��ي��e�K�����I��r馆Wi��Tct�A"���B�C�T[�NN�k�bY@b�=�@��y�ɦ՝�Z���ҵ��$��������⺦p��ďW�f_�ٸhئ�e���Z�x�*kŧI����b�.u�g �d6�O�ɞ�	9b������iIP�*:HrEd��

�Uf]>������CeǅFcC��$�ގ�)uf�P��ŭP��Z��4P��$gs�j��:|�R)�d��+��p��
�׽P3��������>a}��uZ����|)%��M�ws^�Ӂ�^�iq[!@�w�o��d�<�Fh�5�M4��Ϩ���-�Q3���JI���kvA R���eȄ!9e�����oG?6&����;f\	1F�g;��Pկ�ߔ`�����0�ň)R�b�ؾV������;��dX��t��TS�\�
,�p��qĚ/vAX������1E����tl�Y*Mo%5�w�����b{0+��u�����+U��I/ōf��HF�Mx��ZJ?�����Km�/���L{����=P���su��6��:L�<��gA��e�J&(A��#��=@��1[Ƌk���'��/�j&�v��h��. ڿ��5�$f����Ĳ�d��h�In��'��k��Pm���G(4��kY�v��
���"���n�B��1�ͮ'G�]kL"�Ǩ�^RǱ{�!/��0@ ��QiRF:wR.�T�܀o��Y�L�����.���f�ͯ�����X��{>�\�#�`���ڤ�:v=z^@� �BB�&ө�Y�H���H�Ӟ>�7;ߕ%>Zm��;�y*ݐ�G��.�H��cY��~D�[�Qƕĩz$�aK�dM<te���
7-�kN�>�\Be�*5�h�bm�a3� ��5�/�t�)=e���������D�9P�3�Sgw�M2"������L��]�k9������m�ݫ0Q]s���
�l\%�;�7C���S�ܚl�.�e���Yؒ.9s�揺�Nŀ�rh�ǰXC��mj�C��35�q��D�#��-5��a�l{�6�R��l- �W0.%D�wT��ci�Ig�:-��/_3ݵ�m�A4x�g�v<mݖ͉���n|X� �����
�V�(�Ee�[�F�tݼ�;[����L��Ɏ|����u ?y����ϴ�>��o�]���Aq^r̬N���5�8�I�h�c)%py��6���;!���i����(��Yzp8��jw����*}Q��#�-E	��T��������x�hڑ2��I���.��l�CwH�4�'B�9I���B.`Y2�hH�^�M�L�H�a+����¿lFԽa�#�.i��P���~t�알��� ����LX��F���͈��6�ִ����8r"��U���0�ƕ,�.{�_P��t0�B;Vx=�RD�S���XZ/Cq*�z�%��/ݦ���>[�-�ߌ[É��^X�33����������U��z�J9���&�3�~�U���1�['����7�2N*@�K�u�dL��vR�rτ�*�U ��}�f�b �6+�u���4~{E�y;6v4�L�k�M:շ�Q���D���� ���+�������YO*�(F&|��sz�8�n�f�Z�o|�7gL�Ӄ�����5������2q��c���m��K����Z"k���@�]l�a�o�ң���c�t�v��̆;#���v�FQ��2�Ì���|}*<T����`��G%' ��3�h 
\B0 ��B5�w�Y�K�.qr��o���Rt�Y�u�v�R�]��>�[��&ۏFN,'E��*'��b-��E�J��o��&�.Y}�B#�QPw�޾�؍~bٗ����eeU��l�㪲kN�V��h��N,�t1N$���*j�p����)k):�@�+#�E���/&�^�|���&�R�ndb����E1�y���3�	��Ptʷ���	�C�t�#���\O��r�5U�pE���Du�����6lyilJ��Z3.�S��	iZ��s�Xt���0Ud��Oh��Pگ��1�� &�'Sv��^JW��
�6"�<�����f[Z�,��=���➝o�h���.��#�v1�_����v��`�d�v-�C���"%�_���8ɨȫ�	4�W� �E�U y)������t�E@v;~�ʎ���qyk�AS�t��q��L��/��S֢��I|	;���+Q!�cr`8�(�����Ys?�;h�6U���Tp_L��h~����P2q ?�U2��M�l1�.�*v��F��f��������t`������[�(�@ �xc3`N倝%�ev��@,v(����~�P/�5�'���g�1��K��@wJ21�&}ۣ�R�j�������O(�j���W�-Q�xe�ջ��d �l<n@�E����V�0�(�]m�X�Tf����:W�V�7[[�S���7�^.O��H���
�nP{�d�z?�]���
�#����KO�ڦT� q)x�����4��M�b*R"�j<"�VZ(����z��i�-&��GLtN/����@���[�j���^�mE�zX����tlTB�^@W�r���*�2�X���h�f�eq#��	�]��!x��%�0F8���d+�1]�8�Ϋ�H��	��&o|YI�<Z�A���@r�:+I�fs��̈v��X�o>��Ir�������F�v����y��w��n�Z�Mm1Yա���rŨ�7}\����`�z��M�����M}����3�<"����.�f>�܌���,4!f1e���s����eg�9��?��2��-�P'2�ރm~w�o�����������ꂍ�"g�ᷭ�y�� >,fr�3��Cj�S�#nO�t��q���[^���j�1�ţ��"�R���n�-�dH��1��c̼�s_gs=��2���\.jq�F�$�$�����<��ڵƎ�FO����ş�� ��@��7'/>㢘��ҧ������-bsF��� �jF��^$�g�"�ִ�~��U*�B�s� �����;�m�i�mO���~᤼������Cvk��K������(��_ʎ�Tc��B��2��P.�@�,[�:tK��d�z1Co��N�b._o'�K
2)�q�fZ՞
>ȀWx���5��T�vԪS��:��8���a�#�W��h��=/-�@xL�>�ci�J.z��^2ft�?Syڷ?T�g#��+��"�SاY���5x���ZN|`r�Q�å7����"���yݱid��W[�a�v�����k�!&�&�H�"�.�\*����4>)Q(�I�z�א�Q���<�N[-S�4�J]�r�X�������"�h��v��Q �1Bc�C�^���:�e���������n�L�q<��'4wNgZ_�Խ�8�x��F�@Y��L-��eo�1q^L�I��*0��o(܆S��ΦI�Qn��95�F+������nPU������Ξ5R,Q���$�]����^�ށ�=d��xL�~��Rý����޽���^�G>^k��wG�S7^=N���V��M>;�ű~$tد�p�'p!O�@ۣ�P����ƕ��y�P�gM��=������j�B�3\�LIOt�.��-<���RTa��-.cƋ0��
���[��f3�i#��Ef]tq��ݻΤ5Hu�s��;C�J/5u�tp�pz�mY>C�ܢ�������O���i�ϾĬ��MPbbP�|�J�YKp��bsm3Þ��W.����1�_�y�&	gh�M�L�@T���U�"1��ϼ�:2�3{0"�Y4�hAk��=�5�oJy�+�E�|���$�޶��.��-�.ߪ:@�!x�SH�_�?$��j�`<�����S�b2у8|�ֆ�6�"Ȁ'F��X+��P׈ޮ��!��>��XbdҼ��"Ħ�	r�w���+f��?g��DIs�8�k�#�6���܀���|),�V�z[�<��Y�#�]�﷩.@F5��QA�Cq���e�:�,�:�j�Vmg���g���o;�p��K�x�nLNO)_�:+dGb� ��Pʼ���Ҵ�Me�	8&���
�сu�i��iWH��c���~q+��<�?�daY8��FGe�@>��;�>#B�f4�T��)6M���_\�c�|
�l����X�KKq�Y�� �8/X8�5�$B`����L�P!ː���
�/Q+u����q7/`̿é�/j27�%��� :�ɓ��\��N-�Of?o�`8�]S,�'��]�0�Asy_e����Ic����t"�MKv��l7l�dwA�b7�u�zw@��鸬ZޡO�T�f�I�c�W=G���$�[�d��X�@:Z=X��r��	^��(ǷG���3y!�>Wӯ�(�R���-ȊIk[?��V}*�+	��p�Y �Y��0�]��rϩb_@r����v0
#J�7rg��+F���{�������23Z����wp�i�J�qQ��!ɑ7�
�/��kRg��C�Ҋ��-~MO�D�[/����T��v�i�PV�uf�v�6[��t�;��>݅�`�P\��1q1�t�	���*�I&�7�S�+���45]?*�QQ�-y~��1�Q������=:>g4��$������2Ga���pYqCӝ�_�mr��,�e����U";m�5�*�@%�Bs��C�r����C:~�P���4���W�z-9�I}�:F埴�^�O^+/���R?���h\W�Z�Y�B0��I'����J�~á}��"���(QV�O��R��? �:������� L��w �1hN5{�ǀ���E��Tvo�Q���������K��7�s`Ğ*��Y�?Kv�8MY�Tp�ɏ3KA̝�
`�S��"YeI�?�'�Ĳ���q�`<�t#��9'7U>t�o��1' �i�Pu�J�������ȗ��\�蚗�7���c}���F�j���D+9��M��F�x���c�,�0Y���#�U"H��h!��Qk�L�Jw
�ū�Q�im�m��Wm�z��vv�ɉkqS���n�����)����h��A9 /ȷf��TX�:��)�2���O�8��߆xq��ɷ�X�O=�������;/w.��f)
$)��'|{�ǩ�z�.|�%�%��� 鐏`k)�n�e��U�oHs���q���TGW5ϡ�ܼ�e�~�\�I��jKNm��4�����c~�s���^����od�^,E��3�'�B]��N��KV"m<#��u4�W��Ρ_I7,�w~��J���L��2�,�^�����!���`o��h�$h�i���H��d0����P8{ꗐfX�\.=d|���g�{%��ߒX�܇���o����4>&7ш�oT��[�yqӻ���*1 t�3�������k�.�CK
����{���Q`gg�X�2����tl�#����^�ӑ��g�)�$D4��[v�A^����{4 ���=��e�U������#!-��,��K�`�B�B
��82�Q�"���۲�����|YQ���F���CeY��*Ѿf�������8�Dv߮m�p(���ڤ���h��垕[�O+��}�fܺ�:��� �4\����F	r��t Q^�,'�b�%,wVvQv�߾�&W�M5��1~<��2��k�����"�����?��A6��zPʴ����?�� ��x~�->˃:.�0��>�@D��L�b���7G�RC8�"��!^�R��_:�j?U�¹bdo�?��Խ��eC�K�A�֞�V����-i!}:�b�� ��\b�i< Ť��M�����4��Ġ�=]C?~F��ٓ��
Y-�ސ��ebK�$T{��8��Z����;�J��s�N(e�����p}0#Uv���I pM���(/�Lh�Zфm���:�ZA�Ψ������n{�eRn�x玿��V�t:1�ʈT&5H>U��&�������H�����݅�i����5~}�J������&���7��F_)��(Ω!8Ŵ�YV{3"d�����[�e=��5�PU$$�QQ�Y<r�
��'q���೥�z�� �,�!nRg���\��_^����C�@^-B4d��N��\VN������.��
�@�eY߫�I�>��2��$�vٕ�㥯��*R�Qx Zj�~)��	�+��zG�5:!�~�%]
P�+�� %��ѶY�?�HhrC�^ʵ<Nd#�D����|��^�a�����Y�K��S�iT���[��X����7_9� ���'Ĭ���y}-���̡�8`\��qHգ��)�Ԩg��������&�f�4����T�����P`'C�,�]i������~O }��./I��L�d��|����zX�� ��^,��ծ�ȷ���~ڕ1����'𛪟��c�D67�iɈ�DUo��!�qf}��l&AEx�ym���l��3�,
�kff��h��c2(�lk4���N��N�T�g7&��ێ�� ��{^�����CCL�A<�P����qMX�;Ü%�(����=�L�׌d]˦�zA�7ꧤA4��ڶ�����Fq���#� 1�jc��r�~$����tk�F�cj�M�1�+Ʋ�T��d�>1#�G���4��`�څD~�a].�̬G�Y���1y�O�$�����������R�X&��Y_<tZ���5x��NS-��ی2��J2]�1	�D5��/�z��k�)��k��,"�ui_5����?��E���%>$���e��%�a�X4� .ǩ���e����*?�]��t�Lj7v��;E�<�@��_A�Z��`;�0��d�OJ���������L��V���<Q�o����T+�O�qg�C"�����T��J�Xts����}��j��e��5�|�f�/0����T�����$��-�Q���M"�����a&LX����㤛�f`���$pp4��0w>�_�)3(%�F
6,qw�ƽ�u�̆��\�S�X��bsK�
�d�f]��ӄ ��(�2:[������sgmr2�A������}w�ڙ|"�\��9����=�k�.C�ZS�P	�ʄ�����p�Z�#��~���e���?����c�!U���j�1=��3��p�,^)���9��\0���l���[a�͍�<x���]���lN;�k��kP�@��LW���O'���Qۄt<?"}y��5W�1�j��&�a�t@�7������YyV%�|6��qT�ƕ�������{��bU���QC��
����m�0_R�M�r_�]9�(Đ5�r����k���j��ܞ!��3��[���LK�j*t�S�SI�B0mm�p �+�_	|_p;#Y<#/������{g��0D�o�TI�f�K�O\�~�|��=])��S�"Q1AuwX3©:��_��x�K���k
���2�mF^����d��M�
nZB
�-Al�п�V Ǜ$�����d���@X��{Mv!������f`h ̽_;� �w�2�uS��� 4���ѩ����i��{y��vj���uG��oG������@B�G�Ζc2�M�Qz���O�]>u����yX�7r�Mz��[�Kd���0�jq&��O�����6�����r�m�?��;�A9�KYD��钵Hm��A�r?�P3z��J���[F��2�;�
)�4d�����B�~��U~��Ƕ+���S��~Zh1�c�5J*"9G޾Y�ș$Ɋ����ݎ�q6f������'B ��p��~��[]�UB�Cw)3�O�z$$c�X����b��N{x�Z���mˎ==M��BM�F�@3ę!&)���ɔe�1�-�P+�ގƵ�+����J��)6	�i*�c�����aR�Ax(K�E�/�fcfo*���Ԥ��1אM��cwڿ��s�	�gygC�Q}V7�|��Y;G{: D���"��0���;��E����W�)��*m��<p�����7*W��;��2�����rE��J�3.��ҹ��H
Оt6��+*gA�o�\��2�p�p�}O�):��,`����5���J������sR�3E@6��R����>OG֤�֌�Ev�A��TfG�-����Gt���-R9���.�`����y��G��) ���:���` ��<�x�}�w)RT4�h�31�(�N�Wg���ߦ�R}���j`z��+�l�����[��F�)������l՜�夔��d�e���H^&L�������\:X	��-y;X����4�Q��5��h�56��)�AZ@�N�GJ�D\(�*´�>���#_Vy�e��*&Kd,XR�a���Û�wH��0�Mr�j=�~��o|k8�������fO�B���C��?�Z�ԗd r1��ǩؐ7R^0��7s�g�� ƃ�D����!�Ft��j��D��ܘ����R
w�1f�6�������<�!Cn�p�Ƙ��w�)���ꝼa3�����X�fb����}pu�����c�
t_�� �\�s�h��.��4�7��j�ww�i��lG���vп����v-��cC�
�ռΡ����Gc���~N�=����o�הD���	�	=��p���`��\9~G���������v�	��.A[l�}@�:mqA������	p�o�7X{����I���W����5�}r����~W-�w]%Nݡ��G���hHu:m��S�Fŷ�<!���=��� w�Lز3^�N 	������I�Y{7�)��r��H۠�5��Z�>�+�uЦ?�DM�N��0E�?��F�I1�HY�]�f������� ��ͪ$M���P7y����3�[L#�h(F����Ў,����We�`X�F i	L��[���(���%�~��Ξ��XW�`~�`�6b'&w��	��C���a��_��5����j�-��MK&}x�4y�a]�#�'G�EC.=�Y�bG�ˋ1���2ǣ��jy¬���ƹ��
��0��ȸ"����So��87�Pm R��SR�� [��@���tW�2Ib���OE-	��>E�.*%"j�U�A@-�2:km�P������n��I��f]A=��1�{��r���h�	��V_�&����ܹ��Xr;̝jAw+�ڐNR����g�J�8Px%����CQk���.	��;-��f�{��H�&�4l�����DL�O����]�Ú�["(CC2ﾃ5�:�a&@]�1��o�Ok��8�.X�9����"�6��hW���s�sy/-���ѐ	3%�-؊����[�m���GS~w߆�B[d*�H]@`f��T o���H�@��Q�<�>TgIe���~Z[���\�TxΟ�? ���@���'Co�����<>��/n���1upPR�@Z&e�� �y:N�����*��:ߵ�._*��5y�@��nJ�6Ɨ��Fr ����
)��a�?58H�)S�Ȇ���֣��p!⟦zj��Qm��\a�LE�oA��J��g[�Jȼ�lH%x�t�����2�����\�z��55�.̟��vNگ���?��`�����?�u4X,yU��D��`ۯi+�n�t��nԓk��>���]���C����v�4���ߴ��_<�
�D���J)J�y�|���e���z`b�5���*s��KK����n�7#�N��ő:Mh�2nM��<cNC��!4�i� �W������cw*e���4��(_�z9�Y9w���KݏP���wv�VQ��X��Lq�m�
<��dق�s��@t���LN�UjF��+~P˙�v��dOusg��ʠ��d�6t� TY:@{��-Pd"�B�@�Owy���'n��?��)m\\��[�f�n^8���'6�D��^���kfn}�ߣ���G)4B�ڜ�q'1Z^�=���ŏ����H1�1�?r�#��x�K	�V�#ʊ� ʕ8�ꚓ-=�5�9;{匧�S�A�[��0={)��h��
���� �%��M�YW&~ه漹�*�ݩ{E�>��cu睥]N��vu�������i�������*�Aw�)��cMO0�|H�|T��[Ut�`�������Z^��s-�j�O����ae�N��JX-X��ǔCT�QhQ��F��զ<�鬿]� �u��D& ������OP;n��>�Qԋ̴�b�w�`-�m4;w�Fy'�ȁ$��t\�� -D�4�%��{�F��?^��N���3�jf�`\P*?�oy�m������+{�����ר�{l&zAh�5'BX>v�Tu܊��k�������,b�.b�=�+�er����a)�~���.)�U ��U����W���(\�J#z����"�,]��
ZS:g�n�=�<��Q5�J_Bd�G�B�w
�r�������RO��� �n;�Ptzv�L�;�����i�=;�h$؞�}sYd^m���ĉ���m?t5G�`ntD[���P�Ad�^ a��9yr
d�,���Z��e�����C|�@Z��O�RN�"ǯ:$Oe"��ln�Q2 �(��G5ws$D�łb�2��X�V����)6��%��UC�/�a1�R�H<WR:}��ۈ$�Z´\c%1��ڼqyW����3|��(mDi�LI������%��w�}˯�V9���j
? �/]�V��qd���\[O>AE��O_S�����k��)O^Zj��~oT�5�Ѝ�H�+�+���ȕ�Մ(VM��+$n69�BR��,mS��\N%XD��Y�j�G��Y��aay���I�f!-4����v�{#��ys�̃%��B5�����4��#�����Z��>�X"�=�z��C�e�5�B�	��]@7X��"�N���4]�{Bs�[��ɐЭp���&;
�0ۏ�K���Z��n�[_�eOE곕Y��ka�!,�5��X9X��Ӏ�#��V{[���}G+�6R/VU�XEa$>�Q�|�'2��D�W,16���)��ڍS7ZW�N��D���px�ˬ__ W���B/�%]�Dk��i�tI�W4��a9w��z,CC�,.wW}�WM�����;kr�4�3���L$C��� ���!ȀV`4��z�B9=z��\�}K��kmfr�	��Sϫ_�d�������K^0�ŲLf������Ԧ:Q���~�����\�D���OzSU?��WկO��:^�ߙ�-���U.cቀk�>vwo� ��ٚ?xIb��Fy��FȉP�����_&f{�i^�	7+*� �A�0V3���xQ��a��[��d�p�QH��fT�%�'��u�B�^*�O߮���Pg�n{E�WUu���?������F��\��#��^��������YFա��c�����^��e)�W
��'O(�Z��r/^T����jțۘ����p��d���V��sf���2e�]Nwb�S�S�'����r�cJ�ʅ�?��l!���Z�#Fp����a��ѓg���h���|��j�����.`�)jd�ԙ�F܆,l3,��LJz�Zp7�}s�\T��Z/J�*��$�4����8{�wo{8��3�Wv�6��$r��Mz�f����Z��ী$d2g���BZs�������s��f����M
�]�'������ڿؙ�я��'��t%�ڡ|�:6����l�%��g�i���k�tS��
����0>F��n���T�m�2��K-hH�ܨ���(�Ǆ�՟1�G�%����Q���d҂��t�S�k*���=q$��!�LX#1+T�2j�0M�� ��H�l���XsC���Ez/ތ�?<)��}�bp�d2���Qv� ��6S�� ���z����r%�-c��a�ha���(�9oFO�V ԏX˾���`��b8Y�࿚p��� �y��*�կ�+Ԏ(%�K��ʴ�E4l�<��R��~ћ=�ރ��XjSҖ]Df�С��e���fjx�֙����QU<��zL�l�ȼh�a���*I������ZO���^l����M��D������}U�C��3/��U���c#�wy���W�1�y߄%���;cm.P���@vKrM�:� �&�Qng��� oUG$;?��8�%��%�.zL^%"C��z�:=��kN�����	�D1�$k�����|��A�#�4�L��X��L�NN��͖�$�t�N�O7�R��7�.I1b ��(k9!n����$�Z��A�r�Bo<��_/������E�K_G�Z&�>�3��2Ilø���Ef�j.�xx�m^f;$������n�ꌗj��B2T�����E]&t�h��D��:$Kd� q֡.X�)d�`+I�hC��>�%o��u�r�\�ՂJ�Ai���p	�:35}S��7*""�Q�,(Z� ��ԐY��V��L���<�'T���R���7'T �p�e���,����D�����F�}��1uuեĕN�j޲������x�jQ�3��ڷ�����6Y04�￀��z�7�E�}2�Z�Y����9N# zO9p(�sV�:���s�8;e\;O�*Z�@�J�>����ر0R�q&p�(U>�:�������@���������@��F�_vT�XZ*�,]ݔV6��tk�y
G� �_:�8�|��I�W}�V�[l�U��,L��#~ݻhj���N��p7��o��S`�^&�x)1���N�;H�`/���e��h�~���0c಼o �~�_t'uv�y������0G,=N%���OX�H(�jо�JlS�=����ᩖ�v�d��)J�oH�z�M�H?�w�HX$��>,(�%�%~J��B�%t��Yot&�q��0?����ρ�ɹo8��y2���l��0�r�Zn̨P��.�)�����C(n�v���n��@u����7N͝UzL�M�~�R�����oM(� e�l�,��LP .3tnW�-}
 ��y�Ӕ TR��XL�����g+�{��\ ( ���
2�^էɈ�5�ɀ{��?-���G7�����7�S>�?��;���k�)w�zq!`���rt/��UYx���(��=m��a�OO�Fٔ��	$��v�4�㚥v'.7�gψ�|_��|#��xZ�Z�Z��Gw�r�!C�ճ?��U�q�B�fR�A_���K�#�f��o$�(tO���M�"E�xA��7��8LÝ�z��VҴ ��.�X��~�������ߚi�������%(����J	o��pUR&ϖ�e��'Ąhk#�.�[��^��-8�"=�H���o6�g���O ��a%��^cQ����%v��VN��	Q�h����b��U� @�8T� ��O������[���@�eO)k��_�S�^#��ۃ�au#�hr�%�Q�x2:e�v�O��՟�Ɉ�&��(o��ڍ�S�B���	kQ��|�n�a����l&O����d�����z�� F�$���Y�[���Ҷ�7���~'�������@'W'N�:o��y�ha�)���KT�|d�5vl�؜ɵ߳Բ�@x��>�}�L����Ӏ���R���#G�5uvE�_O(��|��EP�:�rU�����$ :ak��&�>I����O��m�F%�o�3>JP`X�:�⩍����H�G�T~�2Qe��S�l{��n�ƎH wT/�j.Z������l͏uwc����$�$�vDQ�+駋^���9\,��4��$��Ӫ���^Y�b&�@Ǭ��bLtN��)��Q����
Z��Ik~{�d���{�"��"������_p�T"��Oҙ�)j�<��B 	�l���������W|h@n6n|Gm��>��k�
?<aj�ȟ���޳
r0yhqYU�-�߯�w�F��������E����Gl%Q�d����juO��jPs����+t���,;�����:��Js����	6r�	f��#́�X'g�F{�ې���Qp	ی�R��:�z��}�H�n�'-Ų]2Z�:��:��m�Ч�1n�G�aۄh�s� ?m`�9��c�
�V��#�q�Z�4'P\ב���C���-$)�=S��܂�p���n�����i����'LK�,7���4|��NV�<����Z�]9��q��fn/����?91�-����87��\����w}+@�_~jVđb⩁x�'�ܸMF����d��uK�f�`uռ_�E����/|�����@H��e�U�����|Ǵ%�_B�Z&Ń�׵jD�u�q��{�tU;�Q���ެ��]�al)����-�Ef^m��j�0��,�6����\�2����t�����*.��)�ʎ"jb�- I3�õ���!�_���f����S��d>M�aU��&�#��L�Z�g�J�%�����%�>���H��s_6ء�"����d�S�FbC����lB��SVhp �^VG��I��bNARJ�����H�bߴh�i�\s-�_v��Ư����{^�T�|O%Q��������:FT��8��n��&6	�R"uv�>s�u����6؟�T=�א[�3�l�a�}�}�ݪ4*�yCZRN��&e7�4qyxi�±J�	 ��y�/�4X�[O�p�Ω��M�q�8kRk{�C����gfU[{�u�����}��׭e0����z����ku}$F;�4��(qr�7�Tٍ�؄���0���O��JVu������WQ�X�v�bH�mIK�����\!v��� �#��3ŗ+f�j����r�D�gto�U���^A{0���%F���G��$�P�MÀ��Ҕ>���4|�6�!��ˬ�81Tu*[�n}��2�FL�3�_*K�1Up@��V�<~j����
��=�T)��~/�<�r��x�hC��$�©|���o�r5"�6β���v&z�E�W�+�=��C��<��G�6<��Q���&�0���iP  [���}(tDA�)�����n<��}R>�0[�]9⡆!a�y���~7z�׷��m�*��bGEH-�c��U���!ܧx�D.Bu���$c�F\���\ZXW���%��n�O����>������,�74�}2��aVu(9fp�M�ɉ��}�����(@|[���i�'����C���6���?g���B~U�VO�M�r�v���t�*a�;<^!�d��V.,�;qb�^@.���a����q~�a���H�Ouu�5W m�Lw(�B?���7�H@&�n6���&���d���o����5k�*�'�Em@O�ԭ��DEȣLD����5���n�i��u:���6o'V51}H��1?�=�ɪ�yq�����md%qB��(�-�I���#a���!���Ij�z�4}�Kf�l�rft�Y �!�6���O�ާ�c����Λ��W���M�#�ȃ�z�`[s7�XT0CT�9`�0"Ƥ��Z�]��+_M��(���f�� XF擒5U�Ԛ�GG�C�K/K`L��o`M!S�V�����\_;o�t�!W��~�0|):$��ys�p��<	�LM�p����ϔb�Z���G=V7W���Wq������o5��ŝA�6̎3�����������Y��{�{�>�� �Am�Y��OR�;���瓨����:'8;�4�fQ='���`��}1J�;�ԗ"m7�ځu��-*�e�|�lC�,=�"���P��������+A9�D��LO��1s�а>������]Y�6���y��Y������{zìk�%3 ���}�!��1�i��3��g쁒U����K[�'!�%p����1�)����\|��ҩR#l�#�Y��l���m_O��Y�[��h�O>u<�^��T�C%7q���&}��dz�n�I�L��7���Z,�O�PLX�b���R�I<-;~��V�כ��m�R�g�f�Ri�#3t�������K�y�N[�N�=���^��:M�4�2S �Ә����V�
��!a���vgɒ���p���>�0䉊�D���������؋1�44�M_�E���5B����H���xq.��,.o�.#�s�x��94rP��̲��<$�.�����B�[2ʖ��n�e��r��w����v����cM����@����1�vFz��[�͐zw3�v��^�̷�K����B�Dl��u�]b� �n��c�W�,��FEZ�PU�^o�ӯo�V���.����P*�>j�0n~�;JU�)�1@n0d=q}�>��h���8�a��XݾR��r^�WE��&�/�{6��l:(�L{=�eA�w�����i����b��rZ6����m�l��Gd]2j�d-���;5�wq� Y:�\��TV�Y�3?�_�js����|��]�V����G�Y0�����몯0f��茿�({Շ֠є;e`���;S��쬁����U~lmF����?��ǿ��1_�6�
t�zUw%�`��S�)}O0%Xy����䐩��W���	�-�ȿ��x���j��c�%q��-�Xs��?�#H>[��,-���q1��#\�x���r�=r/�3�[�2\YS4�E4Ws.I�V�~� �9�<ϼ�'6I5�W�|ap�?����p(Nzt5�h�L�V�P�sb��2j��8��U���ߑd�p�ζ�]�b3��>p7�<w�g�N��Ζ�?��B	��b�b]c|��J����-��X��j�s��w7`LE$�(��{�s�'�y
�:�N3gO�e���<�F�F�3��s*:�cv�&�|��<jk����Bn�����ѿ�1U�O���hN��e e�A�oGv B�dY�N�y�t1Kv�ϥ��>o��v���7���hȊ�٦�;�{��Ã#7j������80�������7F�D���r��.3~m ��T��/�'h�$�5p5j��5�������$�Y�KcN�%�;�O�O	�|7�+�V	rH+��۝ԥ#�;Q���X�ͪ�3�ґ�	)��Ck�My���3�(�T$�8���UM��,�Y��Wc�����>�Yn�M��vd �(�����=��[��
�<��Ȗy�
%���BJ����O"c�*�r�� ������c<J+m�w-�?�W� �j���� ���\-n,�?��5��O���(wj��;Fy��Tۚ����\�:($
1m	D��X���Q���k`E<�٨4j���P���M�~�쏃dh�7�Q�gE���3�����0�Fꡟi]΍F&'K�@�y���#_���0u}��Ę�F����E�7��"Ɨ��b�93˗Pڑ��M.�%�h/��@�+��q��C��3i�e�y�A�q@�A�`v�!��M���g�cȜ{���$4z�q���׌�dj�Sf(C5����Q�X�x�E�ځ;Y��+3�u�\&==�f-�2{=�*���S�)��hz��j@��X� &�XA�4�ѣ����U���}���TR�E���<��/���(D�S�L�|PN�)r
 4K(�,N4��}��������/�J�zQ_����KZ�~�?��ݠ���ۈS�x� A�%�'g�xP�_��=B�@�[��ϯ�u��p-��z�����
;��1�H��O�+?;�?)N� ������_C��D����VJ/Q��E�s*8|C��-��j����aY��;���j��A�]��J�c��+���	� �5��w�͇��[��2/3�j�]�XJnr�BQ��ID#�#.�Th� �^fD�f���k%8�Ux^vRsw��S-���N"Άp	�kt����sct"faS���"L ۊl�!�+,QG��a���vd�T{(�J�s*l�l�<���:%C������s�j�e�%^j���{��&�J/�7I�� |��;�њa];�O�V��,5��[��P�*S r��&�'���yL"��?/ڋ�'�ٮ 0)�Z!d�b@a�(
���+�%�����K����=w�����&ys��h�5�8Ψ頚w��a�ðלȈ8�][UH%jg�mE���?�[tU��Dg��;�K?��kdn3���!o@��)	�4�;� ���狱��7q-%K�!�<�����Q��3tu�\��"�r����gpk�-�(��B�[u���i堠�_��x/=Ʀ��5�(V��R0R�)�#=_�,*r`��҉ ����zc;�4���7�
������l�hu��}�u�-���_�������t�O��X���dR"R��?��S�>�Ż��"?�}"�����ݬ5w�cw�P���5e�z�����;	D���]�?ßF�5�/����5����]���;���;`�r;����r����������.4�F����{�Zv���bx[�
<��ȵ�wlLи b�wkop��!ݫHY'�粥u��9&��J
�h�N�����8�������&���fC��v�P�2g9IY+Am�����D$���k&��|%n��m
�J�2�Ou�qVt�eB�	֮��D1���3h,�U$��q\CX'�����ZF���:6��iœL;H�vc�c 8&xw��E���r�'ni���r��y^�#NK����TG����Ȱ��V#$1)6��v�j�	���^&��/�\ j�҇���b����)�>��X�d�yF���˂�o�S6]?�����|H��̘?D��{��;�-ON�R��xXW���� aD���U��#u_�cwp�(Gǐ�v�l�\��ڧH���hr����I�b� (��y4���)�n"Q�Tudٷ���r�R�����f������2��b���C*�?��(�O���,��q��Fh��媜������-pi]%Ƴ]���͉Կ�?��|���Au��I���-��V�J\v�е�(:
���K�OE�m,@*������Zԣ��Lq�Y��r*�m;u%v6 ��`y;���7�A���1��d�K���X�$�H��
����g�ږ"�߄�s@3�����gaO����PCo��[ҹ�^�}̅g���d�7���|��]�+]B��縨NW�$���7�K�����P0q�:َ(��zi�i�ܗ������`w�qC{ҍ'�r1Q�GA6lp��Tq������*�}�7��T 8��9ӓ�ג�*M� r�8��tU�Â
ì2�Q0X��	���;�ftLx�ػ.j���ī��bS��Xz{�9hҚ$?���i>Ϙ;�0���?Y�r��@,�6)�]D�d�+z���gy>]-E�M����Ԯ5�:rZXWa�����ԛ���]�}���uZA6?Lm.���rͺ�;���8��Ӊ����E8½����.�]i�dC���J���b�2�k�#8x*��t�e�4�`�E�P-~�q�}u;�U��Z��/	I�v΃�>���I緲^`"����XfK�� �����9�^|�f(7JI���\������ެ=���f\?WG��:��^V������7�U��n�6��P��oiJ���k�3lk%�x���V�)g����Q��H�R*��}�fJ��v�:�������1�1Z�%h��9jǲ�`Wl9� �p��C���g�*Ӣ������Oj�f3W�5n��|D`.4��}�g������F�6�7�4X	�HNP��v�꘻�t��b��;�j5���?���I��������|�_��CE!u׊(��"��*f_Y<���i�=�^G&(�?R��@8|���?���ה����Sٗ� �uG�����0<z�1	��-��e�N���sބ9T��)��|^���>�T4%*m
@�'}�c��u��N�Z���/$��:j��v����y��b���Gsr��r͠:`��L�}�G���TT�9��cv�*�c��fQ��j�Ѐ]%x����O5��Be�
K���"�A�П�Eh��\�m�n���hI.@�В�:y1O�P1�Tg��&�P����%�E�x`+N�9�9�[4Ie�Z�S#(-�_1��x�e]��rA���E�9/f��G��@���s�����E��� A�M�����K���?,#rX�x�Wrf�Ɏ����O����k8EdX
��(�sZ���q0��w��Ph+e�ex�r/�҉~�Ϥ�
�A�S��H,�SE͢�G�J�@H����U:��f+�}=lp.4=o��0�8���(�l�G�*��9�E���NV^��n���0t�vHK'�g*�E����J�9$�0�ťĽkN'�_��sw����B�����f譒������_�u�&��|u��f�j�nt��y�`&ڰQ˪�כJ�ðV�>Y��F�t��`�&ʪɋ4wD`���`��� )D`��e��d�U�C4�u�g����)�r�䖒��.�#�䁮���ۿ$����yOC[G󚬀/�
tl32�.wև�tX�j��>�y u������N�q�Y���3r�K��;N�&���k���7w�2Y�[��u���o�/N�H�F1 ��3O�sZL�].|�.2��!�I$w���%�^��'��Σ�Sg��tm\jkq�{���(���S;�+�}~��I4�x�YLu��H^*H��pа=ח[&Q�!8���_��?���ʖ@i|���*�f���~���!�C��%+�����d���f��!'�g��]�F�m���D�6�}���|�Wa��L���B��~��qWL�D���%4�6��I�d8�]��������D=���"��<��y>c��Ҵ�q�L��?v�I��]��AE��UC╯dF�i������I���֮O����~6.6a���>��\���/�	 q���]�$0��; X�$��l� �5SHΊg,�T7�ֺ�ɝ���C�9�WJ�ߊ��wT%�`��@���/�N�����ܡ9��וy�R�@u�6���=o��]���h���7�;�w
i[86V~$�OO,��şyB�^��j�,�V{���	� �s�?�D�� Z��<�}������4>�m/�zC/��闦_��Us�-X/�z�����ØtƦ�FVE�j��R��!�S���)�-��>��U�������w��)w���4k1�2���ʗ�0�{&e�;Y��#]d��瞈��j�g�%�
l��F���pH��:=�A��$v�V��E��)�aC�(s�jH��[;�o#�����G�1AW?�w�(=������c�`ā鏈��>�J`�VtV��J+3��/�o<Eb�$�����4�O��*h��)<�l6�H�
]h�g:ڈ�T��!�Ȭ�������/�*��_�`�4A�-m�B��I��������¡C�ʦ�r�X�F;2{����_!0GҤ�����2�,>�]��8��.�<N��w�q��(i��������7�)v# ��5=n��*�9�c
G����yERO�����ɮP9mo^������AK��(�^��˜����1�G�s�X�!���[u�܅C���f�����ƙ3|�A�-�-z���^�D:�z���njz[��_�j�@X��M%)79ّRs̔��2y
#�B�c�N��5�1
�d_�5��'7�Q�x�/�-�~�c�Q	�5�iT��!M>�\_�/��f��dxӦ�.����`u��X���ӵЋ�<;���.<骒�<���8'U��3�X$� ͺ��\���f�r_9)�W�[�����+Y�¶`J�=,Ib�ӃU2A��TZ5`u�ֵ�s��ߵ<�m/(�uU�����a���h5�d�h��l
A�R��4Y=�7�ܓ���7�xV��gv��������l�������%�*��gV���$)��=D���2���wT&{�bB;K���y/��^h��"�7LB� ��l���
�~�~#@j:{�u��W0��+��m�9����zfֶ:�!�ݤ<���B4�vs��zWr+�Paz[(�$���Vcm뛴�3Q }�d�5��^#lӂ����@�k	}9�&"��ֶ�Oͺx���Δ�d���"�����o�A�i����]ga����} �"U�$��m5�tZ����E�/o���T�\�i]�Y��3�yT'Q0��񃳢��&�.���Hh
2{�Yv(�u��|D����� ���Ÿ.bĉG�3շ�(�Y�Je�2�oh��v�Ԋu|�����ǁo�ށ�ʢI��m2.Q?����T\���lA)T�ۏ5Sn�c�nG =I�GZ����W2�?��������*/?�v���=�����N"�7}A|���ܜ�j�'ғ�3fY���L1����b&�N�����Q������� � ^R��Cǋ��|��a�NR7Z~���4��=�d,�w��K�T�N����

}{�ݟRb��Ӿ�8<�K��>�zF=�G�|��^� �!V/S��Gf-�J������\4gs��Z06>�w�}e�п�z\=�����gxT����39�n���ı�b'��1ClN�+�Oޯ��XH���(�O����^����l�١# ��/�&}X�v�é��%��!DV���o��3�&9Y���9O��Vb�b�`�ٸ=�[�j3�S��,��\�)���8!Ŗ�]*7N��vV�C%�D��x�ʦO��J]��z���Bv�t!^���2�#�g��&�T�a������S76�4� =[ݺ�r���y�Fy:�*Ae�wY�Q�����p(k'&�Q�<����ND`ถPuH3_�	dC�Q���#�4
��p9��8a��ŅD��z%�{rTl����2R��#����A��n��"?3K�?�ŋ�p�$���j���9i���M�-)���+��:�f�B*K�1U%(_����Whp��JY��RU�Ȑ
5�"��n���0y+�+�J9�N��B�P:���*_&K6Z��J���+��Eڃ���r,i�gC��?�LKq����;�t�N$��c�2V�S$le�����J�w	Ol���!O!�� ���b�G
�A�ݜ� �c'&�jF���a��� q���G`}<I�vC�c
������i��CF\I���|�쬿�u�g��#�vQ�/WS�pj�0�c��ԉ=FB��{���^�f.,
�(]/<���x8L���.����U��m|x��>ȗV�p�t�����A3�N[�%{���b`����{R�&���b{H�'a�����Ľq���-����=	»���}��V��|�P-���:k��nAr��V�(��Ы�R+L4�%ep�$S0��Cy�^���M�>���1�4�.ͺrP�:�l��C(o�&զ��pF��gS "�o{.�;m��\����f�z]]�\=˜F�m�qyqÀ�h��I�*g�@��j̢nr�?�פ4_&��?�t����I���y[C�s�@���R��ѷS���6�zMB
���	Ɩ8��v^��d���	�W���:�B��@:"����\��QΆ!���3��9>t�	+IU���1p�;�jkxt�_������� ��O=��4���g��~X�������i-�8�lj*>J�>�'ۘ~b���v��wh�X:����^�;��S�����#F�C*���3�3d>�7���{�&��5���w��Zlo�Y�Vt�7,�9��V<�[�L��6��MGz���jL�,/ԋƉ7���e��2��m��-��s֙/~��{r�X�����ߒ�<�ؤ�ĉMMi��ҽP�Y�Ⱳ\0&��>N uY��b	N��e	*�@Q�˿�m茯��O>H��J��'��h����T�t����
���(iy*޵�;��3ƹ2�,�����y�!p�ʡ�Jf��~���X��a�&��wb��g�ocb1����(h�m�ˊ6�����}Ǚ�ɊjS=����ȧCU�v���'{��_䃲���^���rE���i�A@#*(�@�Ac�M�xDঋi�kk�HP@Oc�����k}�oފy��?��f�r	��n���;�z�;7=^�q�Oo�H,�f^ڝ��G�����4�������w�y�F&3Di\^v�y�E:��q�g.��Sw*�l'��6t���l�{�Ը�N[=مly�=jQ��F�ޖS�2�Z8��ː�b�,y����?G>�g��'f8�5fT�cCݕLA���2qn�jA���)�b���X� ��9[װ�l�];�E1ɼm�ß�ب�w��(:?�x߅"͕|��)�Y۠������rdw�S� ��&��E����5N��\����~[�e+5Y?D����.0(�d�̍^����|�8G͓�?�PI/��~�ױ\ �K��'ͣ<0��!���/�~�{��3˜��!^����c�ƌ�9�<W�0�T:8iѸa��>p�@�r�ᖈ�PI	��[��R���,2���lMbf�i�����$ʂ���ȶ+"�yo�����s�X>�#D ��{�|�z<��v��Ap�E��y?��
����֕�cϢQ�]��h�
r�����lY�`.�i��[G�?�I8��S�c(8r�ۘ��2n{��uO�A�i����� �/?���� l�t���g��K��Ũ����g�%��j�:�%+6�}� ��6��`)/�-q�Ht��0�@dL�Nc�Hr*: �Q^�d�Oo��s ���:.WJ��:&�	�x�%=_��Ȕ*3��ۿ}���}��[��T9�J#1��g��t�i/��<�]����4n�ȠBS�I��tʂ���[|?����k,[#���>�(S�Q1�:8 ���!;�.1�},!0kɱu��b�R�ש��H��d�Me)�CQ+0�y2o����0�*�~72^�n�R�|'i;ݬ��l��z���4E��e{d��uD��M�i���)����t�+�yr�g&��P�w���Һc_���9�M�OG- ���V�T,m#��e�]�4����V�&Ϛ�}UXPhr�ĸ�-\�>ji����<��^�����Ձ�',�F>1RUN-�H�Is��D��Y��G校�Cs�d�7`K���N<T���K����Qr�!0 �0����o*�:`h^=��"�7�]_�����V�+S�M���\��l�ɠ�ɯ��6�����dk����� m��4ی$;"��5�;IBxIx�rX3=�r�������P��Y�Gܬ|LzjTѿ`n;IYv<d����"BXk��+� �ә�-��H������c�8ǒ�rn��'��Ņ�����%q��c�n0�B7�-o�"�}ё�4#�oP���d��kߦm��|N�(���H��4� ����(~&����H�A��%O�^Q?��4��A�h�ŏ�%n�1�c�XȺ7�	X0F�ohz.��(��g��R��wҴ�}y�	�̮�'�N}<3z&�����&���J�T�(nJ�!���c��\�LЮ�ePrQ�=g�v��y��HШ�q���f�2gw�۲W
�b�]jR��@�&� }[ P.:w��8�W-s�1Cٟ=?������`�Sд�f���H�3�j�V!.�6��Yr��MnӼ��|�*:��8����{oq��U���B�ڥ���k�֒����,�8
 �F9X_O	BN��\��⭧@�hda�6��+z�EB�䭗k���e�
�#�6�u�.c�V`{D���C�hE�3~I9��GggD�L��5���6���iA��<v��!a��l(����i��$��MźMgS{�����B�����}��| ����Y,ݭ�&� �q��N�H�ӹ��t��j��!M�5�]@��9]A��7�lIAB@��K��_y�Ժ~-\�%��S������h�l�g��-Ć��F��������Mf�2(_ ϓ;㝔�t>�@��!N���5�ۑ�Y�p�(��j�Y�S+���9a?�/��9�L�U���jkX� ��.l��ݯ��>E�5�fX��7���T�������|^��0��Tz(X$���@�MA�����xBw�j��xe�&�����b�Űj(��M�O�/�'R�����'�ڒ,#�.*�|�M`�]�}���=�\X	��ljGM��׋��*���k���D�Q!�Y=�ÌW����ڷ�i���	��ĝ!��B�4V	��j��r��_��J��`��lN��"���zjS �ߕ��M���� ]��,�'��&�˩����i��T>K__80�G<��+>���>N�^$���%���7��X퟿����w�I1�8'Β�I�E�>9���繘��0�����3�^�*��a��Σ�"�h��_��nf�w�AYic1B{7��Ϗ��0�p�6���>�k�^-�b�\;d?���a^5FRd+���H&�=���1
X�~��I`P�^��z�~�J�i����">�}Q�RH6����=R���Up竼��0���{�����E��m�<�N��E����$��p�s�����˄����id/�g�~
�&�=�s %�Ʊ�Q�B�p��!����k�k���7�-���v�a,4rZ4�a�(������M��O��=�.Ώ�c#�Ds��mߵǽ��K��%x��]���G�K� ��6~�@��ˣ�W�����-�y�&���sL(�G��4�ʕy ��#��k�%��\ �dX�l�઀�U"�:uB�����Ɗ�/�{�7�$=�ᘫ�K�����I[J���3=a���3){P�4�D0�C�|��@�:�R�!6���ۭb���������=��^K	�u:�$�I�
W)�U��J13B,/MA�`��*ll�rv�W/Y��i7�z*��E磍lrhc?01��<����	�ˎ`���E^0�+��N/j�:Eg�7π�����IRWt��cӰ����>$��^���~`�;C� ����,����u�Li2�󮒉�����Uk_p�%pJo�l���ь���O��[sq$�Fb3�/���AM��P�j��6M�ŏ��~,��)Ez�5�RE��!��l�ϙ�`�H�\$�0�ՠ@ �?��ܞJ�1�ߩ#��Qj�a�m���-���F�q��/� ��@Fg������sxIaPV�c���E��.��;w�8��v$�T:���r�X�t�@�|����厕�ei ��0���U��k�M�qD�o�s�;6�����Նa��2�Y)܉����� 4�SwHBB*q�K	⏩��4�-gd������W dj��	�N�>;�k��ʜ�g�}�0������wNٜ��.Ⲇz��v�~��Q�E�5���?�մ�vdUĀ+�{��k�?��ȡ>Q� #3FN(�n��=�������pB�I��S~�����>̒��2����;�9��z�}��qT�H9�GW/s���F�!���9���#�D�^l53��j3x�Jm�!U�dqݺ��yۄ�vp� 1QBn�5�;�.��؀��u\��埁�ͧ�j *�F�N;Ec�=��y�^<����
3��l�3t/5�����P�賁�J��@)�m�l������j𺽋��3�,w��c%�$���0���L�R�a�2-~�eVm �D.aV�Tȝ�#wCW�e���P�A��eS�l�?=R꽟+_t�P�)U���_�{!�lvh��IGb���;�h'ݧ�ͯĄogN.�ǽ�X���}��GG>Y�^�6<�\	�f��&�e"1���"����S3��J�u٤�^��YNʵ�W�ԍ�+�9��5���MB����R�.n�f-�Ua͖�<Ĺ��s�up��#���9�i�ۍ}��$.�3 �:̎YıH�ȶ\�e@%�������ն��\�AMg��6F�b�(��g=��h;�>a�'�P�]�}oh(�C�_�7�+��b�H�$��G�r,��E��l����TCfޥG�.Y_�⃒� O�Bz��~.����k�٠{K$ֱ��lR�*�}�g�����NL��C̅q��J��פ)t�Z��,�{��!�z���Q�,7~zM����1*GE{P	�(���\��2�o��VH%��wp� �~�{�eK�]�FM�FG��m��y�(N�<Ԅ��ַ�C2�D2­�ʧ�x0�&ZL���z��Lx��;15�-��B��T����7ߧ>�r�/pz
���1嵲x�_�.i����	 <vF�%��=����v����L=�l��g$��e����5t3�C�>����'�RAwpTC�ex�ۭ���D�]�S����u��Gc�Ԗ$�"��C���:ki�����Ӣz�iB�x�#��Tb�g�[�o� K/�X��>L��y�&{��u���R˺�
�������`5�tߊ�%�I*^��:(���$�\�Q�&�����-�zj�hr�NK/�1�e+�������&M�V/'O&�p,b�uֵN� ��i�¼R��ĥs�;��H�:QM��A0CiiR������iG��2"���j9��.�w�z��xy�]�sGKSG3�.�%���~�q�wG����]��iƯ�;��Q\H�E�R���f�@?���z���ES�&i��t�|�.���0%�w��9��QYK��^�/�^����Sl��B� �J\xِ��H8: ��p�����^ן\���gcaj�B�\�k�� �5��Wf�Z�-�!y���[e̝5U�U�k�������@��jܨ�)-�M	b�mǭ�a��.;<'>��n�}+�h�yft��Q�M��ؔʂ������W�؄�B�$
�F�;�zc�0J��Q&�'1$��ʝ�g�0/!���>��:vSm�t��V�(Sj,Ѝ�=G�����@Oi���,1�o?B�'<��8M`�jj�/q�7_����
�ń�|Ԅ��w������B�S�J��"D�DJ�`��Ù���Uא{��=�|��H>""*�n�YV�*�j$���cB�S�(��K���o��jIAֽ0X�ic[5<�`ĘG�!m�t|����q��0�Gd��ePN���fZt3��12j���%�?!��]����ՋR��BYZ4��g(3O�#���E����Y;� w�!
�r��=w�`}�O�=E�$uec�ſ`�8>MT�����%v�,�e����h0=� �C^���U�?2Y$��L�-K����7a��uu����@%�*�����8�]���"1`Y(��gW������w�R�M��ǒ�Xh�iﲎe-K�*�u_�pf[��_2��[Q�L��~��q���l/w�b��c���\��r��&�P��P��h�!�vTM�g#��s7�v�'vˠ�ݖ.�L�us]�Ql�?k��n�B��ra�B��_VB��9��{�g�	�oMš_��p�q[p5�� 6�}�R_��wq̿�|2��Q5�������p��U�Q��3��B!z"3� �t��}�}����px�#�B���{�XI�h�cK�
���7�B���x�;�p�Nm!����V�Eqy>0�������$�u`f�ߚ4�m���]����*�����Ty�*�h���C�T�������R�e VP��=$����0�/8�X����4�IW#^����c!�����qF/�A;�PRɚak��>�G)"�"+A��S2��^5
�{��=vfg�~�mr����)d����	}]�n0�ϡ����B;�a�{��9)#t�H��B��[�sn�)���q�.áY�5\�ed�h��m�j�����Xm�"xל⠸p����e�H�Q��OD�<��U����.�ڢT�;0�����-���H�]�"�!�	��O������4;Y�k�V�Rm�����Fs跘�XU9�������m,D�dn4D]��N3č~]w>���C��	1L��Կu�zv�x�m}o�o�\"�����ׄ��,M�8 �>�2����_Y��F"�~ �C���FH�xB֕�֍�'A�DC�o�~�/�����`^@̯d�3��Q�`_Ud�d#@SO�'!~�w:B�\QQ60V��eqJ7��A�}TFB�VUEI7*��6�In&�*�jiԼ��2@��ȳѹڣ^wƎ,1���%,u^�,A�ڳ2����'\IPZ�Q�V�0Cː�5L����Z��5�쏯
��5���=�ՈX��*��ar����￼�P�E�#75�Z��}�ȹȶ�a�#o򀅧��II��� �5�����J<���`0�U�8.r����}��mjgt�EeM��z��5�!�r�9(��w��A�Q	�N�+8�n յ�9��&=��L>%���ɸ�$����sg���?|�CR��G���Z���isn����	����N�^,"Ć ���7�/bu]Fi~KZ��F
���l��Ƽ4
����/�@�3PkM#��|4�֭�y�L�g�~K�\��H�-��f:ߵ�隆4���)Hʀ����/u�p,!9��W��.� �����Y��Y`n���5GqׁO�#_N�Gg�xڲk���@�O'銌�>�1�v�T�F7L�=�!�>	[�L�IG�'%9�-�18<V0�M���|z)ӟˑ �6�$�� �Ҝa�4���^�75�Ǥz.���
�y߰�����7շ�U�2�ٖ:�4�z����]( �2F4
"( ��a�� ��^z>�*���$�z ͫ���vZ�a����I��o�q�4�����f�#�Z�t�Ӈ�^vW6��7����5�eo �_���9�TB"`�\�h2�v�h�מs5�=�N��k�G���L&����`���G��8A�������!Xo�����t�UО��<��I�E��M�" ���I>�Q�,�P���t �ky��ב����Z^�Rc%=yʎ�VO	{��}�Ƒ�������dm�{tE�^A-��d4��d�g:�������y�ҹd���^zKP�T�i��e��)�v
N�����Q�0wGyj��v���wl�'��]�R��x�S$�]^zi=H���ʠ��*�y�0�_I�?"���4��e�4���B��~��簣9򆸩c��'HF̠���#�Q�bP���ԃ�d��QdGn�CrUw}=ú�w*Kv���H��frD^u$}�#&E�$,��ur���!�N����z�~l��ʤ��$�`���� vG�"���7:V�PKj'!axwr5��zw�FP3a�]W�%�^�%c�s�4�P�n*�;I]}	��?e��*���έl,/,��DB�����얕���yl�oo��i�H�$ħz��(b�=�$Mc�h��<w:�[�w���'��]����_���;�1T�\����;T�b�D'���kTIZ�ؚ
ܿ�Q�<�wW�_�ޚhS��!K���"Y�_瓑<:����H�� d�O͝-W��[�W�)��غ��E� �	*m�L��Y���+�*���Ie�0�q�]�>>^��-EV+H���z�ϵ�F��SKG�ea5�
ϧ�iQ �(6e�NAE��5R{��������˄@��ٵ��<��;�ڐ-y���0�eqJ���)�%�����#�sLB�ۖk��Nn�(���%Gr��j
Zh�}�:��2���3!�@Z�Tg�^=��A����ƻA9U@�7�[�=��
O�����[�F�|���%�"�J+x�3�4BL���MJW��:Ќo_��-���X����3 |5h�u�fn��*���@�%(� Xy9@[,��@6�do1 `4��;_[�6��f-�u�����N��f�H��; xվ4�b2��鮪|��FS����7���֤���ʱ,o��ݯ���׷F=�;"���P���c%�V���,%��]p5H���dTB�κD)��!'�mi,o�G�'��}b�uz��zf{��g�X�ǀ�� d����.� ��<Û�~�IN��Z�؆�FD:�h��0�Ȝ�"]kHOէ@3��Lq^����^���,	(��5��ZB4�5ƅ���(�9
e���.t{C��_�2Q"��E�d�b�T�Y_���^��щa�
��<�m������$=G_�����I��L��\_�M<���m�&�;��ؼ�zu7�kR\��A���usj���D<�vM�l�b��be���4-�����=dʉR���W���U9��}Ht�t[(���g���3I�WMFH������Lo	a�1��I��!ݺ��ŅzJf��x+H��%&����2b��P���wK;�k��OI
,���\���6V�N�0�t��h>�����H�����,Bj��bUDa6�k�%U�P�.�,�^�R	��<	���P��R�5vخYV�k��Άr�5&��I�kk���S�|�5�>{���a���r�z�P�s�V;�����ٲ)����r�w��֪���7��'H��
P���0Ex�e"�����j^`q˅A���e�jB���&	�4/���E\�aMRP
hl�Z2u;e[r��b��Z������u���/���Z��쀇�hQ!�,����<oi�/,��c_$IE��B�\�vȬ)t�B��V����º-/4�ѥ���x]�u?ꃪ�^D@w1rM~t��J�ɽ�'IR��"��Ċ]'��AuުN����X8U��Z�TW�.F��}�������R�	h�.�6B4Le(C�؁*��&̅�/j^o��$	�u
.�*�4��M�g�v���-O<�\�L�F�<\��L��A�>��t�Kv$�����&��Ʒ�8�ųDm?�l�<��K������M/RHbub�����zr�Zo'cx?#��Di�	�y{�=�_�yo�7K�+�z6
_�_�
��M�I�2���\\3o��{���6�����u��aCv|ȡ���|-�U��9�@���5y��FB�� �&J�M%�K �筯���WI���(,�yrDJ��h{�H�rTZ��:�gU}���������)Ó�b=)��_x�ڶ���?[�"I悇A�Vn�ۧcA�������e7�7�0��}�Ֆt��t� �86<��;��Ol�b�'y�)�CT�>����u�P���|x��qB-�D�?��N���W��<>�	��A���$w�M!�q;#0-;�#���A�u[��B^�d�bx�\XGd#����c�w=y����D˽r��<:/qq���J,
�ǝ���P'y@[�f�r@&������N�~��i2�PJՋ{�6��*��u�f*'k:���kȕe�|#�`�U�A���G�޿��K�WjP�X���ְM�`}����j9�қ]�(��;�L�1h�MP���̀���{�K�{��w��x0�G��F��"�
K.�Ib7��L���M~K�"���ɉ�YfHU�_~h�	!��AFI�d��a��9-[Z�0�mA��]�υ$q�����n���N��T���:��s�sq�Ӫ�|�v�-K��Il�%�ǐt�A��tJ{�=i���[�L�Z�E�ڄ��Dް*_��Yc�sتBNY���<b��)��k��o���`���"�d��|<�<��? t7�U--{���냚�C��c�@^���EP���Px�ɵ�)����yu�n9�o�9��"�<�㣫lm+�����:zq��%)�s����J�2�g��a:]���12�&�Y�)5�@[�qsm������؇�`is��X�{���@�M���6���F$��쥔\���Vg��3v1���7����]H8�@��\��c`���û �f�����Ӧ'`�01�s�7�0?�C�#d��{�6o��7%���>	��vJ�G����XRJg��Q.O�-�?����L{�s�A/C24Hr�*��H�Z�$�TS�������&�Ɋ��C�	�	T�b�{WJ-F}�D��G�^��h����2�~��c�}dEe�d��
�&��0�hw�s����E{�����%7���0���u��&O���X���e�Ha��L�bp`ٴ�3���� �d��+%}����šo�ؑ�J�)o�Q��P������p�(�3(E�]��y�����)��]~f9<W&?��Ɠ�4U�c[h�=荏m�=�hqv"�)د�E�eF�}��jB+�����/mնZ�nj���\�)`�*�K� c��^���¬�b�q�˩�A�}@7�2V�Z��a�?���$-��	��6M0��>M��6ʁ_���;�M_W�I�T���Ih�\������=�8�x��9d''g �z�|��"1[���D	�WfUx�m�h�~��k��F����1�5�seX�!�n�]j����q��e��6�������ss��LՃ������G@;>���l�t���-&�p��M������Ց���`�Nϟ��0?����q�X�}����'ŵj,e�"�}d.��_���	�����\��~�A�<߯�i�eU�m�����gI�}��y^y�tEd��f{��,��<PY]^h8�RE�ڃ���S�o��+���bd'4b����4~=�4��ǳ�ė���!�y��diB�*|(?���0�I^���^r��o����p��Z�d�\}Т�5-���y��^����ox�W�Қ�y&V��hHٛP�ZǖV��&WS���������u�
3�ҋ>m�ܴ]�/z�R$rU)m	V'}�����|��1��]�`""VvDYq�k0:zV�;��u��p �~3N<!4ӷN�/p� \�#Q픩��8����E���~ز٢M�!�O��o�k��%�X:�2�2���������]��\L��l����\�lLM��H��oV<T���(���,e��<��(�o�D� �E6�{����l��7�׃�5f�@kf\ ���E���5��(���#4�f1%%�����Dܱ������֝=�]e����,hg'�K:�{)�t&��V�~$����.�cE�yP���"�Qv(���֏r7TF �`�K����"�D�D��Y�uO�P�E�J�M����k����W��2����_.ryFPkb�u��-K�!���*��63=���C�̓/�fp�T����IC]5��Q�l���C1��?>9nf�K�Sp2�(.g�G�`�2Ԭ��W6,\��7����T��_zG��Eo�z�-{
��VM��f��Tz࿇*ȮAM��w�m`+���<���r�ZՖ5߰,����
f_��P]��iI��CE�-?=�&=����r#�_��W4M� ��|v�f t0zkgR�"�d��!$�}����7'9��@��W)M7:h�x� =��䭬��ཅ�t�)f��D�te��q�Н�P�K�Q�]Y�_9ћ��,�&:Tx۸?}�R������It���"ʽh}�Q���l�����9��`i�Aڕ#dd$S(~����AV���4 �Ϭ��5a^���xq
޳Z2��J����֮���o Uq�]w�Z�V]��<���~�?�gf��mFE�)h�h��n�v�a��,�*�i0k��V�fm� �r8�M����6b�Ťgo�U�-�e�2q��`��r�H�����tl�ˆ�daP��q�	e�;�TtT�~]�%l�)l䅇B7��h���Zo�ɢ �zAǕҁ��y]A�Bꬂj�#.]t�oX�9�����#�v�I��O}�;�hoM�U�:��'�W��Pe����I3ԣ�؁�'�ξ�}y�k��k���x��z����3���c���coed��6w��1 ���[cG���d�H2kx�"y�
AOf� 6����Q�*����x�{c|�c���U���|w	W��ok"���H��ҡI*�v�/r�0��P� @�T ��JVmp���3N �i�F���k��&�;�)��j�]����5���j܋���7�� /5@���]љ!�s�5��T!�=R
pjp-wLLv5�{����)�LD �
��aD=D}���2���z��xR��
]�M�B��t`�^`�b��dG�����h��].�=�oz.�D�ȘoqZ6v��i�Y�����r\*�N)A���UI��W+�y}�ɴ8+ɱ���$K)�}s��������43��$�s�`�ܦ�!�3b�:����4[V8s�~3Q��Ύ �Y����h8���m��!�>��u[ˎr�p�1������S	d���Ol!ydR�q�67�&o��!R:���3j�;� V�;�̚K�3�jR4�����*�
����{�/P�b���ꖗ�d�gt���^YW�mː׺�kcα��	<��KG���9���܃�@5�ק@��Vv�4B_��� ��kV<F�>�����9����i�4���Zb�2�b��9��v|�V~-�f�s񇊯���xu�d#�uZ�A�\��[6��@R�F��n者�BlC�z.�aN���R��5�R�<30���Cw��֍��.����a�ȝq���h7����vL ����v�Eh�P���u��@��4#�h���1']��W���9��O��Ѷ}j�5պ<1�*Q���%�26�߇��)d�6��ى;�0���u�.jۉ���c��5$]a����%9�c6o���;݀�P�F�m�����h3��ۚ&jq,d$+��TBo�)}}���(LQ�,�Cs>���m�d��eD�:��V�-{�D�\+a��ɜ5�����#�hp͕H�ȷ)�������r߳�w8�\��D�(�n08}ΙF������-�{��?R��io�`�퇋;��
"l#;�Z���
����&�v�zH*:����@�[B넑��w�q:ri�(3Rr�EhK�c�r�j�N83��L��7x��$>�I���$����|[yh��|����V/��m�~���A�{� ����g�Hw�.��x�T\�s�C��j���$n�<�ݦ7�"�39���1�d��z9��8�l#c�{��0"#l4��8��L3�������JI1d�yb ���8�y.�B�G����L�sZB�kU
~}�9��M�)h�)4H����/�P�R)����TU�AO�x�p޼�Y7©78���\�{�*�<�DĀe�;*�o��1Nw
�VL�{�����׭�>�ə��Uk5�k����Cd2EC�Pd!Ä]�
��JZ�6�D���L��4�A������3:���N�-yI� ��g�6�"�/�6������i�")=��1�p��S;��0�����b�Ujiw�Ξ��<�Rd���q��q¯��s�#.y�d<�c���2���W��<y�Y~�l��N,q��S��Fzf-�/I�#�/P�N��0U���ƹ����[~�+�V�U��D7�FǞ��]:�Pǰ��`l0P?/�����|�l'��P-pꍟ��9��oƉ)�NgM����K�
K��*o��$C��W;ٷy椩u�_���pXd8�4OyUr����P�M oa3R���'	�Ů� ~xŮ 5�h�X�Crf4��e�-�Lh�75Y>=e���*�]�붕�����d��G�1��ƅ� ����}�ͺ)�!o�/��%U���g�����e ��{���b��!�i��N6����Ҁ�%��ks[nS�)���0A�d(�x��:�W�iNx�*(�OrDn��uL��Az%^�r���J�qĉ�8"��S#���צP@���x��O�z��,)�d���K�n'پ�W�fo��"�Ft���\`������3��o�"��\2�F� !L�#Yq=�sv[�&�^�e�v�"d�>U�Dm�N�W3k�7�
U�1=�_�o�,���!uS\�k|���)�t6ð�´5p��8j�R���ϙ�Bk9����Q��
1a�T���+���4�c�'�E�u��R�6�i�+�u�%՗b�ư�#4t���A���	m��Փ����0ޞ߭(-�tf�U��@��ؗ�f���7,�����}:ju	h���1�ըO��1�7(1e�\�MG��&����?�`�!�TW(����0��c14� 4�Å#n�f0*��7�b]l��E]e���P0ٯ��?����rxˇ�Z�SW��չ���v-��璱�x�N���B��-�S�"�c����* �'? ��ֺ���rhF;]�#�q���7�� ^�r��q�W�:q+���㼨�;HH��}��D��x����:#�G|�����	�b��� L�^C�`���wpS *��Z��Z��:���xf��~+�ސ Kϥ���\�mмa���~� B<_��H BP?�S
��K?4�+ې%D��Pj���y�?��5���7���oN[2[>gy8zZt�Q}����/g�j�f��k�w���e�Li8dMv]�=�I8�3��-P	��;����1�)8� ۄ�A�]��IݍUK�����0���J�U֗��>9����2p�\�B�n˥�a� d� ���P�ڔr��6&벝�=����'��wuV�C��?��-��Zx��[��[`��o�0�3��{��.Hi��A��|m�ȍ�!+yAd��`4.)�H�(}�k�J6?>P�J%T(Hp5�1pq�M��e�ǣߚJv�4Y��ɉ��F	2ߖ<:9��l���+���(cˉ�H�~L���<��g�#�v�:-J#zE�Td����Ԧ���@b����G�JAb&�͎�e�7�Lhv��Ƈ�X'xY�X�֦�rv���b9��0"m��O��!l���<�Ŏ�7-[j���Ũ�0�3�\��V[?�t@�\���V�;b\����u7����BcK�r&�X���s�ꅄhu��J�j�,��)=�n�k;ca�V���fOU����O�bs��ghæ+D���2BWߓ�C#GT�Ÿ5�E.Z�����()��@
��u�凵��~�=k���٬��PO��\Fن׭�%1�ud��h
���B��种p8eM�MEM0��T���u��=�D	[�żF�,��:���r�w��n��>٬���Y�G�~�x�G��F�}�V1�=�:�_����_��R�TdD5����0<U[.+�U��� o�tv��V��.����BX *H����Ls�>��K�]��_�=׀�@f��ebǹ6�8�k��n�QU�0G:>�a�c����.��	�y�ʯ�&�W(ti����]�T�d��*ˠ:3fb��߇�Kn�o(��v	�<��y9�83<P�b�2��#=h�$�Fl��7�~�|�m�� ��c�����f��e���� ��bt/� zHO5���r+�f�v�^��b��w/����3n����e;)��.,�R���ua[�8�	����Ss�+�=��������lZ�k,�E]�α�Q�(ۀf���Rbwh~�S����k����]����@�MP��k0^B>?��у��S������d�Mp�+nR���F+_��*�(���� ���C_�N�  ��y��]��u��I�����+S�4�+��B���	���Z��O�ZC�i���x_���q��y�Ʌ�`cw�s�0Ƴ�_H4�|������K]�px_/1���B-n�T�ʏ�૨�s��h�,�S=4r�-�d����+Jk:))\����l�!��u�V����Wt����t=2 g�O�:4��%�RRU�<�YΖ17	��Z~�CHv�3�~��=���V�R�lʬ�y�-te�r�o�aM��R���h�]l�(�|����_��7�h��
LiG}� �E����POo6�rj��E�����v�&�7�.��~ήx�� ji��q+�f� BH_��.��ű*j��O\+�V�Lf�ЋKz~$3[-d5;��)�2��*��Vm6���ّ!.{�y	��Mћ՛�d,�����ߢ΃P�oә/}Q��]El���OB��v4�U�v�����L��R{�+e�9s*�͐��HW�fG��)7�%YC�P�R��$L�T��,��Y��cN��S�d��Z�Ā,��,�aa����e�&�(���6B��Y����-֓�y12lT�mQ��*7b���4��S����������sz�|<
#3����)�u�tA��ñ�Kl�m�1�A������ `�@��zr nj������g�3J���7YƎ��8N��+�#[	iq��0���@�/���33n��u��t���s��sw�wR��8 ���2�dO֛H99Z.���]��>Ɠ�LU�l\���C��[��Pd�]��H-�a�/>B�m!5#�P�xe���s'���<X���y��BV������*�I����s;rMj�gw�W��~�}�J�Y�C�Xw�knX34�W�e�̴��t}��/w�+������,�6�������a~�,ކ��P,J�y{bx�.u�t���8L�u|D4K��Ǟ���K�n�$��L=�,�5��J�� i���o3��%]�"�V�ر�sk0}z�F2I����D�G���!�A4�j�wҕs;Q�H	��!����7م�Hr���a���F�CuJ`c��.�?�b�O႓�{%wK�^b��$&���z�>�*&ku����W(H��ڦi�^��%�h�}J��A���':۩a����ݥ��o������9���8��r� �r�,ik��)9� ;�8��p��5�f�S��8�>�&K%�',Ce磸�{�<�E�:?�_V��x����)�|�A��<AG�f5��1�м��,`��w�f�$�1s��q�)�@IKn�?��:���!�����I|�?LR
��� m��zS��PsA�ƫ���j2hZ}��58��������t�~�]b�tI������:^P��)��f��C�,�dN?���M(lVv�f�eݜ�ƞ�E�w���<'ߟ���&�S�l�{w�O�o\*	��x�	����|_km5����h�[&lځ��z"E�El�q�(���Lr�
�0`A����h}�|�K�OឨFNJ�����dO�f�D�;���Ѽ �.Xk��WW���0>�zd�T��T����2�z5llϳ��SlP��m����c^[���>
��._���T3���K5��Ky���ҁ�>�`X���vH|Z!�)��i?���P���t���)[���^����m�P��O���&���̤zmc�;s�������bp�:��MS�66��#����P��ӆm�.	�Hlсt���~dbڇĖ2��j�x:�^��+?�<�aG�)	tpg����S����i����p�/:Y�ʞ�Ӣ"o��~T��c�mG
� WC��W����@�ګ�X�h��1�I�w��l��~%����r�Pő�V��4��V2���E�F�XV?���_�%F�Q����%g��_���H���w���D~��oV�_���p�a�r|'!���:�>U�d��tD��y�*�����1�wr�M����3�o��D})տaPS)�#C���  ��RQI�ߐ^C|B"�8Y�A�$΃)F	���z|�g!��EI��ϪG���12]�B�U�aTT+R��},z��8~�^��4�G�k��<�`^~0�ӕ+���l�|�<艜��Q-�T΄�}!��dR;�o�� 
/�w8Z�1��L��Wz����n�~!�g>�Fr'�l����X�*�M����+������΁�{�3;�5g�Jt&oVP�x�+�H�gƔ�,Hl>���I�b���3t7��>�#�ts��g&�Y��O�'a�Н��;g���+ŋP���J'Z�:��A���[���7������ :�֖T�:��S��s��<s����5��M��h���vԾ�+q�ME���CL�-�t@�#�}\�ϋ�e෹܅Xwck�~vGH�"H%���4U^�,�b4T��P���o�,��j-hS�Ҩ�lDW�7�ѠS��˪�)k��2{f����'�]�~�s˴�G=�	e�Q%�\*�� �uKܒ�(�����-��
�pI@9"}��v�#�-ޞ,
�
�#�-�ũ�4��D�����s��I��p��/�d���������«5��c�w��}�z[�DI��@�<�G�O|Y-E\�I�GN����t��$R����bU�R�hܢd≇��(<5U2A��f��¿D�kq5X�vF�t0�B���!�0=Ͽ���H�
Y�w�	C�擉�,�Fx^���"��"�Y-"���
D�Al���B�4��D!�v�?���\�/M:� O'Y&����
�� �a^������!ʖ��U0�r��!�y�@�Bþ{�}�ڊ�?f�]��g�t+1H�K����%�Iź[J�(^�L#��A�=�|��8+�K���"��N\F�u�z���6m����(�`�Y�Pm�}�6j�%�`�m��tL��n���?���jc!�j�)�ӪUo�S��L�pO�2�s��ˋU�4Zt�L;�J֫�6��������n�E"5M�g�}��R�?,�ogk6"!�D��[@���!:�,K�a\'%�fNe}��R|;T�c�@Df�4���]�ɯ6���ҝ/~#�{�#�r�l��}�n��=j�ƃVS��|'�b�ob#�L^�V衟��{�|���.[����Moc���7�U�8���PK�l���̈́.��d��~P&r+3z�����8��m��N���A�f�-oI��^2�hi3�������:#�4m�|4V\�X3��X�`u��x�f�O��|�GB�ڝܓI�3���m(Vm�}{� ]9>�ʩ�$sv���YG�ŊX��R�4w�'Zr�!�����׺�#��xH�h���3�o����*��l̳C�O��vj���<dL�`�������{�+�����.f���1}R;�%�Ln�(�c'	���(�|�5��їs�V�3>a�z�)>��/�"������lRX��)`[��zr��(��T4�W�M��|."w9"=[4m���B�1\̞��S@Z����F����4��7��p�+�?>~	�7ؚ!���k����ү�Z�O �)����f�	��E���.&���ě�7�6�r:�Ϗ��dߒ�~C^���	��B�q&��'/�u���(�'0���YۗrOUO���E[�r�U
׹��o��E�����P����<r����`,�c����$~�B/n�(���q�[I�V����T�Hjf�U��y�,�|��E��2�ťȀ1��;��H!���xt/Kd͟v�+�_����U&��єԧ+�$!-puf���τ;�P[��orB�����$�_3�C�����0+}�<z�QD����7�I���"j����cE�z��/@�[�$�>-�L.�<�	�I���}�%�R�
��a�zI՗t�Y��G��Ķ��wJ�YBe�<�z���~��K��k��7�}i�lSw�
O���4E�/RMJ����3���,]����N�o[�aҝ�� #��x��4������T��~�7�j���[un�~�mM�VM���G0��I�Y��h�9.s\몸���-Á���G(@Lx^�:��r��6�����mm�{w���"D��7���6�=��))i|=�ϋ�9P�2�Xѣ(�
̎�a�n!A��T�g"2��V\U"8���ɣ�x���]�����4AFu��F65�H��L��~�8M����0���R�n�Y�/��@27�p�ғ7�/1���h#�Q�П}��<��%���g2']{s�	���xH�����m�@Z_�QGp)�6����i��%	d�u��!�>5˟#^Ί��
J�]��!D�6<�6�Af�N��:�i?�K?�Mvj��2?/�M%g�܌�&ݬx�p�7F���S���M�/e����AK���V	w�Y$@�@��y�K������jݲ�%^���1��4����)��~���ꄘ�G����b�>�KF�_������Nw��tE��~����~������ݮ���E7��@��� /�j�̍_��^���T��z��Q�e�8�K��Dr�z��?'�Ȩ���Ĥ\�C��R��2�ʁy0��?�X��iϑ�Κ��-���Zs���Y@��d��W�<�Ab��Q��{L�:�y�jy��GpA���+�����q���Vc�~ބ|.�y�	��s����!-�S{T��C�y�|{اm�ih��h���-��o�Az&lS������Qe�P��m�i�8�K>�3���� U��R,|���g�O$��`5��� �P��C�*m���)�*�Vy�͇9�y>������#���]���w%��T��@���%H�f5���%��wꞣ5��MZ��ǒ�a��f�m�Ϗ���#N��Х&OY&ң�@���� ]���R���1�d��+��Gۑ8t:�o�S��^��"�6�D��,eF��
(�!F7���gu�|��[ϳ�[H��g{i(9�qI*n��Ӎ�%�ώs5� �:�y^v�0~�~]��e؆X��3B�س��)��_0�����x�����]"D��IH��ϐb%!U��/ت�K?]f���n���8N�� �������@Ϻ�]�A}� F�2dM�6��P��U����Bt`����z&f���<���U�*��l#= T��f�� E������S㷄^��}*�Srq?��}�F#��^׬�R�Z$��>���3�������C2�v����EM�����^�>8���Z����%5Kna�+Q��qڻp���P�29����4��jrr"Ch*?�Yb]�E���V>ʭυsJmQ�SO�_̟#�Wò+
�(=�����/�;���:
g�K��L����p�Э�zC��ot�W:������+b�f����M��B��9g���W�-��# �՘�pj�l��v2�^q;m�FyO5���,&ھU �	j �%�B7e8ʉ���w۔�������ɺ�>�K|d[1�0Q���y mw7��t�[Wd��Vgd�2ve�O,n�-
: pr%�q������C��~�h�߿���Չ�jj��<�KOſ��1
-��H��F:�P�? �����M�c)�������LE�iߐxBm� )����MD$a�셕�7���зo�٧!�v��/T�#	!��!��7�X��1 �b��qa	��P��I*�-�d�4�735-O�����%"M��D�{�;�A%�&�e	�o�דT��W�9U�<�0fg�3��J�����	�ͦ���nH���϶"�#j �JGH��V��0	�AHI��*/������^�wP�c�Z.g�d/��?�/�,3�Є�[���9��W+I�ü��{[v�/2H���J��	'Z��C��c���u�v0Kb�6\ֽ���{����P�?O?%��v�t0H��HbU_�z�?��߮�#�WG@�⾄��PRz�&Wx)��cR/S�4�)`ﲆ�7j���<�M��(Y��iEiט���,�#�^�+#���:4D/��f���/UNk��d �*
� bM𽢘%j�,L�W��"`�q�g�]�`m��خϒ�^0Ёˣ@��^���Z������XtJ�JrS�{���a=��������	�����n���Ȼ�X��H���ʄZU2�LH��@ˏ�\\%��g�F��D\cF@�8�ܞp���z٤��SR9��3z(�Z�4�Ze�Z��R+�񊜦gɘ�rŨPʬG]��X���q��5ݐߓYOw���?�~����s�M6�e�#r�Q�N�ND̖o�r��+�zѐz�	,�S_
T�>���<nؚ�1�x�'��`�j>���Cnj=e�Ѣ/F,lT��W�B�,�3{2�ª��3�;���x�\��#�w����cx��1P!��>{ajj�q�>�)��<:ۭ�\T���e�?�ՒTS��0wt�����ج��َ��Z]|v��IЕ:3
�ڮ��mJÇ�v�������}���Cۻ�X{�]��E���`/%`e� ږ).%�20��4���cҾ��)�0V�TƦ!Y��f��$y��=��Hr	�:=.}��z�A��D��6���?�����c��0`k3�_�V��P��[�6�E$�'�>V�'X7����_Nu����x�� Y��b��p_3@������Cj<�'��k�"����m	̰���,
lx�*ɺ�M��9��r�|zO��B��e[-�K�
!�F�7̌/ �zL�{��/&-.�_����7�5y��� ���T�ڇ� �yE]&�a�Q�r��o7���}�gC�L�n�b<`���7<�'j��G�Xu$��^0n1m���4k��~9����,����|>�"���c�7�G�+��|M���H	���GN-Su�xjP�t�:��mv��L_ko�/�Ja"*S^6b���U��b�lcs��Y�k3�Lb$8��>]����/�!I뛌!���"���ϠثU�r�V}~�˧��@8"�#�f�o�rK�q���.l���'Jl���Z�#���-B��޹'�:U�\;�D�NAoJdd�'���/R�����Do["&A���5���(K�(�Sd.��۾)�/r���#�[��S�\���i`�|A������^�����)�?
n��u���a������.�����g����h��Usu��8j�1���ul��G�m�����
E'�q�0p�k`|�m��w�9 �C d]�b5�-���_����ץ0)g�E}�㟼��c�c�EC1�*�M�g����ի��~�N),Ro,�4:8�2�jqq�JR9��/ؐ,{B�e"��!��+�B�!nJ�o'�4�������AJ�E(��	[tFc�ŴG��*�xД��<�jˋ�C��m�wφ"��>�;g/g��E̬1�� r)�f�%Α�fm~�[����j�4Q�/�|���P@�+\-����]��
�+H��3b~�f׼�� S�����ǐt�J�*+�Jے�7W��2]����VF ��e���:�n�e2�*2����V����?&8.[(��)�~&�^�ڕf��Kx�-p����n�olZ�-F_������WU���AZ�[�����gS[�E���>��"�c)�?f6yܸ�J8�������3F��X_{3�/:{�Y@����ȼ�����5�悺[4�]�z�b����ڄW�P�'+ef9[�*ur5|�8a����k+�D�� '�J��T&K�����#�)�qR�߉�9ce���W��Nz�������u��g�_�n�l|{Nh�B��6U�%�*�L8�f����J�]��[ַ��t�)y���Ehq[�������Du�*6U%zš��S�T! �~�<�;����́|7��	vL��g�qG��J_�*���C�����GKF�1"���{)��
�<�5$��"p�k�pH�Q(���_��s��L\K˓��[�$׸�xe�}T�V[k�h�4l��6޲�c���~��H�>�P�A_�^��Ҏ�4���~tqI�`�*jE��2z|�t���3�"�wx+%�����bA}Q,K�	��ǜu�k Z�f��/�>��O�B��&i��l4Op$�J磟�
�vY�����F+`�������g�'����|�Ѕ�γ�/lU�_d/gt&��yu�����[-��QV$d�F�z�f5�V������S�Гw�j��靹"W@��V��ի�r;��	���N�H%�S��Y���B��.{n�z�6���5�C�}����&�w��#rۯ�G�G[��)1���}T�A�Q@��9ߐ�2V�g^|D�&l�!�uG��`됵�!�T� ��XEc D��f�\�m$HY�Xr$g�P�w���`r����3.l~�b'|E��X}�\gVA�˘����Fzx��;v���`ٟ��"U�:�/�M�ZҸ��8@a��M@�y֛ﵲj���-ȯT{�lk��������\0��J�Qf�f`��K���v'�Xf��>M�y�ቃ:�sVY��iFõ��Y߽79�Ý) �q��;��E�����GqH���h�zE��["3^��[��FӜ��w�#G��$����	!�yQ�e����R���-B0}�rc+1���W�V�4�Z
5"+`������se��
���b�Xý�/�f����[��	�J��H[m�~��#��t��2�����0аd��8M��G�)l9M\��y��35�?ذ���C~���1bs���j�.�/��o��0; _�O���������38�vC�Y[x5}H~�S>+�YmZ�r�B���\.�b�3�Goޚ��D]�B�俍&D�$;S=<j Z�	K����P_��7ik��� �N)e���xC\�	��h��B[�Ñ�|>���abuawz7����Vq�V���h_m��N��e/'$��뵔��ڽ���)��?�kFU+�%� 	���4Po��uc�g�Dj/�z3cŐ��ً�?�f}��~U�l�@�F�y�WLR}�7���/�i6��T)j�x��DgP�D�&�$hh�M%v�邙�1��y�i2ooz��p�ͻE��P���&�i�q+]J ���;���	b�,���~F�z �khj��@��ȳC��'�aT���̄�vw<�?nǌm��޾��ͨZ	���΢�u�h�$��tW�q�D\� �O��C������;.�;[_�X���:��bмR��G��5�+e�)���og���_�Jz�2e��3�����)���Z����o3�ԞfQ�;��Y
F��&sK�֤�o	�CUa�Ӕm��B'`�����yQSV�����as�a�@M�4������+Db�� ��;<)_3�ںKT�\�V �@2�3�A����s�� �@c�%��+(��3��=Z�x�2��`���l��l>$����#I�=�x/~���-��\km-$�j�/i�Z�V�=�������Ĩ�Fh�7�����̻�&��.��r"��PzdmwO��]�=7�jf.���N�#���i,#�AR�E������ؤp]r���?!��j6��+ؖh9�4�y63�$��㈎&��.���^.�3�5��j��w��b�V�T��X�@�2�h��rSC��ɷ����+*^�I�LXRb�Pz�>2|�۸�Pi�ui��V�<2 ��� f��.�Fz�Ց�z���#0C,�B.���̀u�����$Y@�	`:[��!1q%�3�1[qE����w�_A���q �Ql���s1��߾c[����\V�ɓ��nB����$���?c�oO\&ذ&6ߑ����#j���zI`џA�����~ޓ�"F���y`g*�����6�� ��f����\S���X��a8���k7�)n{]^<�z����Y�>Pm��߰R�L�=�C����&B����O�:Â��m�n���� p��#m7�����Ň������T��)�
���6^�H9�No���x�kDNt̏�p���k�������YK����l�0��j��S�:y�� ���E��ŭ,�p`�9U��^.eBn1�NX�~�jE��agB�y�^��Ex�"���5<C�^�B�E�d�ͮ���o�_������J����#��7T��TM�k���ٺd}b��n�����7A�o�w�΀A�C9u�A��m.	�v��њ@��
!�� �*4e��
�f|hGh_�'���h�|I��8���d���=0fu��%�NKz@>���όC�l���a�!,c����Fe#uk����I��W�8z�GBx�6���� 9͟�pAW���]ƈr�jt�B@i-��-aЇҨ�e���|�������S�B�F�}nog�+Sp�U핟��FH�3���3���Ȯu��&�����cX�V_YgT��T�����kL�h�'�ː�������\ �G˰H�bn�S�S���T�t_'�S��I��E�)R��y�7wRv�kI��v�T�t�X��Ԋo���3qު����)G���d���R�%�Oic��c���X�7�_"F�UV�
��(���?�io1�8�a�`��o$�C le5C jJ�ɢ��(�95��w�h�B� ���Y��6{ � 2݋y���a���
Tg��_�-�^���c��`��a����BM�(����ꦨ:��KIf��W\c(!���Y�ނKg@.�IJ�� ����Kʡ�餉Ɂ����:r�����	3M�y�ܨX!�/&�p�#Ӹ�wbq���g�]���9��f��Ɵ��0�q1�%��cn�1
r���'��;_u��"?��B�?6c>ǘ��2�I���^p�xӓ�Tq�Ȓ��c�$1��ͫ~�3&��#O�L�|˘���]���O����H׵�=I��/�[��o�U
N��e�#Y��;6���V�d�q�l���\KQ���g����l���Xʘ'Sæ8�l�ĳ�3-�oٳ9AH�t��������G�ٕ��Oœ�O��h��'��>�W~a.8���~���\6����i9edo)(#�7�u��ᚌ�\I�D�4W���|f���j�s$~
�Z�>r���O@TYݪ�𼞇D��f��f���E{��b��t����.ۮ���|n,�� ƞN���47C�T?3��������]l��Re�.s>Xr�_>�w���`�A
'rQ�D<��?�s��/˼V�=!����xZ��Qk��"4�5n�K�A�bR��l�*��'Um{ꠧ�X���������.����Wn"
��g)��<R��v�s͸�w�`����,����6EN���߳�=�T�.f���fme u�Xz� r��$�;���^?'��T� ��Otv�r�Į�M���v��7����W�A�x�Z��Dp� =n}��F�b2����}�����X�K���r��2�q�>�&28�:�P{:.��rL�]��'�a<[�^9���\��-�0Z_��3�i�v�2'_`D���n�H��H���3U����|�b�6�{��LbR]�*��B�ګ �Ȁ*��E��q���e%�u��ZЊ��X�BE����r'�K`��k�G�ئ�N�E~x��E�rW�"�-ŒB�$��fI�`f��q+�|'�-w�
��c����УL�zۦ3�`F�~t	��������.4��Xߧ
�$)R�&<��&SA�J}f��	V�=�"�MVlOZ"������vY��H�iW��g��v
��ȧR���C>��{�y��+�@ہ�u���B���}��k����1-f� b�<�_�d�p�P���&@�AɽC{����Ѿ��#y���+�G���zY�.l{�N��0O�A��N��NJ<����a���a��I��G��%�4��Mz�r$���Q@3ޫbETc�K3٢~��a��ϟ1�+[&����m�1��Awu�M9�����"ߝ�y��Ͳ~�Ըʀ2<�Z5\�}��g�D7�h�����*�UkbҾS� L�R+iS��ocZ�+N&t�y��A(�^� �'�L�(]C؏2��~(9�`/�`@�i�N4�2T��(@���B)���L�iA�-���.��'��T��O��7S�Ҷ^�(�t;���x�AЙ}%D�t)э�B�AY��z^����dzf�e\�]}徛�)T�����(��w�9��G�E2a/!hã���	eGQ_Y�F�NKBsh�yZ���ק��MN��8��ti�`��0��\�"!�r@���[P�b�w�D�X<�ݴ~��{k�m���ϭ[Ԗ�-�I8���ao�[���L�?m-�IK�\�FFƋ&�����B[mF��N�b�?9e�m���^��ha��;hEq�=��$/��_C� ��&����=cl��^�1���HC��Ե�-݁�="6N~QHP�+|�buAg������/��JC.9�C�=��)��N�!�w�g�j�G`�K�;J�c���詼�n�x�,3z}ey����Z��Gac1�B�P��~�����]��;HD1������	����a�|	˪[Ӎ�>���Y�Np͔`@PA�-{GD-��{�>���	��7��H\����
��3_�ң��C�ai*v?���U��^ *O��
�;B&��'����	��p��
r�����Q0��i`a61~�,��;��I�2�b���<��t �5�k���gAz;�#���P���"���QM#-S�r=7�h�K�:���������b�bG���!1iS�4$�Y08>��"B]�`�A��!�y5/X�f���%:NO�A�C�ef&q�e����G����I���b�%{�2�����Şo���1��ȑ��m^�Tw����ȦU��2ֱ��е��^�K��
����B���:��9K�ۣ��l�>��<��l��f�m�>-AWڂB�z �@���v��@����;�{���.6�VO�Ʃh���%8A�<K�DPW}54���$F�L�u����x�''8(j�E�_y�Vmx��>�i�[�UPܮl&�d���n���"��X�r���xVe�)��kU�w��E�3(�s����$S�F��B6.�ov���⌥ZhI���V�Ha
�ZMXS���p��G�bNd>�l|O~����y��-0�jqn�k�m�V��'�9yD���b���Y5�,�V�����l:�WE�e5Ι�g�$�ފj��P�λ{ԟ[����@��-���a�0h�\<o���E�.+�K�7���س��;���+�ł�8�q���d@�f�R�}}�����+,|h��l��iH�l��mdj�� fm�iZb� ˠ��FX�lA���އ`��J�����pk$4��cx�n�g�&k[g�<�#�S����`:$ �շN����@X2Z���f�W����#34�ܑ̆{��8����6~�(ax��j��YG��ka���!j�-��Vw�o�)�c����.�G�'��F�����Z����^���/X5름� G�0O��^��k��n�f3}t�~d�HV���6�@��y���Z������ĵ�d����<��a91ͭ��1wY�RN��/����i�ۆ4<T��#ذ�c��U	�ǌ]2ʮfL���Z�7{���c��VeÖ�2�{s{Đ؅���PmOb����L������%c�)��g��HY㽨{H�F�1�c�m�c�4�$�쑟&�|��+�Vd�`�4��ʌ�>��v�y�f\��x�k���D \Ɖ����oև-����/��9�?�C�W|���А@:�6�g���?aJ��O(Q�߱{���x]���s&�Ʌ�9d�\���M�(B8�����*Ԭm6�Y��R��m�,��/F,*gːm�#bkƇ	�u������[R�P�}�|��Z��Q��
���\9����5E=9�ʶK>g֯�#D�@8�t�~u�4��~}�Jay�%D��7g���^�ōQ0;H�@{��Z�YC��?Ǽ�r]T�oI�x�ƞC�f�)Q��b�(�}J��=�I�����/����*Y�����Ĥ�8����3�
�f�$-�27+c`.��LBM�&@G��H���W'��r�g��ab��8�����A@�}̽g1q?��a���!�i/��A�҉=�j���UFi������K3��%.��,��F�)��3=>���S�5�dM��6�"�v��R� ���98F&�:"&�A:|�H
�e��鷻�[������{�3D��Тc!�/�(m�mx+�����g���:�'�2T����HZK��9���Bۄ4>�fٲ\�7+$��T�uJ�UߨC���]�G�<���"9��9�_b	�.�Kp��|� �U��iT�gh䒖vDna�������+�i�*mp�*�1�㙲�;��\�Vi�R}#cn���l�d�|�q�����>4�p���w�s�W%��%��3�~�:��9��� DTح�"�b�z�,�y޳�wr�)t�IB߿�D:O��G��H�;��}@�����p��R��^�g�2s�0@L�J�c�?���:��:ȕ��F�k,
��,q=�1�y�[<B�5�K��B�h"�p�m<܉�H���6�e�ٟ��9vd�aU�%�CWX }`֏X�Μ#p-&�A�A�ޠw6{fa�0�����,8]?�5 ���ر��&_�Rh:KWć������g�T+/������@����H�r�5����k��Gg��
A�	�:��s� 0��E���~o	�/8��.���%���o��y�S�c-���+F��)�� 2����߷�8�p����dTj{vbN�$*�Q}���u�ԛ��V��3ngC��e��U�m�����37p���/?mU�F�G��b�0��| R�TE�&����aٶm7ü���]:���'�X2��ɕA��#$�_�g�9�u?�Mq�~�O������ ~I�Q������g��Q���>�q�Pv߽�G�X�D>�f�y�[C�k��?&e��14�]FL���o�сP��N�\�������}��`���V-"Q:)z��9�9��Y��<sk`Uk�tZ|���>�-�qO�)2,���c����zxd�
-."g	gMv׏)Z��j��9+UN�E����ZV���6���`{�7e��&��"ۆO�xOl��X�ݓj+��{�L�S�GG�%��`�.7@kS��a)G$�zfUU��<�y��*�J��Ĵ�7��0F��ю��S<u�9���8q��M��Z�/*��+A���n�Sx��*��/D�Mߤ�E��I|�^@�����p#��L��KXIҊ�DԄ���<e�������Ȍ0�����] �qvw�F������ɞq��:"t��5�6tPh�N��"����P�t3�5�E��g~��?�cv�Fnq�P�V/�c����4�O<f��	Llv�)���=�֋ο��cc�@IJ�s�lɐF^!���/���&�XE��L�,"N��M^�▤ ���ufXHnsRa$��b�����5�4|�B�s4����h�-$OՋ�8��O+tV�`�E�r�6��Ւ	���}�8�s�3���鵂����Ht��zYz1������u��w�w�՞6 ��y��T6�F�T^iB ����b�](�s�{�����jKP��	uo�!���`hB/u���g�w�0��|�u6��n��}77G�Z�M���%�C���76��W�f�#�ޗ{�����oY�(x�����I�� �s*p'���@K ��@!uD���اA�b`����.�,.~G�b[�_U�S:��[ŊĶ�ȡ��J࡙%U+�Ĉ�(�T��b�*FŇ?��5�X��{rE�����n5�Y����2r8�`K�/�51� :��/������y��6�Q�#<���P�Զ�K��!��]'�k5��5o%P3�_�����)BI�EcRɅ	Ll�m� >lJ���h��z����M�ه���:��1��� �e������	A��c�(_�:x(�(�I^,�����!D�X8���L��p3��f�e�4�@K��6���-un�S5=�Є�"-�1�".ycsmj�{�ۯ���4��-�	�<+�\���r�`��'��-��Ws���fF,�qB�}���S��?.�e� G���Y��F��wNy?#�Xm�p����i�ld�W]��A&�{��� ��xz�⭸�mN�)�$b���2�NΒ��R���*�o�g���wo���~�a�^��.Ue=q�'��ك_`�n�������z)��i1�q�z��Y@$���{~�N�J��p,���q������ƀ�b�B����B�W�c��Ii�I�QRa�*��J-��dW�2@���??�@�OZ>z�iJ-�D�O���f���#`e�������g�T�1�TE��=v�d�·�oT�=��q:�m�w���.�P���@߁��:b�N:�ĉ��슲|�:�.�l��:\�_�w������&���]���X���o��jVŴhc��	^�f}�ś����yu��o�G��K�ne�"���!�7��MP{�6�N6٘!'=���~�M�`#���n�LB�?�eh�?F�~uk�p�%V�.�4Ja��A�-rY^ ��y(@N#L�ɍ6Q��F޸����7��^(��<�P��\��@Ξ	:�hf����z���7���MZ�u�Ց�l۷ d|�Q�2��&Ww����՜�M��ud� M����Kc�,4�&[ b�,��`(R��m=`ق�a��L��K�ͪw�Z��� ��CE�"�qva������(��L�c�|���QhJ�3j���p�d�Kf?�S��ĩ(88"�A���$��������d��ZE�$=>�`����U�|�������X�&+�G����n���9�B]�o�+r(��n�wr*����y�C����=cUSMB�%��� ����� 5�tFb�]L�+�DlL����j�t����q�Y��.bB��?�=�L����'~�'����qG�WH��z�tK9�/�}��tW��z�����H7E�못YZ�.�b��4�mT�V��ѿM	=�J����zn�n9:�x7��;�ƍ�߸×����4/�}y��y������Zu"���Y�4�I�^�h`�_�p�3��W\�`	ܞ�ݩ�����a+�Q�#�eN��h]� l�����4h�P�4���d1������r|B�ܒP�m�������G���7�/�-֌���>�����Ŵ6�ſ���d���/!��["�K��f�(@��	�����z""՞�İh�S��#�$��m��H��M������>H�X�@�:��Q�&<4Aq��H(?��C�6������A,cPAY��6�BF�h�	�D�T^qD跁Bw]W#ȁt�HQDh_�֌�H���H)������
����]�mSMQb��% ����W�<��y��?=��
-;�e؇����@���P��������}�DP>6�0,CT��k�bŐ=аIΌh�D��><�X�E�O=��Ʒ?��a,3�.�T�S��~��H������0���'�4>k��v	���Əd(�~�Ja�g���`֜�,tZ��͑-�̺�LEd3x�Z]'�w˲Z\�& ��x,�5�hݍ(����P=5�|���+�'�x�̔b��N�1m��'��q��5�R'?$�2@3C�IX"�U�"X����aK�0,VA|�=jN�ʡ�N��\���u����u���e�&�>���F봄a-l8�%y:5A��#u*p��Us@X�U3��9v!_���J������;>���D%`����0ih�Y�������4��l�O��GF7ɾ�d��\,2Ǫ��E��r�	����DD[���`�[9I�y|�0O��m*hT�b�r�M�w�XՂUV���c�EZJ�i�Be{��_px "r��@��#�)�3�~(!n-�
ݞ
�ǃ�,����/��֟2��g-�i���_�R��ۄ�(Ӧ ��Չ�2�MA������KTx���2P�s|~�%&E d�R�&sHw��礂+i�K�a��_^/d���;=��3��B�Ϳi��p��΢1:�����ײ=��OF�đe01�kd�Kl!���h��@mWؚ�W��!�W�~7g�}�� FT����u�������
<0P���xCJ��2z_���"(60��Pdk{��_����ܐ0�:5��<yRʲ5c�k����%'�I�0�֓�?+�̕9�L�=-wnqI��^>�E�;�e�v�����T�t�u+�����k�}
6��{xʐk���:xi�~/������{=�W 5]�lpS@���	���^֋���B]Ҭ�r想����8;�"�%>r�Jُ��Bm c�9��f�q�L��.��wt�@}�zW.��^�"��vy�u�#AMn�$*EǬ��:��3�͈ߥ�Z|#&iW��\f��� 37Ta��А�l�,��k(��:��0�4S��`�6E�1�x\����:�_�6>��X�Ǻ�K=M��|��������7��W�����ݺ�ъ=��+y�5^g�F8dU�0����u������-�*��� &�P3<�e#?b}t��xH�����XQ��t���EpG�-j��A���iUޟ�	��c�2�sh�oMj���3[�g�P��Y�ɵ�if�S-���1����&XJ���nQI�af	0��&��o	q5Y���~�*�p�����ݕ�(y��l��~ʠ��i�Qõ#��O>h�qߌHS�g��%fW�
��
����~�M��Z&���k
��:����A�UohL&e�8���MG���/z׼
��^��z�Fz��b�;Hi��$�(�ŉ�*GG�&Uf�B�Ƃu!�,�1��B^���I~�?ۋą�Ҏ��3��~\�x!.��-�m1�w"\��8�J#�ХZ��vzTfĎ,�����R��;X�Y<��S���O����6��nOV���:���ڍ��8�^��|O�if�ޥ�"Q��u����©���?���."{Wr|�I2����a
���	W認9&\�P*�äM���6x���b��g5Q�D���
�/����$�HA��#�)���P���-F
�ǹ_�O"4S `o���*Hrr�m�d9�*���[^6S��K����J�<�I��!8��V�|��K�%�7#u�F�R�+iW֕�f���\>6�p�G>�h���X��JbiY��-�&���//����>�H#��t�o�c����
�rD�(>N�笄좦���]�f"�hoЉK�®&��{ �-х�I����CxÐ_�Ql��l@�zv�$�d2v;O/kq՚�k�^o��o����H�������%��"�KE���^j8g�j3���<Π�-^�2�d�~\Qf�{В�W���SQ~ډ �F��;�-�/]3Y/pt�c,�=e`���$Rmdt��}���/5(�g�V�jI��#��z-Z�&���ü��F�Á}�7\��`8���b�	�P�H� �t/2���*jY�R��D�N��J�a9u�\�)څc. �a;-��޾6�r�T����mZ�t���K{%�h�u�h`���]l�͎���'M����x���oP�SZ��
�_c%��X�x��|f"�⩫���d����4�+���<������Z���h�sD,C'� z� ��޼Ȋ����y&elL����P�q�=nf��O��[�_�_)�m�ҙ�2��QQ�0dDccJ���]`<����X��dɡ�K8���W8j���I-��5�/*J����8zD��z�p�;��#EIb�"�!	���O��1�$������s��������m�F
�D�h�r	���O��qR��5�٬#��e+��͞	T*"�����M�p�~��뇥i�
�A}�bY��a���ɾSI��OX{o_<^n��b+�-K�jϡ��Ҍxt���H������ �UV�}{��svv�� ��;c1n��*�>�ch���v�-����g^z0Q9�������ُGR��t���
d�K�B�|�>��_1ʵt�T�#��x�HbH�o�LD��?�%MG��t�S�wl�m��M���Um&�r��� �1c�q,���09�Z�����qu��lS�=����V�K9���J�fhn����bTȔ��}) ̖�Կ��g{d��S���!Q��� AA���(4�{�����MĄg~��b<�Q�]�e�z#�D[[�IM���{i�!Q/��K�{NdNl�9h�e}��/`ů�����c��7�sԪ�2SjYdOk~|W:_X
�HOe��ġe�x���7එM�[���W�``���M4u�A7�)F1�VQm+�j��Ph���񪕮
C�J�{��5�xfx����v��s�/[�ѧ3��-�9�h��J��U&~?������`�+��4�t���7S4��*$Z6jt��|3Z��1H��i|%6�?�h"Ş��3Q�VL�׶�SO����Q_��&�cX�0��|���Ʋ�s�S�^��9����Ll>4{Y�g�	F��f�*�YO,g���^�>��̥�+䓥��^�s8Šd�D���Q����Z����;�J�?�ب8�Cݶ& \�yx�5��ǝF�Q"��֧\'��y�|��m1�����W��}w�n�-�F�\KG��TU�0_�E:c_\���/^fC�0�ږ�V�"Cֱ̣l>2ޯ�)��MK�y>��t�� *Д�~  �����*��x��X�D���)�V���5ܖ�LC7���]�ҵ��=�SH���[!'@��l��@f��aƖ{j��]�{��=�=��%��wZ���e���5��)1d7�be���n���='��m}�
�M�_(C��t�(U�����u�t����k��r��A���_A^�'g�ݬ���b�vo��-<���H��"e`����%�|6,��$g��R4�;Dx��@�N�� uD��0悿��Z�(��B�n=�8�;����/��;���	�\zvM�J�&y��0�,O]�ة���'Q ����K�7�̼�����ޟ,��a|7p���ψft9�gm2\�8�\�{Z��R��l�bʯ`�\0�d��*����}� Q�X�<X�#�����.w�'K(�R�U��A�yb����d׈���E!
#�Y�f�Ci��#��i����uL7�>��z�/xx��*O7p���I�q��w��X���auYY��J{R��H5)v��ց�T�u���NH�����C6ؗ��D���g	YL�ف���z��JǮ7I#1�;�U_�;`0����m�ġ��U�  ���|dj#k���r]R�?�Z]3� H:?#ś@��ya+�W�|�^�FJ<(��<�4̽%<m\�������t<^fUg��#"=�<���������B��7gd�a���;��m�Í��Vga�N:����F�#e���^�D��Y!�p]}M
>u��!]��5�ú�g�=j����V7"�;��`�aD5��E���s�������@ճ�2$z�:���^��gN�(BfE�'�ֻ�՚v�Z��nf���V�QZ9W�#΢N��$]����7,y�������M��\ ��|Y"�F8�	��=22�gID����������bȖ<k�d#t��2`ǭf�4 �&�&��KѶ�#~�,���Q��q#�k�IM~n�y"Yiį��N�i��T�GH( Uঈh:��ϑ��&��ɠ��MŬ3Iq�NA[�Ƕ���2š�_c�"A6�iũ�4���
����@���q=��"L���;�0K���ƣ�Ӌعp���DFn>��@`���]��䷆Zģ?���v`��T�|j>�gg!��]�\��*�^Mۏ�'I����ϙ9²	�g�8�����]��8�hM+�y�_����`ʗ�\�x�_o$Z�X�T��mc���Yb��{���Hf�qP�C�Ծ>�|�v��~��xӘ�6�p�y�Rn���P3�<�l�r-PQ~ #��݂f�A�M�^kw�Uti��e8U���m.���������Q8d<�w���j>ZTI\�M���{!N�[T�WϠ�Ya+w�u���F�c�bP�ƹ�K���Q�b���Y!<��e�1mY�v���[J:������zy(Y��q��S��!Y�����T�����Cy�X���a�^w^��t8=���(��[��6�\��Z���\�֏��Y�x�fV�}�˅�m�a�����S�y{�f']~����ϳ�پ�4��'�2�׉�׃dz�`q���]Lb/�H��3�����
`4�1I�{����ˊ�>!�!��( ��E���\�;�)ޮa�}L��[f��տ�AW���暳��l��� v�H%ᴧ��`!�j��^�����/���ml%�=�Sh�h!��V��t���su�8z�35�=t����H�OIMi|�r�+}K��$��������ͼBO�׀�N/g�<X�ABa��ۿ�o J݅��O{u��O�y�@Y&ŭ�k�"�	-$'�E�$1�7��0s���&�^��`ur:�|O�w셄�hlX,b|x�PI|�P��B�8�rZrf:�Ǉ	�ܩ�Ҩ��B%O<�*N>���,|3[�"��L��������j��&�M�u\j��C�&G�M���GH>�C=<j��v�ϚC�G�>Z�Q�/����#���=�b'�!�h����2�Y�I6l.����h8���������v7���w���Ƨ��ƱA��
g-΁��Q��lq���C�Y��Oy�1:��ڎr�W<շ}�{bԿ�`}}�a�<j����ǔU�U�y��#�^�8�����^6{��}����=\��Jْ!��-L��R��s�9�6��oj�S�5�e,�h��u��Ӳ�D��'*��W�^mO&�Z ����_�M}�^��*�-�&�Ch4�.A�B�'� ����OE�V��6t<���MNB;a�iLAp>��k�ǿ�EhM3�:��Ռ��*
v>fv���J>M]�5X(��l�^',=j������󳋧���ߡM�����2����\2����kQ�,9���0P	��?�y۞,.Ǧ���rE�ѵfq�����y�"�ި�C���q�9Z\e������6�5�$DÝ�=ؾ
� l��S��f��2*H���Ÿy��뛏\	}�[0/��v||��^�M�.�<�Z��O'��C!/5�y�����@���9���C�}�	�ҫO������Ga���I�9{'��;��h�����Fݶt�RѶ�MZ��<�?�W��9�Ξ�M<�)��L�������h��a5v=lV�����GRy"���i�:���<|�ɋЪ�����z��W�[�1!�G�� ��N�3q�<����P)����[�=bL�1\�NTw�EJH��{3.�Ҫ�i;j�i���Ů��o8����Ɓ2��L����a*_-�a��砱/5\�T�����dª�[�"W�Ga������vm�z;��þ�ֺ��f�y�j9���v��jnZ��6hl�����T8"H�E��lE8=�/li�A!�ڸU3hj�a��'3KJHC껷ǃ6<��
Ґ�_�k��њ����m���A��R<��7S�`e,��C�[W.��:\2����A�~���DC���E��x=Z�F!��~{�z�R�G�c�=E��/ݱP2|I����&_�=���:+h(,Ъ���8!�=��������g����rlY[��XH�]����E�[�N鵛�l��vf����ᎀ t���+�;�)��@ �����!����6=����4�B#�r�>XX���Y�&��%��U��O��2���i�٩��$x��N��3� H�>�G���盵�Q�;�����},<����r�V]��G��ύ��Z�p�iǊ��٫6���EF(ޠ:����G�*������	%�vw��D��Qkj��[����*^+.��<P�����b��sDLK}[�J�:!۪	
�N�<�#!S΄F�����G���J%�\z3wz��o�]=K���m�!�g�3��T���й�&hk5��a�����W�v/��)¨�tt~����Þ �4(�1��O�o�hbR�W��C1�$��(��>e��NqĄ;�L�N�ָ矩'����
�p)R(��g�5�Տ.��9Y���-��wƖ�j0�."ۢFI_W�e�F�ɪ������=�l��i�`��\TE~3�2����Ec(%�(���1�lk�#�.֋�7��m�HWt�(L`_Z�ˉ�/4+���r��퐷�Y����ό��Ͽ8��j'k���s��~��t���Bq�z��RF�}��l(y]k9�Ԏ4xԓ���!���Κ���>�9���� �u�I���w#e�@��^nL�M%�
�Ihm2+�&������	�>t��P/*nY�m�8�}�L�9-���_�D� l�	�Z�� ;⺉�O�a7qF�*��KcLt�!S������mO!�:5��Z�q���缾��e[�ڋUmͻ�?Ν�\H�x� ���G�Ȉ��ʐ�����.��|u������룒�#>H������,�Q�q	&���l�?�*���A@`��r|Ճ�W!�)&+1�nP�P��%�k�t�G�+
v"l���W��8�P����t+hT�AE]J�����Uk5��^��=�ª�?���2F��M�z�ֿ�m�����7Z��\lЌxd�h�,� �$�H��>B�! �j�[~Xkh.�x)����6�?���2wyu���Cձ��x����W��p��cMB��K�;��$�4{J�W ���o���Q�ٽ�'��Ҁ�A�6����k��ƹ\���cM��6B/�r�o4���/���Rh��'*����OѴy�M��"�C-�:
0.,}}H$��-W%�z��;5�� 3v��75{B<�h&�˒Õj!Aߜ��\���R�c�W:j�m�����o��{Cf�4\Q1��>����'��㙃E�ڎ��N���|h\L�KA�����̿��14�X�]��-�ږ
_J�$WZ��+kU�F�5a�r�u�|Dc���M�_i�ݚkw(�h�P���\;�ޖ�N�&���Ɯ	}V��$̊�:Q���2���%[B��*�����#�t0�I���);�-�.Y��<����v�ױ�8��hG��A"x�U�H�f��2��/�+=Ca�їx3��>���������F�5�Q��_��t{�;��i��� ��(�{�;t���פ�'D�wI��Q���"ޗ�e@p�����4���q/��t`:s�]=�]c<����ܶc3%=�zת۝O`>�z�@9�ez�:��MU?-���C�L}R�<5J�s��l��Y;����`�qM�3���X΃d�c}�Z�TJ�O)�dP�9y$���!����(���αGb���x�������$8���{
h��[)���ީG�yR`��X�C������'�*�Y3d�!L�+p	X�%,dk6?��C/H�h
M|�m��-*�I��5_<����F�]Dc?������3�Kr����À��Ϣ�z��ߩ��'6-J��%���PG�^�`%9�1̡���֠0�_e&��p>��E+� 6z���>�P�n�K6X*�2�3���J~�>�f�|�`��?���¾Ay����j��켼Xo��PB��S(,�m�M��V��o��M_���M�`Co�e�@Pij�4x��&+<����Xm�0Sh��\� �s�G���>�ˋMፎC8��{T)cL����j���WöQ�|�t�5t�����ˡ3�%�xFN��K�X��F� �X�����{���&}��b��_�y��;�t.{v��?�m/��F�-�]@"`����,��NJ�e�܍��!d?��=��ANw����.�k`�N������ �'�$Q��$=w�����.c!Zj��0�*0�΍p�uc��?Au(�h9�;��[�m��uK�M���0�'ԧ�3>k��2�Wi�}燝�3ϩ'囹�}ۼ��||�6��.Rg�c)qg6"��ґTp&����Q�����׎i@�f��&��yy���)�^�\I%-�:�3�`���t�n����^�6��������qߗ�߬#1T��cL���Kg����xw"ڞ�bj5.w���2�2a�9H�XUn�!��>��oGQ�CGEٓ�o���@��r	��w�G�;��`�z�?kQ9�I������7r��\��ںҤ��a���+��2���M��F�m�Ï�=J�?����2x�EtU�j&-�l�oZ�y�'���}F\�'ݗ@H�D��;9���C<��(��$?Hxd��&�A_����V��c���k� Ȳ�;zl[�W�,�~�Z�N��R�'��&?��׍���haS�5�6�+�Sf��%z�m8��>W{|������8�R�A ��ԟc ����|r�%O܈W���Xpo���iƁI=����r�i:B�L��o���,c5L<��Z���p�3v\[�]|���n�-$n6�ZY�0X�Ƨ̤AÍ�G�ӊa;�BH�Q&���iH3:D�D���	�����1n�b}�1�+��G��b��lLBQ+�7����u������JQt|���X�
Lϧ�qJ�'��%�Rc0B�����E����Q6@�Os��V{��썦��'�'&'?��ᑬ��әq]2kHz����Ҿ��'�J���(�]ݜ�(��Z�Eu�����KG��Z��[�cw4Y��^>���gt�d<�S^{�ಟ�V�������rX
�ri��-����$G�*�i6s���㵊r��Ӓ�c�a/&ݼ�X����>�T�q�G4?1sO�s�}�j�r%â�Q��:0l����]�t���7�:�ɰtHDf���9YwK��:C: }��rK`3}���e��G�u��h+�e@p]�b:��氖׿Ż�w���L�T�k�&�Ʀ��e	DL;^�G������7e�P��m� `2��AY�a����<�x�`_���$��Ջ��)0�5�`�ϐ�o�|<���Bg�'yc
6�y�LB>�~d����1�u��Y���BuE�&��P�	��c��z�@d���rM߷d	ș��Q�� ��G��TNÓ�,x�S$�@��s��_$�k�*�q��ǛDA��ll6L����yr�ո��P� 4�I=&w3�mu6b"�h�r+���^3�T���Y̌���!��C��K`�K���W��f��>�A���$�r���{Q#-T��>&N�s�t��p`�J���w���qC���4�<q	�@�5pҒn��,��j���닥vj��=%/�[͸����2p�������6<xj��_�|>�âzl��^�!�c�҆���\2��y����4��R�0S�R{2�f,5�h������rK/z}{;�Q���D����ZbIb_�ڵ��
��pN�у\x*G��HM>~`Ť^c�0j�[
.�yx��ӵ�UfJ�_�c�eφ'1�n
}#V��`��0�Օ��M��~ܓS�0X���C���I���>��mӔՀ�Do����&���f���/�r�V�u���ݨ�Xz'��(7-��[Ho[c��2�;�!k�O��я`�;e��3�p0�GN"x|���I�R||���}3U���"�T&r8�X�7+�>��7�	(&�T/\�����K�K����&����p��Ze���9$�y��_���I5e�c�sV�kL�є/.�ލotR��Xr���M�?7�w�,��6��ib��x����%M*pO��K�V�n��nT�{(��B���?�S��bF:�阉>���z��SKsi�r��Yd=])g�c��
���컐��ݢ
�$���-Y���*�j�[�����6��3�e^2��ݺ&��ȵPYT��
�� ��Q�Pֻ*Dn+nE\A�A��{�m�����Ezm�l�|Q�_����I��G[�ɱ�N>���wQ�-�xmq�kcu�q%��0̋���!��q
4\����NQ�`��y���j����~��W r���W����y���U��@�U0�C,��x$(����[�N�׆���N�qF�4��C�Ֆ�X�J1`=�����q?���}j�����zY��q3��Cff��M��F�~n$Y��[M,����*a8ܼ�_�;'.Ɏ��t3s����wv����^{�!���m�hDr9CS�gCR7&#�)a��|U���gJ��}�21D*�L�D�u�Aʇ��,��؇�ʇv!�7򽌔|*BFWf��0Z�`�u��
%òN@�_�h˖y@"j��x����e ��- ]��%K�R����n��̭�3��Gdȃw�a�>pc�����Ɏv�Hs����5QY�t�Ĩ�$
	��I��!u��Af�������dm.�����^*=��Ϸ�nbU*Wf��E
�蠂��l�r��ʎ-�D�d|�QƝ�
���Rnpe�tT#�]����j�<�B��r{.i�\h\��r��jG�}����R�y�B��Z�|�C��;Mar�%��aT�p�K�Y�*�@c���@�~����`[��u��^��կ���>)�A�eTN]٣P=E�4�7�O+aH݄� .����C.���	-T�YDfd�_�]p&�x��la�c`���.Q�F�p}Z���s���тZ�<��:�jkP��.���ԭ=ݝt�vc���ۄq������ڣ<��CVU�?���lȮ�+�26M��x����*X�&�Ŧ��&8�(�X���.a�ԩ�R��	���5+�/��E5s��ߦhɚ�����p�BI��_�R9@���M���y]
�(�"QlĄ�n�8�c��7�]x���,Քb %b�<�R������~�ޞ�t{O&�v�:�������sq׷����a�IC#D�U})�P�p�,L�K�m���o&V01` �1P+e���*��oK���J�g�ʿ�xJm�&��|h�6�G
�$5t�7��Z@���W�t�fKS[R�l�����1紬�z	��b�ob��$P�9�2.J�	y�9�?Gs��<m�9�!���T�٧6H(h����5�܅�^t
	��e��1�&�ns�k�>�9��z��L�!@^�_�Üߙ��W��NN����Geoy�/	��ϧyb�G3�pY�sxM�O6���ř)'�Ⱥ�1T\�.Z�>�.��X�1�d�V�Ș��QbN��0ke�'��F��9f�FIq�񟰎RW���lH�j�>V} =FS�}P����L�%�ok��z���t��Z)*����߶ǀ!Ey��C�������{�Ed:"�7����N	W!8�B�d�� 3�U��.y� _���xQČ�w�DUJ�N�����}i�4��޴=4@�M2V���`{�r��ɛ x�IZ�����m�ԛ�Q�,`b��P#���\lPF�_J/�-���`V�]���̆�lt���B��3V�y��?��\7�K�h2�Aa�h`0�'�q�	hH�ů��t�����#�y��Һ�gGy=�$I&`NK��+�f���(��'	%@2��`Kʤ����9G�,g��Q4U�V~��� Ҍ��w�Z��do�](�ӄ���i�L�rgp8���"��x2��²P�(�Õ%>�2��)��"�(+�{b�ǫb!�~|�#�J���������fw��7uU��&,�¦q���Y#^�C�ZJ�\K�~��zP���k�؂�:���YMR�08��jA�%3�a*�x�ꢓ��zCc}G_�~.2:���H�8&��{�A��Q<��E统>O��cn�v��4��V�A�+�~.�ZUf��Ǧ̀ �;'�C�qL6�%��{d: ����`x��J#ƠV�����I��Y��^�?$-�EI��>?��� �?�����de�k\
�8Zɟ�i?��M*Ē���kD�(����Q�|�3��<�����^$�����eM���א���&��Vb߻}����9q���|j<��[)�a�H�2��bD������t�NaB��<����ZuM?.�3�X��Z�� �<u�T�*�4�R���P!�v3�7�^��_�P�����po�0��+��Ȟ����V��Z�)ɺ �PJ d��w$�W-fP��}Vud�A�z��8?�{��p� A�=ͣ� ��́�R���/�Hdᙸ�k(�}��.��zS�d�_�A��@�ss�Z��C��-�O�?�`�L<��rc�Ɏ�\ׇ�:���ypr^�����M��=G�����}Zt�F�1�f���		�y����Y���aKI��[��I�;d7�#���FK0�J��p����g|�r�&��=�`�fx��C�n�Mw�g�B�u�/g�>1T������G��-��+��*�ɏ4�Cɶ#�fO����fY��P)��F��`�>+��񠗰�	sG�'��2��(�6ڙ1n�-����@z#ۚ0�a�2=D괷�봲��5+��m���!~�HILN=H�
���<c5 o����	���~�TB-GI���pT6o�W�F��W��ş�\�Mg)l:���j�̊�C��F��-�H_�z���W����^��v̈+R`�l����t�j^BrĂ$��\�L��0=���5QY����¦F�>��G��}��RNh��'���6������ӧRhL�V���e�N�e��}(M���^g��h�t�� [�3����@��ɛM� Y��?�r7 e�ȫ�/����&�z�|�Tl�U��+��J���(�r�"�<�,�ʤN��h�c%rz�C0v0�js
���X����n��Kv�,C m\��zkE?A$	u��c�5������Q�H�)]�GS��ӅZ`�{���UC)�&�A �(�Y{������5�pՊx\���C���'��"?��iI�Uƞ<8�Y��l �ڮ����%:��_�I̕Qߍ��˒�"�XQ��7�4�s����E�!��poڢ��3�|J� WH%'H��I��K���x6Ȇ�'}��3E�8�7f�a����L7F-�m\,��ִ�M5��WPT^�ׇ/Oc��BP%�[��S"�ꦻ�c�u���6�i@�����op��t� v*��DY�<��и9��2��W���W��7�0V߳�C�9U���k��_ҋ���g�mc�H�a�ov��x"��4P׎���"(����5ϝ6S���I|�]Vjc����W�}照����Jz2��RZ�3����nڛdbz�����G4ԇLYKS�rz�ipM���$ !r����&�w#�/�l���:����S=��">�:����ۦ��YT[��ee�+��hvё#�,<�D��'d�pQj�5_��e]$7��Vߝ��AwAʤA�M�d��lWu`T�c�~�C����K���UW\
���'}���	�b
Վ��Z޷'�	�C��a'ޏl�4�c۸�W��Hr�LJ'Z�q�O`CT��ެj��	v�|�˜:-�zⱾ
K� |�e�;��`�f1rqg�/�h.8@��o<�"3:��G��vj��Dz\��|?n�!=
���=���5�k�3!�fN�/Z���t�f�dE[�t�i��/av�^���^/�h���Z�����"�g�ղ�����$E����{v��#��
�Sv(�77�PS��o�NX���+:�L
�1C%M����b0����
:z���X�(]� :،��>V�[�O��"'�/Y�J}�a#�+ee5�Z6y;�O鎛�ˤ7����(�>��L�]Ǐ�Y�l��)+W��}�H�i�>��3M$B�	�G�Ķ��'��1�%~XO����Έ�FɲW���$����
���S1'�E�  �N�Z�C-��7&��徭��� 2N�����!��h�E��wDm��Wh�o��p��"���.�v��XC3a�c���S�� �K�愠�p�}�"HG4~�	�p}���$֦l]� �I�t%��Y$#í'n�䢛q-��ζ�	�k�J[/��y�߀�c{ ��X)��\�"QBA�T��t1�+R����������-L�����kϏv�C�$ܣF �\�j�i�>�u��S�uR'������$rkv=��p6l IډR��F,� _o�!g~䯒}�}Ao�?#U�OV�D������)����l�I@C�.$�7#�mUG��'���"�������p�$�;$M>C.�z�l`;D:l}��c�v�2K��-<>�3
ƆN>�oW��pX�qł\�����>|��O��XH,���� c��X�]�� nR嬸|�%ZȚg�(iw/T}����>�D�ZC�# �k����A�D�Ȟ\K��*!Q٤�Ot}Zo�2ge�������-HI�I��/�O��Y�3;���P�4т�B�y/T}l�I8r��cC�ٌ�a�+�
�v��t�Y�v�T݃�j��y�瘔s��E����}X'�E���6F�����"��}�4Y��Yz9nk������|��5Jόï�y��-�+3V�����F�S����9�$G�6u��c�z�m+��� �( M�T�| �I���Fs<��}��[	~}����w���Rӿ�+",�xr[���1��K�&����6��)G�IS��<����IĥIƭn��Xm������˒�t�����N�k�C�F�?Ӝ4��z6�q��7?���F\�v��z��^����ca�E�� t_������F�{�����x-����Uә����2j�r�P^~�o�K��3��t=��&L��/lv3��:_k���C��;��8��
9�ĻC�8��}��J�~S��*d�0�*�����{6H���E�i�Qxr}iqd1�B�{�?���C�ū���--�ٱ�l�W���9��l�X�7�7����2	@<��l��"���{��������E��Tt��LԒ��ۙ�a����E;�9�gA	��%���srr�e�A���LS�_	�Z��e�|��c���Nj]�r����A�+�[9��xv������������f���>����^�8���|�7��Y���{aXV�F$�d�XR�����5��C��=���� �)��ݥ�&S�Z����q[��C�O:�C�������Fڎ�,t"ge�)�)�� ���|��Ho�
��!:��z|qp����������O���]��J���;?�r!�t��9��G_%E�s7��׋I����&�@W��br70���7?j	�m�{�P(Z��F� ��3ru/����$�Z��
���zh<l��XAۜ�@m�u�L�C����v��A_Җ��� ��֕�u'n���V޼"�Po�q�k�*��}��������:��T��d���f��8"���/����S6KZL�05T#o�$1q�+k������w�U�6ǻ⇐!
5}��(���'kF�z��FJ4Q��ȥ����бZD���EYe@9,V������W�z�^�ަH�\K���#F(�0I���[F��$�>�7fEwySm�(��Di��c@����m��_�<!� $�l����8�7�!��YzF���x���24%������cF����'6��qb�$�E��� �9~>��ʶ��]�]"���D�ͮth�	? ޞG����z#s���\n��m*}���E"��B��Xl(�ږh��^[~�}���̥�W�@?ԗ�w�V�'J�i�nw�5�/����A.P�.���,��x����C(������������^d�_z��ھ��V,G�>���9ؚ��+�z7���0���	E��dTD^鰙��p��l7�n,Q��-�,D$+ɛX�8�[s�g-�V�{���t6�w��vb@E��Z�]G�ޔ8�ɓ�Gg�GK �5ȕ�x��]feμW�;��[��".+4!+0�]ws@|+���4P��4^�u���������`<�V��� ���vG;Re��78��:�a:�;�G��7Zߩ�7����k�9�L�y�fvT^WQ7'�6�J�Q�
͇�?��ӀX*ڒ�$9�9=�{���esg�+�.)��`� �F�Ѿ�-�g��r���6>`τe�F�w�w����`iS-��
F�LO�O���L�!�����Zu�e^�,�z0(j�9/zߎ		})AN=7Ɇ���=Z���T��k_Զͯ�.��.�i;�b�\ ){����
q�-��W��6AN�5��p�����9:�A��d�X������ B�v�����67��d_��ȋM��7y����hk �,����hR�&��O��I"��NF]g�A��}��Pvu��dp	�A�� �b��^���e" �<g�,ufC\��|۲F��ގ2���㉮.&өm�w�[�������v��KP8ShO�7�*�����ц~�ʏ���,�(��eIdR<�Sr�����E �ѭ�Cq6�c�W*����yCo�FkΓ����֪���rw}�xj��+��#�2N6���b� ]�Y����sp���Z��Q����IĐ��|�$���|G��d�hL͓�x��(�߱��t��}ԁ�(�N�|����aw��
��@h4v��E��ȱ�e(Pf`�9�C|_��[+p ��$�7�4R���R����FEvu�'���ޚF�K�N`��t�#&����t�V��9��W�](�q�#YVF|D��0��y����l,_R��?�T˧�F@G�3��M�.�7q�]��du�񑙿vV�@:���b�};2h88i���^���\�&��_bVM8��޷bp��KL������\ɳ3��t�-?���C��[�2�X���$����>�>�Z(p��|uѹN2�=�쿰81�BU���׳��1_�[�JzB��H��Vc�|�����O�H��9�D �^����f5�����]���4Kb�WC�e�^���8�����r���<��ƽ�C^���������2�(K{�Դo'�>��;J�`n�@Y��;%I�v��=
Sa�YvC-�:Y�7�o�P�S�$����4�����	��9���i�7``fO*>�[�6qe7�M&���6pm��w�ё�Z���Cy����O��ё������>0�SK��Wi�H���⫙�/G?��A��Rw�S۹���U�(�h��� "�%�����Au�Lx��\�oFmP
�zKZo����Y�4<'��8-���HN������\d8ͻ�1i�RD�8���q;,O�NCW�+�'���@��w}/}q����!��I2�J��d��nHя�@�i�5�$D�����rM!�J}�K=E([x�3�S�.-��G��͗p2�^R�gs�����7k�.[r2���
�N�L�S{P���e��Z�EF�'�A.�w�A�J���I���C����+Δ�8<%���սK�h%���hl'����X��;��̈�zgߘ���Q�t��VwN���8]!��H-C�F*�6M���s���P�0�����Cc8����)��Դ�,9yp�$x/��
/�D9&�jI)���W�*t��_����?��$z�������A�u�L~��a�E��#�Em�w�gvȲ�fH8E$'�F��-�7-NHe�qkU���K�*`J��pG��ĉ5��1��J�������6#7<����t�_��X�6�e��x�a��L!,ܑEޔ544���gJK3�zd<���R,1_~ RQ�o�����qI�=��,���!7��-SM�s�2^�7�`i<�uxM�[��3�<�8u~�E�k�_���."���NdJ ��o�Ax!-��Q�,3�;R��tF'��/�f/׎yX�IA~C��݃ܿ�RNV�5�k��t�m3���䘀�a?����#��~��q�r�Y� �%j�����f{"My�,N�����l��鴳9_�"��ME��:&0=�g�5��c�zAEG=�m�/�O�ʺN�����M՞�t�i@��R�:/'-r�ٗ[��͘-�S�o1,�֕J����@}g��oX%���VU���$ÉY�[ "+��Y�/75���j�H-*	�v�cY�ik.(���r�k��H�-��Nk�FT����R+��,	��`�[4\i��W4S��fj`�9������J՟}�MQ�[T�ʌ�.�8��t{���̖]�h��9�gk�×��_�(� �P�pԟ�!���]0�_;GZ�>�X2N�
=�t+5V� ��;s�m��c#�ߚ�}�.&)����CXgZ� ���<�O�Wl��Y�LY21�d��������)B�t�[�Y�5F���G�Z�zK��So�u�1a}L�x�k(���|'���մ�������NE�cS{i.���_�X<����i�E���a���D�Jg+eS�F�6���z���B���b������k3}���1�����PV�r���t���b�C֎�e���X���\�m�1�ѠP84J�r��� ˩�b`��ڏ��j�[]��C����&����ϛB�K�~٩ϊ���g����)������eU��ZҰL�b�8��[K�Xܔ�M;y����y���(	%Pt��w���"5D�6j�t�Qe0��Rp*Ŵ��nw	�������aB����ד�6��ͤ%�=�E���Bm/|͠�+�������y�"9}�j`y�za�$*��|�L&\���jL'2����v<��ׁ�nA�_��z$�r)�H��4������aּ'ɽctK�1�X�	��=^�
2&�oAw�Q�G���אr��ISm#/�m�������F�;�m�-wo���@?wa2��P�����1�{�ϒ���`wh��Ҋk����G*��%�a�^ɟìf�ƾ�v61p�C�Sy��s�>]�C}B�Fc��D,��=&������)qaO��x%|�Z$���O_�����H���VŬ�*|��}�V��R�?�Grh۝��`���K���_'�	=��,��Z�Zҍ��愑��E�w�M<E��F!�NXi�У$/ߴN�6N�%�R�@�{�4�)�����5�C`?�����	T
ک�Shq7�c�:�B�US��B�����W�jb��k�(J�ȄN���>�-K ��'���KJt�s)�p2�A+������Q���+	�6���^��=P�h$�Գ��Dچ��~@���ɛ"5z�Ď뮈��ܳM��*b������g��pۖ̒J�f�]X�����'��E�_����6�w�yb�p+L�`իG�]_��$��7��n�᎕����+;��_z��7�l2�*.y���Q��;�TMf�-���`g�o,���ü%j� �H7�l���3w|-���{���"��(Y!���1I��Y�^y�t3�d�GA�6�Y�L��P�������0xō�4�m%��ۯ���5�KT���:����MD��b#E�<�kыl<.97���}T8��L%+�W[1��� 12>\����<��ə����B������.7Y)|bwM-�KtZA�S{�=4��+cҍR���ZaQuI7&�m"�+�q��[���O[q?sB{h�(�n^��>9U�k��$�����'T��k;{��u���н�p �΀�R�,k����(D������QV��x��<m��������r���?�s����<��E�/?�t��GA�i#^��3s��Շ7��xf���hE�s^VU~ �ST�1pʅš�������u���l�;<�PL(Ƚ'Dx��{;��98S�@^�aak9�]oM/p�nRZ�8��F.Κ�� ��+fm2*��d���Vv=Š�0k��a(�ax�\��\��i��U¶�A}�1*��7�W<�E�S��1�r���t6\����?���_�ϗHk��\�~M�z����i�cd��H8�d���)@T�$�RX��
����ƽ���Y�G�cA��`�"�����G ��|��4����c�<Ι��6Y���H�+В����*��/�� ��ӄ �d� |#P��J؞0�	�c�$� C�-B��:0����IX'-���P�E���5��ȝR��;�#�Ch}oL9� ��=b���k+K���評D+c���J��P��X�eRin�D�N��i�=4��ϟk���~��G�do��O@m�˗������� w|cE3ZE<j2����8K�9]�7;r�ߐ�7�[��R'<�t�rU�IFb��u�Y�g���ԝ��>���<��NB�S���h��&�W�����`��0d���I?��y�ԚQ7cV�@�G �E28����:i���X+J(7��4�E�$h�a�C�O;������3���퐶,��X���cF��L_�����N��
��y4�ؤ�(ܒcS��3-zF��[��a[<�:��R�"��tp���0@,a
.2����0Ȼs�ĸ��/Ӟ�K`X����4�7�����@.'������v�F�c����.@���a)W�C�֡�6�Ul��]y@��÷"ko����@��]$3a]�DV� �@��J6I�=+���3��{��ss��\}�	��3����(O��x:����0k�R����$m�(q�[X��ǧ��ŏv�vC!�2��*B!�_I���=ċ.l����T�{�O.��
і�<��ޒ����x������P#�H'T�u���!c�":l�Z0y�Pq�ȫp-�<'4�,n��p�A2\l����h�K\���X2��f�v���_O!������a�s9$��T�H���?�/
����|��oT �
Û�~��</p̅�ߊ�yaq���	NC�ſ�4�c�~&�e�[�͉�2�=n2VK�HTL?�� �N+��c�|u0���� �d�i��u�⩈g�.N�?8aЇɢ�t�:����kUJ�pvI�^�>�wAO>���ƥ�h��MŶT$�wy�o�:9������r"��cLD�璚�٥�@���>@��D�- Jނ��	�?m��z[y�����m���,�]dtn�,W��L���i+�
���u��I�m��ҁ�<�o_�y�.-��;�-��������{�]{��~��
JE+��P�q�^!dI/vv��J��yI�~E<�*Z��"FA���Gi�'��֦���u!	5�Ǐb�����O�+鬁��t*��H`{��)�.����sKB�����TG�b�x�<�̠��&��&۲�Q�����n'� Y��Ϫӄw�6����q9\~Tj��}����nHz��/FO��no�ې7؏cL�#*ґ��7H<���S�M��\DǀU�.��h����%����%�w�ے6�MC^�I��U��-ˮU 8Y:{�Wp�uB��=N��3����RqX-w$^���<=�Qy��=�~5���-�������z.>8��Fs}�T���U��T��(����9h�7�)��e����g����i?G���ӄ&�@�M9<r�=�)��!y�:�m`]�ә��եsb���w�J��oh�!�
�^�� �oE;�qZ2,�p�a����K���>xB�J���HS��K��M"����=����.����̀˺�e�êx��.�!�Q�t=iQ�?��g C��^&�F}����6���57%��F�J�N�q<��Y����J�4�v�x�ՄU�(7�Y��E|8��OWd���AMu�=���u^�:+5%ƚU�
��j}n��ҹ&�T ;Z�;i<�r	�1p,�"�<ۼD��S�{`[������?F��,��!Y[x�X�n�[Cr^<��xaMa����'��	����>��gnG�He�H��2a"�hv����v�}�K k�e���ʓW*f$a��'b!�m?��m}vsa>J��P&�E��1���Pجd�:T��%`�Q2�v|�Z���iþd���C��ر��X9k���?��\�~�᚟i#q�*�%piX�i��E"S�C�HM�9�HgF'iJ�y�(h�IUf�ڝѓ�2��@"4�pΨok�U��#�e�f����s�H�B�s�a���B�1�{��5a0�������WIV��&,Q�.�%��X�Zh�7b�YiR|e�d�[�,�ԉ�_ٵ��ޘ�V��o\��&���J�z̢��aV�����FZlg��"H�V/�U@�zǹ�e��7��bm�"����������%]*��B%<��ǩ�_��r8�tb�������N�������I���+��7�0�|Ë�8��f|��="�B9eh4�p&��t�zN��s�!�򣅁7d2Q\Չ߮h�h��W�*B,h��K*�N]�BBb�t!c�=�~5����D͚�M��mi9���P�G
0�H��)	K�7�X]ƪe}؁��+��8e|�&��2W*��7r=/;L��V��M�g,/���!wB��w?9:"�Y���@��&�3>�'|��Z#>�D��]���|w��"�8dq��BGh�P�8oߏ����>��.{�o.�:��m�z�V�pW��|��E�j6�'I��d��L񦄐ю��<�xοɫ��/[�S�5u�o��?��Zڹ����z��#W�F.�&9�-���eF�\�ٶ+�\�ʠc�4�#�ڤ��l*ϱMYWi?j�afG��n����^x6�p�A�+M�{2�|T�����4$���V��]��Kd,bk����@�?�ee���e3o�c��띹4�=�~8�A��h���mF'�cCO��]����'�ķ�}�6"�������a�'����vG��k�*����()U��bJ-�Mb�=� 4�wc�裂���'���e���p.�?E �{@1���\�m�Զ��E��oij i��iē����ܺu�O��'������v��m":v�q�(~z�{�~�C<���J�!�.?�aϜ)�0��5%�g�^(�Z���q��ݪوi����U�v��y�f��Ma�	��QZ�T��U$��wu��~u����"$�����䱩ڂ��� ��-�6�%z�Ȧ���ń��5��e®�[���Tg��Z�z�w��s�9�
9��an3�غ��o(7\]T� L��.Tp�@��H��]�85��a������u݈�W����t�=3Tat�'��7g��-�6�V��TГV8�Wl-\!D/�Z�~�f��h$��@o���4W��a��`_,�VI��'��3�8�����F6ؙ
32>��
��KW�����*=5���]�|ݸ��n� m�C����\^L�������j�o	��?�o=\�؆Sҍڨ/��A2t���#������ᤎ��5�%9�!��v�~�:?�2���W�8�)f���M�8���]4%�U���;�3Y��*l�,��T�?�馭s�-o�i=((��&t�cf�	vM�/���t�B�M�
-�0��v9�v��ɩ�;�9���L@w��\ǒ2/�RC���7*g�֪��眹�:ao=��<���&zn��P�@.f�z�T�B1'@�#
j�/�	��d�p�c��l1]���U>S?Bd!1�z���U��{^�rpC���d.LKp�Iw)Q��.��L�1��ꍐ�.�Ih@����Ypr��A⁠8DJK��*��8l��n�K�a�O^J���4�)�}�l�7-�bg1�C��B��^9Nl���.���-�9�휃r��!�F�艍q�;��gM�hO!��^^zܽ[�?o�0'�������;/��!���������on"�_b9�V��5]��7�G{/��]j4=�\�ܾ�O�2�p�H
vo�+xS�sY�N//�XP�靁ZX)vK!�����mb7�΋�#93^z����>��#�'u\�t�ˀ��E�[�N��u��J*�BY����WD*���'���P�P�o{���l�8�����m	h"ľˉ��~�I���k�FR��3,޺�4W~���寛c7׈^->qG�5�ܵ��>	�{=�K|ztB�x�}�,t��{���j��p�m|%;m�����K-p�ؚ����<���
�%
.���E��iHYm ��ba%�h�\��{��|��S� �z�BH�8��h���:�+�؅�)������41�W�a^����-u}���-7�|���w��X���;���l�>��Q��>_��@�!�v4��a5wf�/��]%lpEz8	FלClU"dY�LN�~��?�%�B)�}�����F�a���@����lx.��z��¿�uk�[n�}/�f\G(�U7n'j@�6������Y��Ee\6���C���$��haf�P�-LN�_���%��yaK�7�������4�f��A �	�Ҏl���8@�zk�y۽I(�2Q��#H,�b�:(<�I���u��n�#J����x���sO�La�e�Z	����1Ɋ�!�@zO��  c��wSt� ��� �(Yѻ;�8�"W��)����ٽ��?���DIYf��)�,��0�̚��K��4B1�!iR��]�5�n&��x����s���M=���|��fP)�85z�`��k�jά&��,�.�̉v7�ū�$�6�ls�#��� ��ȧ��潂T?j|˺��V��qj�S�8{�M��EU9S*�ެ�U-)i~����C�jQ����|��n~M�t��E,@w���t�y���\<��P�D&����Ybq�]x&�_7pY�&�8���I�ޙ>�� Ս0{�I���pCr�Z.�<R�R��lVP��V��5:����k������ț�e?�%c��,��+;0H��ֺ�]�}�������NT㼙Z�T_p�	1O9o�1���
��6N��$���j� /���C���=�_F�]��<�)D���=�m*�Ӿg�j�����<��3�Np�t��S �#��#�� o�%�w<3�8�+c�a���s������)B-���ıX�@��ooln}�=-Ƣ�lL(r%|-O|��������+S���u��_�V)����x���8"+94����W)�2С��6}	Ф_��C�dA՘�CB$D���MUc �:V�l�)�kJp뻈�x�����G���_ ƻI��F
�¡������%+Ԯ)�󡅳�,U~v?Z�[�;�$�݋4��F�T��/ҢB�JRЈj	W�4���wU���ף����Z��������j�+QU��쌖�� ����� �%�}e/�Ux%�l��QE3�hVnW��EG��T��0	�ԗ��^|�?���A�]|ʸ����+E5�:	��;��i�4��Z�6=��*�>�BXf<!�_j����ŹG��2��y;� �3E�@<��S�S�$^&:�Z�'g��XR({X�wT�_�w�EI{VY~_�tʍ7��ʷ8��u�),$h��D�y-�`��<�ٛ��m�����%*0=�:g�圁7&��Ʃ��:I�l��"�VHf����0����C¸�}o$�� ������ܖ@�,�)m��+�9�a�NCf�-����X�����EMc@�>���@%���e}_q�RMD�/>'
��):���#q|��<��1gt�Z�XT�6jӝ+o�K < \�VB-��$�+�G5�c8MNƃ����:�P�ڻj��o!���! /[�(`����et�F x��Z�S��Ң'����b+_��`F���)n��/U�Kv�A����#���5%3�t1�̖���R��TDC���F�L��;f����v��Gy���^�L�+��5�!�N�B���s�+w�|P�����ܫ�3��r.|ᥤ�����I��"���۵�U�ꢫ�@�#�mA���������<ez�}\�6�5����ޥ�j��E;�5���qIxjR������㞓�����0���mY�daT��Z��V��b�Xm-��I��uY��-���[�Is��ף �S�Q��O��������������^;0L�J�¡J���"�������:]>E����lI���,�l��'��%�[u������={�<�"+�y����%��)i�/ڝT�9		�ƅ�p@3W��K8~~�)�����?25�,�����Z��A�ת�"PZ�u��)Z���L�X���}a�1�\| Ы�,J ��_[�H��OԱ�,���j��ɋ?��t��������"L4W�m��r��΁�R���D@��e����#С��oE_��j܈�P��	����E�yڱ)�ٍٰe�6�=%U�w��?�9j���-�x1�U�,[�g�-�a����e����s@J��y��:�0.ʵd�w|7B�H@=H,8F�:�*ޯ���	Ǚp��k=��) ���1�̅:�����7�s=��l<\����T�G[�d��gin�E����ٍ,*7�����5�!�k�I�&?ؖ��n���x�遇�M�ꤊ�T�R�Y�e��ych?B�
Z�P�璢���U�	��C �n�S�"��b듰d|�G���le�4����~�|�&kg:�ٺZ
.�����u�e��YL�	?wDrp'<h�	�;��~?�mέ�L�M�	��7(��w�X2۫Ff����A���"��@��j��6��w�́�b��\Q��l��M~�-ʳ��g#�_�8s�1,+����f>}+LV~��jqE���*����N+�jW#��7�}���]�5uX�����Y~&wn���%�S�>��ʘOr����;�&��~�T��1�E�R J߹�$�?^c���A�_%��������C��S�*�YB��=�5qv�8�B���_q�S�6q�2֠s΃�̯S��Ӣ��A��IW[�Y�K��H��.��u\M���1O��2��Qݥ��^K#h2%Qўs6����`=�/���q�Z�B�7��BI��2�#��[9�9�=��=
�Z�ZO��jbw ~l��l�ߋ��<�����Q���,!�G[4����4r��fy��2��(� &� �:��FꦃDJ��xa���Ų]���V>?߼ʔ���U��d����ѤV�s�]��t��*~�>��[{]늆�;�G�Qj�*a���C�C�-c(�=aY�`�2
�B���e�r���X/{m�*���go���c9c3?�)���}h�kߢ<)��c0�e$�ݒgeG���P%���r��מZ�/�pEWA��
��m�}ҭ�1�^I�ZM`x�u$���i�osP(���n�C�O5c�ca�KwnN�;���w�p@Qz#+2t�s��6�N�=<Ho�̇�b�#
�9� ;�Oa?��+}q�.P(�B9���-����ǧ��t���.�28��7�Q�Sx��#��\�"~�DPE���N�����Aϧ���#\��+h"V�:�j����p��/M�����}�����`����U�!w�.�����MV��y����B|=�R{G��{�ap)x�^�Yb �0�x�%iF̻O��ii!!z~�\��gP9��CG�s��m+y�M��5x���^&��%J�wizQ����ِ��ri�s.Rn�A7���s��d���H+S�Q�2�[&�*�b�4M;���31�U������g�]p��	���a����o��.�C͆���{���ʓ�eP�I`����� ʾ:§s7w����P�{1��/q�'X,*c���/���5�&��@�(�cf|���Ǽ8�n���.���խ�+��F2����>	t	�U��� 2��C��R�V��"]�<�zH�&s��c�x�(�0k	)���N�� �a�/�bVH�׈�+lw�(����/f���wV��rMU�E~�$�~�����Y��T�OW���0�
�f� ^����u�Q�9W*٢RVư�8e�(`���>���W�_��3pI�Q��bQ\?�?)R4�$cs${P��v0��"�X]l�v�����#qq��C�X�Ey�`�u�����{��m(��������K�?�2ղ�����]�i<~Q�v�77S�t�Q�3�2H����m�|�CB�h�|ј?��a�
�� jM��Mg��{�� ����K��C�(;ت�Kx�/���8�N	{�Oa<������qk:��٣�y���41R�]�k�MJ�:��9Xښ�%�R�5��T�ԟ��#~�}F@raO�X��XwɊ�aѿ9� w�i/�@�%'qe�H�2[E��}?f�e����P�n2ᩣn�1��ԑ1�ɉ�s�o/ט��|�a:�a�az5�P(C(�m\��z��B{��!I�L�I4�[6���[w:YF� >�D�!���k&��#E�גky���E\,�2Kn�����{�vzHE��K��k�?oL+��W"�΄Tdʬ�Ù�(O�8��=b�,��@zj7Zx�>1&0s��:�?�u��B�-����?�h5����.��Id�����W�FQ������C��kn���܍
�9_Ey���{�gq����b��Ǯ�����B�G�X��u��%{��"�J�0{�N>ɼ�PR=#�������d���ψ�%B�A�V����C�V�R�?# 0��D��w�s��s�M̵.�ey���@����-h�zCƴ��>[FL\g?���Q������L$n9ɯi#�O'4p�x��Z3�E���G�d��?I��-�k��2<U��!�m��`�sV���ӯ���.���aY>ۘ�9��
��W��4�R(�ή��=�ǁ r�b��#g��+���{�F�!I)9� P8�iu�!��61<7�Q�ɍ���FQ� `($���7�g���qU��!��ug�:D�����'���2�6:�k��Hb)08��/�Ч@;nr^{�?jMI��z.YA�3�4Pi���ۻ�?\��u_�ˈ��cڛ��\�ҙ�?W0w)ց��i��ݪ��I|V��V�;B�1h�IVW��!����� ���C�r&���\��l(�ã�/�db|j�-5� ��g�8��>A���Syt�K��=��I*R�vgصlZ��0���MCS*�G��!z�n�l]��JX�(Ϛ�<=l"�t��A�4��U��O(�Z���M����+j�龕;n�� $H�����pjGb*��{�(����>t�>ނ߼M'����蜦����k�qO���K��ԙ�n>������oO��䕜��A��V�$�dW�f��b���F&
y]V%O:��� ����-NaG�,e�=LD���/5�I��1N�Y���?.�N ������։��<B�N���g^�h�)�-��\�W�����^�L�(�ac-�奝!sC}���A��������w�x&_P�@�MZqt�+�'�r��rA'�ٜ��Ȟ�0ӣ���;,\L�`�n���kjF6���}XS�/����R��М��ع4��=M"���
Wb2��pϵ1R�^r-�Ԥ!��#����}����`���3_M�ɧGчQ�3�o9#��rL��q��SJ�%q������R�W�����S�O��$����Q|Z���3�X�go��4���Vh�jW
u����׭��9Mf��ib���Nz� 2��jɬ,iƥ���-I݊� �����]��|%��8�t���1~`F�M5k�v�"�����^6w�ft�I����-����q�ۥ�h@Cw+�M��a���7��ke-�H��q�܏��I&1�M�ݟ�>�jv����Vߒ�R��4HN}˒b��}�:�y����Nh�1�~B�J�ht�ށ3}��^�����=�K�<*�
9��7�@ހH�.(A^�������!����e=���?J�e3=�=�@/Q��z�%cYA�@aWqv�aj��o`�?��	_!X�J���	�ȅ���΂i���T�
a��u����Y���D�	�ȁ1�C��k�];RL�o��pFku������d�jf^�DW)k�`� ��j�"�I�,}��NB��V�˶���g"�Ѷ^A��8�z	�v���<mH)�75:6���{sѻ�͔\�6_A��J��'��ۦ7�xx�eŤf�#݋M�y�N?���H2��ܾNb�&Z�h�x4u��{����#��[�"���|�V���u��ls=�ꡍR���_
���Y�Zk�R����Arýy�8����C�h���LҤ?��-�+��䊘G�͵g;><�Ztx(�$+]�XB�4��N=x���]�	^ G���zM2��,a���jΓA��Ѵ�c�}�l	&��lTOe�UˑANzq�;���	��u�w��dt��t:{��Ͱy����mvki��C�U��(���o�լ��͔ɽ�$�e��_-Ͱ!k,���ଽDcH0a,�.\�dp���d�[�i=՛tw����ߤq�k�)�Q�����c��`TI����I6��=j������$֐|�ꔌ|*M��>�@9�)&�`7iN��.w���T�M��o#ʦ�����l��Ǚu^�1wވE��J���8���I5׮Lzg���F)Ii��nH_{�/�l$�wK�����aQT$'���qh��w��v�f�B�9@����������
�}�|v�UM~��9R�w�|����Edab��6ZK[Z��B�xϠ�f�?T�c[Sx,wE]q/�X����<���0�)�#a�`�:g�>�<�2)�4�3H�B`aR�"�lf�6vЯ<��'L�{,�ڨb�&��inP�)�z�Š8U?����5����>��i�X���ܧ,h�i�'�R��!_D���ҰB��/���súb^C���4ZNO��T�y�������\�7���a��e�<g��n5��k>G*�c���Y�4)l�"@J����#��Y=���m�S*`������`A)1&\��K3���<$��	�.i��t-a՞�Y
���f�@�y�^�1=�x��;^�w�ei�h'|y�yi(����}g��`+=V-H��?�!�UE���{-�ռN1����R��èbb�~��D��;>FB>n�AV�=~n����Y�X���N��~!Ģ�k%1�'
��L�7D��ټ֋3?��z����ly����w.��\�Px��Nm���Oю��y��}?���\�Wl�
�*	�&̴4MR���ͩ�.k���?�"�O��coў-.}��Nhe+(��4!���ґ������/����Qs�.Q����[2�X�#�`�ouHB�z�����[�T��l���p<{�'��Ɲ��`�-���{3.�>����A�J�~Q����:����L�D������
$�����IǏ	��ĥ�&>g�K�.�� �����hK"��a���/�M+,����Ǡe"u�L􈿆-vdim��Z�Є	e�K#�\�^3ٜa+�8n�^��~�
�����!�6��]�)�x�!L����m�Oa4��6X0�},��1邻���>�מ�/n��w���OG�Pт6A�r}��`�8K��C�/Lń �'.N�$�*wď]]u��5#2�RDx��]_
4���:�j���n�_=��f�U��hv1����id�]/.7%��F)?jr�#bч�}"���4��[���w$�ϛx��%��e���N�^5l�MU���1�(���; �=��S��<}���^f����6GF�4��e8�H��M��a��Z>B����K���r���mTs0*ٕ�R���So�v�E�Έ�mwv;o�c���5���q��|t�l�����dF����2��X�13Ǹ o�|��%�M>��a>M�ޚ�Q���("�L��\�P,����(�h\.K�'a#_|y����-��G������e�Ɏ�J��y���|B�r}>Eמ�=�g6�!&�hFr�"fۿ�U��r�Ʒ� �Q�6&��z���[`�/X�KY���yC�'�CHݟ2��%N�׎-��[�q���ױ̍�ӗ�XU��	Bu��=}3R#���Ó2�뵀I�6"��ޝޥK��f�k�4w�n�����-q��܅ɼ˹�5�y�J7FL�����&2݄&|P���S�c&��\���ZV����d��
��ք���f�J'��bX��JiGb��%\�S?b2���1�NŒ���v�<��ˤn��'�SB��@8m;Fn�9ǫa����**�Y1
�p�I���z�����������QG���2<�1 T`��n6$��(Iuݽ��'j�? ��mPx��c�����R��1ĸ��d���:��$��y�4�����hF���7��/"�J*��Pv1p�Kⷼ��O�0Se��B��Y�Oȿ��;\�/�6��D[ҋ�q� ��o���#w�(D�M� r�V��b-���G�e��r����Ϻ4���@�A�Dp� '�JgS4�!m(��m��F�J���d���qF�JG�)�8��m�~r;ܧ0��b�s�ϭ�����4�r��<�����L������=0���[�<'��&������t�����,(���wA��C�D)g�U�,I��P]�;���;�����yߋ̣/Wݏ�����2��N�7�^1�l+��h�h����N�����d��E�8����
~�W�Gs~&k����Hb����=�ZW伮>�Lo�����8��f�o�`1����ʑ^���N뼞�8��`T�9�d�M��Om$�����u�>A�ɒ&c�pC���J@x�"�@��Y��������=������*�O��7%qե��
�yF�ۣE8�V���{Q�-�.�Xo `. yi!S�p-�HU�g}� :0 3�J���yߟ�g\�|����<�cGV5� �'�uܴb�A�Sd44K<0�Cp ��<9Ȁ�2��t�Tɽ��S�\.������ۡ%�,@/��	�J�[��&x�~�N���L)č��H�O����� '\� �^��n��B���/�x��%L�x��)��|7{݀�����{%"iI'��GU��cNQV�ҽ����ҳ����t���e��$'��>��Y;zE��G��G!a��ӧV��1��eTf����eF�^�X)���/4��F��@z2� �j�gKT�#����{'��~�)�o��J��;Ҿ�`�̠�gD�U�<�[�Ĥ8}����:S�û�V��E&,�{����QU$�*a,�̽��8����-ɪ���Cq�o�:)���3qXn#Ǡnf��f�L�J9g�LS�	~����ȕ%<R��jd�R�]��t�?�%�������O˜�,�.pt��Z��2�/�"b�7��v�����7#���IW�
�c%���K`n��C� �%��L�� p.�"�w��ū^�։���U�
�c�_��-]v>�F�W��ex�:[��≴�h
�vD���(O�Hq�&�X��˵o�Snj�u�d��sa����~g�a�12����e�v�Nx�vBF���R!�Yx���C��;�I��[`�V>���N���?uo��q�̸�������
��eeᦺU�ADubT��;��(�D<���g��K06"�M�V�%K���� �v���?b��5e��A<��X���&�R��e���R�כz�w|X�B���1S��g��c$�ő+��$N���\8¤A��
���#({�qf�˱W�g$��2�'ƣ�L1ucyӻLd.b:ai�4�;�4��Kuf+4��Y��,*��At&���>j�B��6~_�H�@�ۉ?����h���BS\�Dj7�"W�(
a�Gw�yF�N��%~��j�
�~�Es<9��ۍy�(�F��B�u��U7�s��]z6K�����������8�_�,1�m�("�ɾ>I�`�l�T	>؞:���TI��-ClA簄U�Q��T]���^l���c�ow��C��^�μ�"X��v�b�*�2�~'��v.'E�iG�X���v���͵���Fa+��m\���y0��R*#���%��� �����О�m2,k f(��a�A�ɦ-r�ܥ�-���I�;��<c��1�=���S�~l|�^��g�-�Bb�0�]eM�/iF��O�)�ay&�:IU���i�^"�몰�E��-���<�E��\qRJZ$��z{����x{JN{��q1����/^g���:�����42y:ۘu�1�����!��ŒJ'<���&����>K����[w�����J�4��C�O�<���jr��m�v���� �d	��-@�S�y�TFY��Q�oV�Q����c�U�u�0�{`��P��k~`��P6i�	��[�	ì�+Q���Bm�td~���<��F{�GƦ0Wd�`����h`��M����l;)ջ�e���nP�1&-�*n.���y���L/���(jӚz�`�:A>�".�)�:?yl���o[6�??Q@K|WUB�n.���ӛ�&�r��z��_dkD���7����( N��8�??A�!E�
����`���i��b�T�F��9Fe4q��8�d��}���:����4�:���P��y�eh��l7�ⴍc���>���.�F��-ǡ���������Yv3�x�-}�і����o��b7�����<�fYa�?�����
O�I�^�ׄtc�U�"�#�#wD��C�B�P�I� �2P�̻\��G��{dl͌���9�q'j)X�p����;�٫��qr��<�,�Pp*�-���T����rD6�"8�(/c�k�吺rj��7-�1��<���O���L�ԯ(<���\^jA ɼZ��7Cc!c>�`_H�(�	M��3�n@�<��I�t=w��V��t3k�I����d��H�D���=@���;�wYŎ��1��������}�M)@�-%r�����-��֒>��iwM��>���~�I�K-.O���V��$���^?���y��3P]�y��g��p>�.��X�D��=�]%��J�bc���bk&0�Ӏ^'�J%�T�� �cܳ_=���_mBz�?8"\�%몜 �D7b|�����~�85��?�t�^�I";�5}`�XdCJ�>�\'�a欄�k���Q���mUv#�^&b�]�ȓn�G<��Vw��Q8Bn�C�j��G�m6d����׎U�@ۓy�X��E����n%�O�Yz��d�̻1�!Ĥh�QXjA<��wG誓ݵ�W	+p8>j��G�>N��`�hEi#;f"���.)��^SyG|I�|��,}�ʃ(�Zf��wHz�ۢ�D9�����]V4e��pp�U�Pۖ�T���[B�ցOs.j��� �}�ٻ��?�W`
��xШ�9	��<F���7^�C%��gu�ݝ�yX:S&Ά,ͣ�Z�#�	�����>���� e�io�b/L1�[��e>��q��p���H�W�����#F���볚{o��'�v���J0����'�q�S�U�n��݌���S5���`e�(��{%n��}-f��&�G_Y�$�VmӱS�ol&`��	q1 ګ$(H,U!�};f�<�-�p>��}P������iY���^<.�C�o�K�� o�&1�U�UkI�&��l(Uw�+tW��q�#��]������c��@�)0e�6t��{�"$�?.�T�I!-P� q�n�L.��ŷ{]�;NT�+�]��(S=�v�����(n�H,�4Aw�5�ㇳp�eї�j�s�Hw��������?��$�`�*��k�(ϊ�����_�=�"x��Û��wq������.������Va&.�B�׸����=�����Y=7ё��^���%�aS�I�kT�pV���
��E��S��cߗq�uU}�B��W!����`G��:�o��88���K��s���գ�jty5i�"�T',�f�	��&8Q�4m鬱��D^���O�m��鿟GG"`�*��y
����Sh�>mJ�Esʃ�&����I��z�ޡ�o�(��d�����8�����fO}�`���;�c �ז�[��b�͏��y��s�L�#rQBNUa���b�E�w���"E�@��u����;Ψ���{��P�G����^�ǕÓ��A��c5�֢��UW*rx?�8�KN=�&���9HK��s#�,9~]����B|��aV��K��I�=rgXH����|V*֏�����Y�2�*Y�o���#[vU�ٹ��$�q��F�M������-U�(3N���,gϭ�O5���M,������M��ظD��+�����['��C�2Tx����;�lG�A���U��]����9ܔ�v"��<1z_�u7-'�DGT(k@\`oܪ�Ɏ/���� F';j�*wa�l�R	��Q�߮����	���Ê�׺�+k��k�q0b^E_�u���$HĖ�7�H��\b8�Q�� 8,
�SЋ]�Sޏ'9;I��h�����<t����z^;��Γ���Ƭ�`N��KmзӛZ�B�J��\;���ΦXܙ��~tJF���c��|z��Q>�h3r�d��X=��ck�pWF�;��y�/É�`Be֟�^��1�C�9ʁsAO+���W�{�y�b����=�j�8��hc0ai{<��+��������`mV��nb�(_�<m������AX�{a�ňeoJƃ�5��At+k䞰�6�L}��mF[��	�'�@�R���ñ���O����|�t�ƲM�6��!�s+�]d���((�R��MQ�r[k"���>GY�Tb1RAJ�3�ϙg¡�^Ԯf��m��%��~�7�f\�4=Ǉ>ַ�3��^���6hpI�c@��sz	�����e����r�������7��u�� ~���¢Ume���,%W��}z��A+��.��q�B;�p�A��\��� Ң��'���>vu�S��Y�]�;w��G�X�y�A�9��Q>��+���N�	mU�	����p}Y�'�$*]%=�.�//e���J���>`8�rG\+b�]ӆe��)�KZȾ�L)�i��<Y߳�����ͶLe��\��ĻF���W4*?�O�`:�|_�j�n�Oݕ�}t7zY��B%,��9�$r*`AN+@�J��=�/�/��K�ڊ�ݸ�F���"��������q�=80e@�a.sN U��@�E|�V%�R�y�KtoDpV���5�ûS�bw(��/�7Ar��-S�-�( �a��x�f Ʌs�T�5	�:�e�j��U���N�1�[��B{GG����1{��b��Lbә��Q>[��^*hRט�j�__X��p�KoQV���L��䢇d�4�����IP�*O<��n�s?P�>��`/���*?@Կ�J�rȌ5tp$�"��d<�,oo���S����5Q�3'ۭd!Rq��B|�Ӓ�<�X����*ۂ�]���!8@ׁ��.߈5�Mp�W��iy��L�����$��>�?J+�+���3���	Ș��ࣳB*Q%3�vQ��{d+�{��Ջ�-#&r�A��`NMqg� ��Y��$z2�	E)_	q��2k���J�J�J�[~�Dm}�:k��1iw� ���<���=�+��s�SQ~��x���]�d2
��ǬU�{��z�GH���Yт1׎�&��=��q6���G	XB�hg$⡤u(�U.�D��W�,ed�B����T��;�Q�ed�ϝ�G�P1L!���҈-�5����*&���G޳��ks tA��ܼ2)��gg���gSpc�V��[���#e��'>��S}��Ey�V��p���'��H	�� J�s-s��������bL ��4��#X����i�N@΅$��p� �nyͫ�0�����ӧ����'���BY+�*;󝟨s�L^�W���0JȬB�Y�QdH�]�6bLBt�;�%�������*n0l������q��ٙ}V?B��a6�g��wmKL� ���d�h�7� �9����3�?~>�'"z��G�SJ���(Ը��-�,���� ��E�19+�5��.U=���)�o������H�z�SwK�_n�j�4m�Q�Gx��(���kWU�uy6���xz���~��Z��A <�Ҡ:��ɢP�d5��� �N����z)p�/�<`��X�,��f1DO�B�t��o��	�F� �I���`:9��'Y�=���b n����omc��y��q��c���,i�n9_��$��efik�CsKT�󛤬nqcf���C��pҾ#��n�9:U�[�n�_��%���ކY�����;�31����>�ф(Ļ�Du��C����[n)��c,>�@����	����~F(u�������fv�.�fG��fQ[����"��gP�`(�I�ɾ��C��H]�ȟ^�1��K�ʇ��2�>��߼'��dc��l}g�~�nh��Bږԝ�/�����O���K�0����;�p���9G+�EP&C���ɻ��ދD�����K��A�4�t�l�(����;���~ׅ����\Me��h����`F=u?�Q���Ra���o��Xh��qDݠ�mz8��1��&��Kv^ ���GHa���2���Wr�)�\��mh/�qK\+L�)��E�c��5B,����i]�>�DP��h[��LC� ��m�6����穬�G��9m^	��v�Ɏ2�B�Bc>O���i(w;�I���-J0r(���[����I0�������3� K��*.u9c��'�6�Q[a0	=��h���5:�5�����������a�5\E��WF���6M[���#V_8<�eo����8��Fe?#���SvJ��x��(1k�ȿ���AECbݗ���T�t���'wFc#+k��b����@����B&6p���_7Y@	C^z���l���c�! DG9���+n�#�B�g��Zp�aH����pIk�����+� $���~����>��4�6��"�+g�ѧ�l�ˇ�:K��,,xث�?�*gq�'E\�i��%�j���oƓ'�Wy���w�������c��h�M�9����!*���+�w��d��-9l��La� R��hS��>�����Oq�ϗ�i��Vv��w�@�������J��c?�"�Hi��ձ�ˈ3<թ%��J�m��),T�8&��[jiމ�H�oSF vx��&7�V u��U[b��O��РI���l���eU1��fyޠ�7�dQ�+m|�����{C�i�%��J�N��L:���3�����R�i��5�~�ݭ�����dOq��t�T`L(���	��e�!M>��������[����3=�f�.��X��R�w��֌�jR��wh��qMu/s��B@}5�k��
ɜkTU�}�B���B�_D�.]�q��`{N_��W+�?e(�PN�Yo9~�[Q򞬹A3{њXR|Tj��b�J��^�|��It;
T���l�`;�Z���,��ǽ���.�u������H�{rf��k��s���2��I��,Q���s��b���֤�� ��>(+z;����~bz>�,�)4e�>���P.�e�?���0�u�I���v���][��R*����3��$�}��Ncl&�JM!Β���u3�k�t�*x̓�lJj���{��0QVޠ�	�0�^�GԿI@߂:{�`s��N �t������q�-R{i!��C�}ߒ�x�#:d���p�GA���HY|��2�&�Y����9v>[:y<�_��;�q��P��؛3k$V�e:sbiŵvLf���Sz�m�P��E���(:6�Q>�@�:n�~�.�%����.e&
f�LZ,�T���3�/�|��M#-����$�Ų	-;.Y�3,�BD0TL��*L�`���G�P92��И';6�{�$�5sT���0zJ�I�eۊ���"�t���#�3Y���RA�0�����8���TN���@ �-b��Wu�GU_�
V�w�+�{Q�O9�#)��"�̢��IYe��@H��.�8~>T�Z�i�\����ⴗ�b��,p��_�A>�Ń�\l�TRf6�o_YE�zW������q���$!_A��o}�T2�&�X�
1�/��B6�Ty���L�k9�����7U��@���䟶�$_�DK��~�f��a�h&����XW�C�G�?Ͱ�;�h�wB��HL�g��颳-�˽���m��Jy)p�~(�[� �NC����Ch���f����ӡ&��w�GkD���Z5R�&|��6<x�3N2^���U�L�*��)�q�E��Y�!
�V`o�d�]�6�#8��Z�l
Q�;an�%����´�X��X��u�Pk�z�¡��\yP��	�y;��Q�~�}��v*ݻ�6~��B Ҏ\9<�Ṥ�����~]��Э��{����	�}��g�m�`ҳ���ښ�R��&��t�������)j�b�^w�g�*�o����Z���B�`k©�@�Y�{	�|+�Zƛ�������F�k���l�)#~(���e�!(Iw�w��#��ՑY{Z:�Y.L|&d*&!2�K-sG"*�4y�Ԩ�.���$$�r���ޓ	��Y5x�X���U<���P������D��eML0&Z��9�n��Y}di�:V����}7�ʆ�B`O�	{$?���������\J��/�Ż�&��*���R�ޜ��XV�����'�	i���%��)��'�Be�I�l	3�τţe�Q �A�G�$4ۡ�VMe��*ܢ�D%FIpMo׼�E���H�����P����:��G.���#bG�MȲ�H!��U��~�SK�3�I��RKm_| $&��9"�U�7��0&��W�NKO�w{� t��#������>�j��&����l��H�<q�b;/���(�����I�� �6� k�^��ް·,������>��*����7]���:>x�謨�W�i�-(lM~�������"����=IZ����8T���f^挽��'��_+I�����Q]���(МlŹ#��#�<(�8���੖��_�1M�iO 5� �(��kL�n�<�hee�o͙#�ǽ��8~,Rz��[΋�ݍ~���ls/ꍤ��?�"���drYC歏���V���bF
(�<���m��u��I÷e�w\�Ca3�D�RKn}Lݔ�u�ܕ�t�&��6(�yG���NQpH����ٷ���(�;�4MB�����e����G���l����{pg��y"@�vU�_���S����.b��q
����r�o��_�睯_��.�A~ғ�`��h*0��QX��sv�IѤ�Ms�ĭm�,�	Siu�rf[8gO^	�iq.ZJ�3Xړ�3&��f u��Cx?:�}2Z�RjAp9ڙ`�ފħe�H3wl�vu�E�vb^nF��3��j����m؞]��ʽ#��t]���m�-iE[l*�B��!~0�fȽW����L1����E��Jn_$B�L���iQ���x�)��!�}����ͻ҂n��������9C$��dg.}���!X���Q	���rP�E�M����-�g,n�ջ [��tM!� ��uw�=���ERxH�h/�E��|��uPLg��q��ŝ�G��됸�頀��,|?�?E����0�K��X'���ͻ�N�͐�b����VK.��J�;���Ӗ�,D���Oi�n���2Wqw
@⼎noX�hۑy����
����0���7�- ��&�rs�ଚA 5/ ��'Mk,��^��j{v�C|ߴmPl���jr�B�;�P3?S���,s��S�3:�|� �
A��1,?BS�X��K��܍��<����%
���c����s��?�Rv	wC��.lk�S]1��RV皼+��KM�������q��F���qH 6�n�!�±�����<)�J+��M�,+�6k z~Z�B³�ݤA(�f�|��K�Z{�����D;7��de�)$p���V&���~���a�7˧�������h<��=��[al��ܳ?2Zk��S0S���mP{{�y��ԝ<�c�i��Щ�����f�$��1nT�=^F��3�4>��+~9�3�� 6�ΘpV�S4�kF�_�����?��� �]+Tai�^{i�����%�-ߖ�P*���I���fz��#}~���U4���
y�O�<U�g۫p�x��Q*�ׂ�H��& ������Y�@��
�~�2�`D�GvC� �����"��"��8�]�y�=�Uw������E�54[��;,wː$�~;/�+�l�[ʷ!���l<�H����i�̊en�Һs?/^u7��R�T���C W�ˠ1Y�}�ދ˯�M↠��.����g�6����jQ+�/U�g��6̿sW,x��8��SZ��7Y�Ӂ����)��8��R\n�!�aQ���+sx�b�B�r����z�0<yD��#��mjz\d; �+�ǒ�j;*;�C1z�K��� ���m�V���ԩ��0�J�")��x�.~��*�5,�Q`��S�S�õ/�įK�݉@�qq����L��.:3�@K&�
Ҵk#Lr�5�5e�L���P�(���K3��.
���M�bX�7�5��N�_�nN������W	��"/�}�Q�kWdtNH���	���_�zNt֠1E��j��(SO!{Lņn�y�P�����>��[a��Sσ�2�+mw�:�' d�g6��yڣ�@ ^�$S(���<��-}�^!��g�.+���T�/���+#�&�@H��1M�P!��b���9�x�Z���j�h��/S��~�Ћ���;�B�\��kw:��{�e�/�Fu��Թ��494mR*pxPRF$���8l�9z��3۷�=,�{Z�&�[H���>�����[s,?�7��&{�Q��*��k�wrI�i�M\@�'j�.7r�حm����g��۴�K'���K��6�HЅ��O {���6��G�!��B-�BrT\N,������~�j2�s��#d�n�j��<-
���CDF}���A��,uR�L�^�57%�Ҭ��/����?*��]���Û�^*_�;>mX��:��-�:��(��U��[5՝	<E��m,L���WЃ ���,���NA��z�7Z�Х'�щ�����K�9�b+Q<3�p�i>��՜w��e������FX&�I`@��y�ڝ�cW޻Y��ƾw,
j�䯖��+�R�|g(�K��w��+� ���M���3`�}��r�l�b��@�/~��$�a{u����Ėnx�?��K27\_�����r�;��Hѫ���cꄭ]���C�t1�Z�H�N����΢�'z�V�E3^�[
�9��jd�|�-:��/��&��O������Ŏ&�Dp/�^(��>>+˯���.Ɖ�joR��z����|ך�MʒA�l�5�����e�-��Q޴@�xY��$�8r�( x،�cʝ����J�w� c p��!�-�S��
+vu����� 3r:��V#n�R%ȓP�`�'�AIգc1�f�U^�A�'�j���<`�Qf1�\�U�86�;�fqo�q��a���=�2�Y���n��f�0�&?��w`I�S��
륨�Y�ֿS�2�ڨ-�G���Pzxb���I.!�;p}:��MR�*r.�.͑sYVJ�%�����.�.�|:��'�TyfOܜ�;O\��4`�(<�sx�ہ$1{��=�q����Mz��ɷ("�%_+�v*x��B��i�S�c>o�' �I�S�����v���E`8��%a�4ת�_}��	?�7�V��-m5���=���f%�l�zm�\��Hy����aK��@�.tw�Xx{�M�o\���ΜRƩ�R�s�ʉ�7�����YX����N�.[4<��'�ݶ�Xhڎf�=�/�+��%����όA��1����4�����g�t���'D�>��4y�K����S�U���c��5m-O����85�V��ī����C�4H$����5 O|h�n]�S�O����Wr�ov<�L�0��{�r�7��y��3z�{d�Q���uhꚀ��|���`��6��1����M�IG��x�M��q.J٩W:i�=,�o�=/��K[��%H���t�{
�"����_)��~�}��Z$Ѡ��h�^����a�OhZ.B���]����ވi��;O��G� 32���y�(-i����kqG�4̀7/��2�n�5v0Ue�x1�,v~TH��"ǂ^��Ʒ�W�sg�lL:,�"V�|i�(��R\"񭉘��	�
r�xROB+]�XK͈[Ⱦ��<v+O:7��Q��h���O�-�Q�Ԉ������rdt}#��g_\\>��mp�f��*��G�ã�%���m���[w�޵ �����4c��g���z���e�=�%�4�v������*��9 �� F��֧�ء��ow&i:�~Ǵ?F;eY[�x�=���_�7)�S��o&�D�PX�jRyhCOGA���̯��D[�w�a���m�4��l��I^���d4.C$�5��ld*�g�xTS�R���l��_�m�yc1��J�7�%޶�;#=��n��fak�yh_�h��s���tgM�{�b�3�W`�;Y�-ړ!^5��*.�Z��9�����_�Zy�68��)]+����ѥasl�i�z)���Cb1m�����	K%�k*��2��"nJ��h���\u(�J��c�͉e��;�S�*���f7��e)(���@� ���N�ۧ�z�|Yu|�Yo��t���A�0g�2������ȼ��	�h�r3�Fo�~�j*��vn*"��%�Q����$C�9eN�Y��|�9���1�:Af��>�����lq�zOu[����D�ɉ��dU�+?I����v��Ԅ�b�%�Y��d���6?������ hFәV�-��RR,D�.�E@�n��$yG�u�7E�h߂�C�:�0Qt,\��K����V[߾n��^BmFs����d2����ЫZx΁]��f�X����/�H�������5�Q ���j�����,EkRE*Lp>zױk{�v�k˞�Sip���pb�1�LH3Sm��ȈvG���b�BU��4�2���<C��};�o�SOK�f#+⽉�S��`|��%�
�%����i��_+t��wA�9���E���d���L"��%�PhL0*����=����^�8M�@� ���m��X�	�����0T�%NP*��o%�_��N��V��v���H�pm,�i��<�8&�&Ƚn����eŰ��!˞1�T�4��ԯ�w�?WF9AJ�� �$����tɭ��EFG�Z��%�͑�^��7}�>}R!@,z����N!{���T)+�܆M����29�
C�l� ���%z%� a�ѿ����u8h� /3jv���וXR�?H�hu�j���fҏw��!�g^��%�.��WQ�o����Ԡ��8�-K�Z��0LB�u۬2�Q����O�������RXk��˰�K:yעbq�3�D,tt譕��:�ّz�����џ�Z�Ma,��=�uE˰��$pL`���Lr�cA@�ʹR�@i��<�����p��>�l����	5ʽ��{�_N
�A�%��:� �i�Al/��q�ɤ�GPXv��x�,��T���@wn�9
Ik�Y��˕���uO����_���>G)�5�4Úc�{~� �'A���bGF�y�����������o�Lh��֝��~l�H��6d�/RP��Pw�yD�:0�I�S��R���P��Ɛ���6}r���z��v�d���2��Lͷ0�cC���dS\`T#5�����x���I(D��Y�X����km?mƈ~��9a`�qt��C���K#���+�x�_]>�K]�=�0��2e�y_�q��c���3,��	<�߂�_E��lEt���+`���5$����N�����ɕ�~�H�I�7�#7���J��m@AY�=S�,�`��%	�GK��$f�]~�x�����b�"�����x�n�ﴇ���r����2Rg�^4�7���\
Fw^�!��Ҭ
��PT#�B�;�T����z[�YD}g�=�	j�lCx\�.��f�ȗ�J�w*��O�@>��n�x���+u�K�(�*,�2���c�o�%��/S�1������Jܗz�I���R��E׶1�謅=��w�d��-,�l�R�|��v�����R���;_��������jn��σ�p[��n�B8A���0�,�M8�.�x,3
�� �|sz+N�g0_���`�l��:�aW.w���_�z2"���@�3@W�/ ����_,D�?�ɞ
�KɛQ;�\�u��X´n�ֹ���e�dz��n��]��l���Pz��l*N:�"4q�)c�s�����׸X!�:������~E�
~NB�aA(PZ|)B���G��+�ٍfM�9&�M�| p�ϫ6��hO\���r����0e������DDՍ�|V���9�
pk9�(L<���d<c�|�u�P��X����9#�6a���*��4L 7�z���nG�lїEeϸE�������3���[�:9�^t����+;�L�x�-?+�՘����hbBi���Ի�AgiӋ
_�R4o�Ra���8��6i����W�L �H��;R�n�����f�o@F�.ҝ��0�$V�ʼ�tȀ�G�!�:K�FW:߳u�8ƴTC��T��yT?�gY�(�*����`�D�4h@[��ͬ�l�	]>�[灑zn2��iI�#x�I:i���`
v&{w��� rR��y��!I&���H.e�N�*׌L~�+d"�u��)���r
�)>:\�2�"�f-����&f��S<f����T�YQ�X���G�gԎצ�υ pFc��(�偸�/�xmpL��r�~5"���BL2�u�⸲�6d�E�]1��(�̠0Ʋ0�V�V%�dW��I8�K�u��)�+�Ϲs�[�(��kB�J���z� j�J��פv���Qq��YX��%/�Q5�u��99Uv������4�qQy�i��*7&ZBLH;������������K�ͽ�W�f����8�a�4=���f4��j�9��d>�� �c~ �d�kN}vu�P}�1#��]A�u���\���pn� �r�	z0o��m���+i�4��N�J��Uv�R^��=���:�Ȥ���I��9��q�� ���m����!풤<�6Y��֔ы�=�w6�ڲ��X6�~~�
���a(��r�����������(��c�q��3g��Y�Q'qb��Q�$��j��W��sꇴH�d����C�
�9N�L8�(k� �����1��>�Z�Qߎ�g/��FŹ��D��g
�Є^����v��ф��:
���u��ω����|wp��+�btyN%�P��C���Wa�����P�����E��T��m�N�m���!G��Kv��[+V0��C�u�t/����c�΋��>p�}l0B�sI�6���QD�M�o����9��~��|��P�Y$p��_p��h�0-��0#f��Q�� ��wa���yce*�aEa�1��S�_1��Z�Q��_^~Pˊ��J���FB�%����1j�|�=�%�!�����S'E.�T�\����5|�a
B>��%����6�q�䤽�Q��6�?���RdZb��{ŝ����:�3+yEֵk���Q���<We�8͕���'�+��Qu&.�8fr��I6�|�'z�����͚��� �j�^x;ɰ�Y�de^�eh�LU3��N�VH�!~�2�ZKRd�l�_9:�<1X�hǼp'A����z�#0����s���Y�sd�6O�YF�
�P��H�e�2I+=s6�A:|c.�+�y���#�:��&DȚ&GZ��>������ȇƒX�I��`�eH��Ѭy6�*��üm)�ݵ��EUe�Q���y�x���Q[������^K���nE�->�Y�Lfr������mo9*2�X���W��U�Su"�sx�����C@�֢��q�e���s�z��׋��W�e�yo�9�2'�{C��BUY� �]��a:�ɘ��D�#R<уwS����Ar��x�q:?��!��kZ���Y74>ڟ�9,���P"flr��=�D�i�4n���Pe�2������L�ߩnv��#��q�]���Hd3!�B��J�k�=1�n9�j�U"���_)�mAi{F���l��6#��(����;�M�+U%��x"U�݈#c�6j��5fAUlNdW�]�N [T��e�K{�)Rݩ�g^��Wb.�|��x����<�l��N�/A?Q������q]��$��L���4��M��)iB!�];��|����|.���l��JL�htq]�4�-�lw�_����V�T��LS�H��0�F �bc���supw�޻g��2���V��GE��.���c�t�O@�9��)ޢ�Bp5F��GHV�	�F�dHv��q!i���M����X��1�Հ-�!���bg�WG�t4RB�cfv�sG�,��n�Z��ZM}u(Q,��U�6�����?g�$ll8x��e��il��J��|�#J\��G=�i1�'9�[��O�R�K�/%�2ԝ)
�s�~�<i�2�e؈Vl5�Kpq�w�pA��@���L玓���	�)R	�?�X����Ɣ>b��K-d
��%fyu�@&��J]����SP��Ѵ��sT�3�,=��������3��δ�TW��e���W�	d��^�E��g>߼Z����w"o8`�p샨íǝ�T �Q�S��q����cD�A�5{j�}�+m��)��n0q5(�!����\=0A�/�}��Ց���#8ymM�[�GPqc����vDT(M���9�6��-���h��;+).b�v�0r�5CM�Z;]�]�<u�c�1�y���;)&�:ʐHTr��L�5��`bi(���c$g��3EWj��Q��v!�D��s�H.���!I��[���0����W�u���d'�D���E�W�E��^#2�4!zO����C�$(���o�1�N�a	�q��#c4�5qi���Tu�A�%��[���Q�R��p�����)��!L�>
����=��抢�[���vֱ�9�VT]I��Ȕ2�]�@v'�DA������~>L��V;���ڜ�3[MB�s�"u������]��49B�rP�(��/uP��e��K��IO6�c���Y�93�=�f�3ܳ�=���eeHb4H�^܂��dm1��+F�D�����,t�N��"`ח57o\�v9�]b8�찇�����r�]���i�z�S�dY0�%N$ s?\`{%_At�i?�qc��'e�k4_h��Pc\���R�e�CA�1�_�q�ڻ��,x��S%�k޵�"�V����6�!��fW��x�����mK�~�:s=��-��L����PkDZmϞ���0OQ�9Y���b2��d?)������N6����j� 1{���n���x���bh���율�H���Q��6�>:-f �����s����橢�G��<KxS�(c5��6^-S�9p�7z���C�Ʃ��)��Ux��	~g	�1xT^'(&�EtqC)Õ���o�M��f��L�2hy�ۢ�x.b.9��|����]��\�[��e�j�������F����	)��^�/�h��J�'�7T�Θ���z�Z.����Z:���t��c�i��/=~��U"A����d�^��|OW/l��L����/�ۖ�f��H���Su�%�qJL����D��G�b������4��_ Z����\;D%��)h)<A�{���p/@Aܙ��&���14Q �=_�1]�I���%�p�d
����F����2=w��e{(^-!������ښ�ޤv�P<r�ҿƷ�Y��̖A�FȺ1��V���R�P�Ԟ�*@�'S��VߛuHng/�2~��,q� ����S	�V0�p�Ֆ��Pvau�����ɀ#0�G�^�y����2(���1;,%T�߂P��� `�*�<RD�CRG� ���oP�]5�n����{�ʃbS������?gMv�'(GH��Ι��w�6Avpih`iIC��p�z��2� ޓI|�`��"���U�UDE�,[�%�Ovn97<I�11'��T_ǟ�Hx��УC7�^�+-�w�A�5M=*ް6~�Գeߏ��p��YZ�8�)��tg����7������&��R,���6�^-����s��rP<�a�G�q��؝-����+�Jq�J@����J���La����R����e�P�ٓ�p�Z�����@9���dT&��{i��E��
Ѽ�n����/���۩[
ۚ�p�#��ӎ����g'�g�5��ML������<�c�ԂhÕ���B
��IN��Dm7��*2�Y�q����i�_m�.(�� /��4�|�3�/��gC#X�i���͑������H'��|/���	�� p��R�� ߓ�P��Z�઻��jQY/F��qv�ɤ�K��I�p�!5԰�/��{��\���H�90�@�w��6,�_�.!
M�'2m͵Y�6��M�hD�
�Ϋrh�_��(;���ߑ����Ҏn��o���ΒŊ��~�	�>�Q���2�G��$>�9�
_'��"z�����c+��I\���^�r;�-pa9��_F�4��V�q��!�g}�B7�;���1rK�/ �.o������N*������H�]�+�6�oؽ(r�3�Q�M�t6�\�gV#��5��9�F��w�~u3G��T��ob/}�>!m.й<h@�z�Oz����^N?.G��L�O3(����hY,kQ%L������3YؗWt�,�)�������^4�ϴ�T'yf|��i��s�U��-P�u�C��՞��I�������	{^J�7�10�_��D���֝դ�dv��뷠8�Ro6뺐���<��7�O�P�,�`1��f��G��6�6��T���Z��y�|�|�f���?ձ+�F·?�vV��a5����D'K=P;Ou��t��v{(�Z&*@.lՆ���d/�}qs%M���/AW,�c=��ߠ��l<;���	89�.N�ޥp�z{X-U����)XY�*La�D,D]���-n��,�F���6b��L����\S��z}-���Y�G�i�1{�O���Y�3�26���V,��T�����f��+ز�[���5��ts休�g\-6 d.롰����( HU'�����0_����3�x#�Lg��ѢL��z�%�41܌t��~��=�_��D�)�a�P�YHG�vD�W;��t�^iD�V�f�d�p=~Ӑ$>и��џ���r�d:���_��SI:)W¡���x��@���:{6g��V�Nv�^y�`�� ��!��zx�k`�� l(��`�է�Yd��9����Y{Ȝ��d��/
��I���^'�3��I(@X����dT�牖�-7�=�jq����@���7������u)�3��|�F˱�����^�������"4ט��Qc�9
E�8J^
�n�G+�*�͕�	l����h�#��]��~2�H�C�2�S) HOl����Hr+P�0Ųu�;0Q��0����������<~��.R�ېK���W���G�l�����o`��91k����j̵�����{�X�2�}6`q��K�dH�����Vs�@�<Ax�9�/_K�����/�};�`s�����P�tե߲2�g�/�P��چ*l�}/π��0jf��6ɿ)ƹ��j��B�Ww���U;h5T[Ufjl�����"�fD�p�Ӌ�[�4��mJ��[�Sc��p,�p�/���Yy�~j#�D��9,��<m�z�%�|كr�=�ۼ�>$^�'f'/]���b��\�f0�&
�CMqtp��I$���>�8���$	�k�xq7�g�B��E���ϫ�6X���5[�%C9'ta��>�U��n����~%ɷcv�Fb7���
I�@���=�ӵL�ւ�hz<>�f{�ޡa�Xk�[�ʼ�l{io�}�s�jNg���B�h9����(��g ��S<�4�V�Hu�G�y�S���5K�� �4x�!���<˔���)���p *��dkRS�9u�،`~C�:�e��y�GV���5HC�7oh;�TB$�?�6N�I1:�%!7��Ϡ��K� pn3��B�#o�!��s*]��)M�t��R+�Ӈ{A��4x	 vjc'���:ݻQ��"���A�D�շ�k�c�A�(�Vf�	�֍v���m����r�`������-(��2��Y���0��Ly��Ǵ���j��4��vD��#�.P����Lh:�=��|���d=��/��Z+�pU����0�8�A���?��`���8�b,�N柩pؿ>M7�ǰQ �b�6�:b�`�u�k!��U�0�Q�6��b�6��l�H!]r����J���`��5X'�r���ަ۫�M˥u:��LDQ�ƌ��$�#��Pա�c��C]Be��("��\�$������E6:�r�&4�:M�W{��dY����_!��e�"q�[ .��1�6�T=ҳ4�ޮ��c�x�K�������t��'�V�;C��xݽ=�.<��aòQ�X�3\YBx��
ճ/�.���f�̆B���IS�R���7��.����a�4E��,�p�yתӖ��(��i��+�VL��&��&VK�&q�Hg渜~�K����7���f�z��,`�7"ST=X ��4P�KTv:�p(�̕�j�UwM�IӢ���p1�*O ��]�oJa.�mUh����RP�l=����3�H�/�Wb_}
/��7�	�����e0��Z�u��J���3�{�4SǅKh;9��I��7p������wh��ox��/�	��|�'����:��b�h/�U�"�#�����2�=t˸5��{��4�����g/��2�F�Z����;V�A</�$A_w]�C ��c 4�{�=���e=��n6zL��?hV�	��A���f0�E�}'٥u�5�����/����X���F@������"���9�ct	#��'������̪�/�5���Ƴ蒅�r�v(��<T
(zIehKn����ȧ��~R���
�H.�C��ú؝��%.�QC�v��>��j1p�W�z���72�vJ�Э/�+��ݯ{H��^m&�1�����#��No��|!�B,-�Mԡ����N����AIǟ+R����9�R��\�k�$���d���6������&��o��T#����M�p�,\�*��g��y���>���cJ���6(Cj=(y^.O��z`=�7w�[=P����D�k��� 5W�	<�g�K���;�J�F�3K�E�w�6\o�fm�Pd!�xX�7<��ӫ0��������gT����K�.U�Na��f��ʨ�t�����D�����ϐ���������dݐ�#�g� ��'H)�S�c�G��-���ͣ_�ٵ�.�nw�~!'�2�vp$�&f� �3�L����*�cm�w�(G�#�fnJz�\=f�O.�R�;Cj�;��"z�=>��:�F��c,�{��x;���aBW§����x�%�r*�vާ��pxf�iW];�> ݪ��G$��Y���Mo�8'5|a�� �,_���?��*��~i����0�H[N�7Rl�C�le,.E^�J�)|����K)A+���^��4��?)��f<;yK,na�-�O��0A��[6:�"J@��G��44$��p��D)Ow��)�b�K"��)/1�#�sT%'ʂ�{���Vy��9��5I���^d�>v�s��f�C��RibX�굞������+~��x��L�^��2�Hh}9��7	{l̆~��-»���3�տQ,\Wy�!�q���%)ȧJn��B��i�5y��C%I
j����H�|�"��?�����c�MR�#!!(c�����\����I덟��<+�J��l�JE]�� 39�;B��~o�S��\�!GB������������<�a3�7rD�)P���^�2��#��1������8ŵ=��[&���Q`���X;�����VE����NUxT�Цr]j��aQ�Q+�&�s��)�9X�O���������W�R��H��X2Y��=@T�gw-�?�G�7�O:��xA����UxYPs��H���H�
�a�+���r�|�](A���-�����<��+(H	cE���38ʤ�,$È�5��0��������Ї�ר���>�����*(w��>.V���S��8\�રS�يj�HIc��Q��;D�� �-�m9�����Q��%�A�8�֭6�u�&fg�<�gqQ�����=��0幯�)�����MC��{w�	�B�:��Z�P��ә���UN�A�G6�����>�:�k�[�"
�{�qR���n�aZD�;k�� ͝Ƕԩ4��@��t�|,Y��� ���٦IUI�F���l���#�8]'�w���@&��@������c�R��N�9�ܒ�O�F9��L~�Y�hX�y�$�El��S��%���P����b���9��5�M8�R�7 ή��gR��e�a��vO_��>@z�"?trtx=�"��C�q�{a���c�:�
�F;�UC�d��H���w�{�}�Q^��.;�Ǎ�}fߐ4����k�]����[G�:f�Q{������`�9���z�dj/��&Qt�h��kJ�@��Abo_��A��j��nLҢ����ŗ�^�騭�I�Ĥ(@���h�X����LgH�1� "�j���$�~���.���$�9Az� �J��󕁻6�6 ��ֲ���xj�72.��?�B��I�s_�EE����V��9�{����[#�B�ʜ�	�Pux|�W����!am�xT�?����9 �2��ֹPY?���p�C��{g�~���,<#8� �rWbţ,�Nvaw-�9��,��P�L����h���jʙB�id��lv��}&Ig�H�X��ο�+̫$	b�3���j��������c�k��QR���k��̲ͅ8-�1O�fWwJ@�E�v��e�Z<hHͿtBu�_ [.g���Zl��� P�Ζ�xc��z�\ۈ�H��.t�Y��k� F�?���x���j[2 �)E���t�B4���%$�,m<H?h{
 ?A*~2�Xh��N�ď�[��l#~kU���8��7:�����K����*��i���������F�LLq�ƦI�k����6 Q���y��"}�Y���#悿!e;Vg����VMmu!�=c�0Iį�P�l~�����
A�=��jȟ@gC�!ϯuu7��h#$Ł��#�Z(ZhU�9�������2�s�ѩ��)Ɵ�?�h��l\ގ���2�_���#]9Y8����d>�Y����z8s����IO�̢[�Åp�*�4�u\�Κ�?�qj3��a��ʑ��Hʼ�#�O�[�h&��4���io�S>�v��.�T���X�D���r߼����,0b��{���|0��7��֐�-g��S��9GC�{0��v���/٭4:.J�x�X������2�wX5��j_{��+bgvVƑ�k��Zº�o�K,$�TQYR�k�kt�%��=)�`ML�ٯG�����E���� �=��Ε���� *��]b܄��U����c��{x���Q[�;_]��̘JW����W�Q�_�~��dv�~��27h�x�2��4O����l�����T���3��j��m�Y�9L���\<������4&���)�	=���	:s̾�*�u�q0�®�Hf��5�p|�]�?�z���O��-���n����g;�D�����Z1^xV��cΪ���tl�8�Ɣ���&%��T|U@���L�P�2��5�.��8�q�����
\�#)S�L�sNx4��6�jb&�s���#7��N�U���!��s�0�3�P Ԝ��k"f'<-��d�8/ЅsJ���102�m���Y�g���Wy�'U��̎ \G�sYV��^_�c���Ѕ+��Z��Ͳ�m|S��b3~E��5Ɛ�H�
�n)ű���ۍxt�\xL����T0$�f ?��-\F���Ӕq��2_�3����f�B��6���`�R���\�\cҏ����0*�M�ټ�|c��n��U����tRL���n��wa�h4��2���Wzhr�@gj��bQ�[�H�1>�Q�D��L�����p���ř���Ea�>�'�t��Ʋ6yA��ZݖW0�4�n�&�KPC_k������y�q�˂�u��%>��,�O�<tZ1c���h��Z��y}����E�Iy{�b�Xi�O�������zz<�nc�U#C
UҞ�k;�Mz{F�]��X�D�L���+KÎ��8�(>�xuD`K�2Tl�4o�Y7[�[,��k��x����m�:���I߈�1Q��0��1�A�]4y,c,��l~|�Vf�y
r'�O�\Mw��TbYs,;b!����8��v^!T�!fy�.�G��2Mgh8e��|�?R�����~ܠ����?q�McgPg
�"�> �ſ���ak�zM[�*�V�XBJe���?�ʁ;4�E�/���&P������B2��@�ۓ~q���My��m��d����0����CW�O�Ǯ���Qۆq�L�~�A���.�O�i\v-J�w�=�V 'a�1�0&F�}��I��2���E�L�0�ϒ\:���,5q���\��Q��
_��}�"F���L|��q�Sa�Z�$��1lX8�h.�<'��T�ۍ@mI���;��4��5IM2{}t��W�p��B���j*M�n[�}�f]F��7x���^��~C��Emt�wH�Û�q�@����=S��$�P:Ӆ�5N�®|+i��$7WLS��P�҆�)����K����F4���O u�.Oьcĳ#��G)z�|~��B��dÅ���;�~�Ԯ+�`�����,�����Vr���f�^�<�ݺ]K8l؊��N,愺�V�.�r?tY&�gL���'������Bp���g�c�T�T��l+��p(�CF����M��m���F -��vf�`e����j���b�W��)f����u�,|m��*W 展����қ\�8Z ��UV�����nj������9J��V�o�b��R����	x��c�_��`�e^&Mh>l! _�\������y
Q@���篳��,5R�mH�&��e}h��aR��w)�cx�B[�;�����_)8₦1��O#^����̈́�H0��Vd2�u�'
Wu��x��6����������N�1��)?A�|��u+�Ҭ��.)�\��	Jޜ��j�`��#��Ѧu�p��f���j�ҵ�Qbݯ.��n���qRJ�p�F6���XW.cܵ����aqu\c�R�+x�!piϞ��i�턇�D��8
Q�#�ήˑ�12ـIQ�b�X�Eڮ�; hh౷��< ��w�d��q�'M��b�x��Be������u��C88��:��<�z��G<��`uc����;��X�9�g
)���-�=�b��BMW�gb�1lq`����؂��X;��yU���HU��4e�gRVi���,�b�b�x����g�K�4�Z,�S�n�mK����y���UP�鿔�;S.�3ݰ8F�US��o�Å����i�Z�G֑�d�K����;�Q�I��n~JV,V���d�0��.T��Z�Vl<���nr�_6
1�Ǽ�C��g�OX �d�8=��W����޺��䢵 �z���6n7�5C���$��z�>0ʷ�׉��~]�-��g�5�|���i�
#�g��w�-�]�F@�d��,�\�R���5��\j9-��C�m������j����c���l���:)�&�m>�F�3u�wY�C�����YL��U����!{�=C�-�7�&9�iҗw�����uO<��0|y�;�+�,��NAL<?��*�t�̭��+��v��������JLP!Z�Z�A��Ϩ��:�&S=��Iڨ�����Q�£�!aDq?��O8j_���T��0�����h1{��p<T(~qI��C�9o=���vպ�!-m��ڨ S�8Ѕ����a6 &6�{��&�l'?m�Щ{ˋPM�@�!.t�\	]�c�EA��l�����W�	����P�E�8�����5^��DKY ������y�[f����>dP�7w�<���@e��J|OV�me�<�/�O�#TɈĢ�C�%K����:B�I�bO�J���-1�����S�:gS��FF��@��7H���b�$�X�1����L�8��f-�������} K؀�#F�x�b��\�꒲ c.�Y`h�
���Z5Ƽ��9��v�WTg�*M�#Uҳ^ʠC:��_y����z
�լ3fǚ����g�w��>-NR}AMIU-���<�l�a�0���,|T{Z��``Hs�O�a�J�ɚ��Y�xdP8��j��E=����R<�m��Mm�2���҇SV�B�������>�R�iPi^a#m$��U��2��d����XÎ�X>B���ԋXhS�>��`��{R�{�(�Ja����f%^$:���%��f)T�R���h�nց��ug38�;Q�3�h]����I9�g�g�ݕ���E���,�
�`��;ޑ|��%F�̣C�+�Ԙ��v��ɧ�"��v��8_�Ӈ�����}�R~����a��A�~��(��O޴�P�'�K���E)�*�X�\�~1��U�DR.3ѳV����'kMeք��I$��+�?	�VI��J�ަ���
��I[��MIYAk���3��ְʺ�W=�iN�q��U�u�z�3�i8����;?1�
�O��x����<� �\�E#�T��B�����x̷h�[^e��wj�u��-�[��j;��L-Hjh{��F����5	pB�,�I�:�BH92���;����Xu֡�G�7�Nx�����|���1f��b���ҷ������6��LF��љ+L��e��e������VH����>�J�ܘ����|�KX��l�Je�
bg�����+|�iR�g���8R<wV����_R��<�>����ق����N�=4dW�FXW:!��g7Ig����+ë~LE<�'�|�)����$��M�/Ne�9�0ݵ�D����N|H����d�t�<؞`~�oW pu�r��m����3|=hI�����$-F�>4��L֜c�fATx2�X����:���:�-60y��؆ָ��-"B����P���
�K�$�B?ؽ����@�Z⵴(tIb�3��b3A0�R:��!���4A��"n�G/�Њ'��>����`䭵m�@�0z�I�B�����|j^7��³^�a5R9�?W|ǂ�pCD�i�ד.wG1��#��Ug���T������?GJ�a�8��A'�����eW�v	���HU����0�Z�X噳%1����׏
��gU��ẻ��Ž,:�sB��f_���f&����MÃ[�h�B���~*��o�m�z~���{�A��7�� 1{�U��PlK���$pީ�n.J�+r_�JSo�;@Rs.�M����F�\�+f)G�6�NH��#�E;�k�oc�P,���4ڜ�[�2*��T��5=�`f#�x���S�� ��w���G24E��y3ܶ�13;_:n�?&�|v�x0���\E��5�qQt��������q{$)�c�e�켅�(�V�]�0��r^!�㢿�g����@o��sH���C5jj�%��T6��ςH��q���xlNi�Z�����;U̵����1xs�o���c��-Ȇ�c�E jI����i��Oj��#I4���e�ѣ7K�b�.g{�&�}��@K%�@0����?�{L��w{�p�:WH�y�z�Ir4�E�E���G�r�6�ޔ�]Xt�Vߍh��IR��\����GO�}͋�����cl�P���kY.A��\`F��-���u�/j��A�d���c.�Ӵ@.�c�6�"=�����W<}�+D`u]��YN�m��y�\hZ�vX���ƠQ��	By����V0�*�0ߕ�x�\�Il���p�P�G;�Sjl%�[�&�΁D�#6ɍ��L�^��ūS��v�E��E�'4�;�[�M3y_���,�k���!pM$�2�L�<�ɏ�RF����,^MbC��CD�O"�"�y�WԸ�Z����j�"��(�\��zuCB��7���� Nt$�dq�ֵ	xV��Fu���"�;�	SJǣ(��N��˹Z��!J���[���o���&�+�i��t\�J5C� �s��ف�0����m�;����CN�\����x��Ff�v�<>����{���Wɏ	K�I"��NvT�+��D�a�P��z�Ả�P���F�����zDx��?�֖���q5�l�Fv��5�ͽ��0nH5SL��%����,�H/��mpY%�½w�b������g�9y]���qе�zǴk�Ŧ@���0M��')���QxB>�vf��8<��p����\cP�p��mug��d(��Cˬp?��y�t���⸲�o?�t���G��st����Bs��V��Ɔ�p��������wq�l:_4�r��P��đ��wR���G閦Ltj��T�M�0R�~	�<#��Cs��'[�h�8_�N�:v1E�6lL��7Qt� �	W:elt!����p*t<���5	g�z$3����\��a�F�a��?szS��*?�����5ҔA����V��(�|Y�p�?�I�O�=��e5���St+�d� �pS���*Խ����>���+'P[~�N�]��Ҝ�����������7*��X��� m	�mʋs�Xi^e���4�e9�b8���y�\x^�Z�@��A"�����o��^y��&��c�$Kfb��:��M�Y�f5<3��Ɋ�m��eEPBy�G��_y�����5�{�xmn�1�d\��ue�P/���,��b��4Q�
�=�"Yݐ"'
$�#�L����3�ې'�*�;9�>�r�� ت��~8:+��G*��qf�~k(i��N'(��?@���J�ִ`L�C�͇o5�5��3nCJ�~Ls^������~LO�n�o�?ֽ�����
�V�:��3���XfE|�K�JB�y�.F����{�T�Ā4�p�\[Q�4[K(:R
wd�	�F��{Ae��)��n)z���5#R�����\���0[l1=�cH��I�
��F2'TRm�!^ڂ v�.�ŋ�@~����Hh��h����A��ȋG�{a�}����t���I��j6� �*��"ځQs��s���	����I�9�1X=0��Y�6Ki�h��x*��|��5����Q�$�xb���t���7��`�+>B f=!��p���Mm���,��!F[��3q�>�˨ǖt�B��XS`�@täC�E��(�~2�U�N�a64-���io#�$(o�r�� 5}�榮rǵE�04�P�7ԣS뜶F��R���v�m�خ�_���/̺����.%�����W�XH��*����)� �_����y��[��J]Wْ<��m��<3���(�@3�2h]� H]n��+�O���X�x2�nR�h���U������Fȣ�ZN����ʜp7������
>�������5���ś�#�ϫ%&�zaJ�$W�!��c೅��X���b��R�f42�'����b��ٟ۝���+�jb�H�dS�ę7j��A !W x�H�&�FY�
�Nv�:%��@�@>)*rI�)nر���ǂU�F~Ccs� uU�eo�/z�&9�Go>���J�w�۶CΈ��]93E�`�)���8&)�=�Eͨ_4��]��_�VیH�`�+S��M��A�ط.;��Ӏg@ʥ���?�ؒ$Ѽl�>��K�O=����U��H#G5�����3#��>P�����=�'�Q萸��1<V��)o䆄� ==�>����[�Ӄk��J���2���| t�
 �]3y��h�����#�[�IT�)���8^c7�sc'�$3_b*/:��'�S�(#�rv����3�;8��$��E�q�m[ ܰNC5L�X�	�n}2�!���'�< ���^	!�[YL}����؊%qҐ�X�~��l���c�T$�=H�}ӻ�*+]ɝ,w����W�5��:^��JL�N�ɪ�#+0?�֑J(.�K�D�۔�����zHέF�<���lt�Ar��5)�]#c��Q��)Ppֺ+<�'Y5��z�����d݄�%b����iE{�jO�fH@=����j��2 *�1��|�f6��g iq�AMz�����ל��G��B��P�yv��G�
��(V�?9�8�VXJ&�l����3���ZŁ���D��:[�5IeRf�+��^����v����/�e|�/g[�� �`��囥��<�YZ���r!%�n\f*jɈ���Jсt��̗�+<ƴ("�\��i�ˀ��.���� ��@�Yn>�x(�[|�l�}Y������7������P��&���{Ⴢ�{��5�3f�ԑ�ߟP�n�k���<�om��L�Ŗ(�!B��/X��9p��.�;@�gK{��W���C��x��b�ޓ���n�k5�?���eRY����|�V�[�o���8����儥7�,�u��,�4�\��0��G��|���������n�<�����J��ߙ��r��iQ��Jh���c�������6��{�;}QK[���	`�-����/�n<N.� �濳ɘ�d��Q���d@To][��mĚv�r������!�"<*����)\���Nl����=K.+D+.J��k�A�DRM�4Mv�f��ǟlA�4g�ž��/(ό^�N�o8�^��bXY��,@��(�Û���ʧ8���<��o+�����;dy�������qD�m�BR,[�}����!yͺ�b�O1�4bɱ�[B�bx��;���+T3v�Q�W��O��0©>+�;��^9l��E$�J��� ���Y�Ծ����d��� ~'�A̤�}1v�xS�;��b��:��[�)8�A������s5\o$Ӗg(ǵ�f��9X��]�r�Õӂ���vE$�E־R��N��ٸU��vJy�
Z�愤�*!#���}�$j����nB�E�M���X�`�A�2H�c{���q`��������t���S�xN2O>!)ŅF�X�{��!C+U�u���
��y��Nig�M����L�Qq(^�.����WO/9�ݛ���)i�0C��
$����,��A4m�j�����y&ď>mq��,E1 �aTc^t���^觰�+���j�19e�����x�d�reC�R��֟�'&.��1w�����4����ώHҕ�10�T�y��e;g`�~�&�P�};���|@�;�']*sه�l|?�V^,�B%�\�/o��:b#��IUR�(��l����e�6��xt��\��t'�r< �P��8�D{5u�J�|;h)���6���G�S�b9{����V.�%��k�4t:Q��I�<a�A�R[5�*x/T2�C�j�^wwt�28N%� e��3w�f�c=�@ �<ۨ�?�m�"�6�d �2�ż��!9���B�xyo�u�2E���!��j�w#�䤟-�ݱ��n(��N�ڨ|WZ��s�?���#ں5�tm}���4CҎ\�N6��zަn�DWw9}�l�atd���L�c-��t9��6��T{L(��6X"�n/�B������í2�f+��8q��j྿�N���t��y^e{ĥ��� /'����)�r�=�,\'�7��P���a
���p6{���!ٮ�-�I����� f��bspP�O����T��+�k�e��qa/����D��4�RJ�־�~i�t��%	��%}��ݺP������e�=�z�l�ͪs�,��Z�4"D|b�� �N���0/*srϷ���;�i�pڝB���C���\MS3�;�"��� ���Wu$]Hx$�Fǲ�^"4:�)Ao���;JLZ�� D]:mL�����\�
=�I/���t�U���xx�5�3>���aX��K����^���y��5Z�@t���Ű؄KDo��e���&�1VWD #S��!��*��:�C���0����r ?Ѐ����!��l3�0�:�n���D�S�)�}������j8���h�)���z���&��^7js|��f���S�6��R �f�b,>��D�n�=1mA8Iޞ� ]嵐�h+O��yt��D<~�anK��m���(akT�~T�ha�P-\�[hl$i2"�S_c��(T�)U�`$p��L�A���n�m�0F��u+X�����7��6)��AN��&�N�|}23�VWߡw:�k(�%�7ߢ� �\��|f˃Š�L:,X)a!��,�n�r���[�q�%�S����Ǥ|lϺ��C�&H�q;r�glm>���<��w[�Ɇ�u�n*�k����vqO� ��{�z^��&��� 

I��2��n���(��Uj��9+�������g�(����O9�m%#�ǆ��������C\y-.�2����`\&��4H��r8C�%���8�|���ټ��7���K��Mc�ε�9�`ݚ�\E6�ؖ����k�D���xˆ��vK\ate�k���
����B�3XW���*@,�)ʊ��9���79�`��f�31s�)q�2�9K׶���\Y��㫬��<�@�k����̟X��@������Mjۄ{ϋ�	�,h�����"כӴ%=� g��u&x,gL��1
A*�eh����o!l���������߲$���n�>pb�T�9Z �I���O��E��r�,jp��+������gM}sC�J�l|Ib�h�Ī����쪲�ށ������ya�[������'6b���6M�a��.WGZ��`�\��/�W�����V�r�b�i�➁ѕțjHޗ���!�e��p��j��Jޟ	�G#nO���b�{"�_��T��/�S�g>�-{X'22)Y���]���yx����ջ*L\���JE`!'?��n�:�.^�����t�ZB4EI�;5�/�r��"D1VS���O�2Wf��J�%��E,~���cq�sQ�����P�m���c�׷�W ��������@�k��H6��>��'��?%�F��֖������ޑv'��]���0�WS��,�S�1������i�|��F���as�QE ף|���@��Ui�(�8�%5��gT�~l��$Y좩c>����"�Ga��A/��}�X{�l�i�v|���o��ķMa�#�ԝ���T�uG�x@Q_�y�.T�N���*�nN>��!�I��^>i��#��^����M:��O��]��+Cr8���%kZ�BY�)�N��gQ�@+J�Uʤ�ok�mlA"jX���gS���aN/�^t�5���h�z�j� 9�FN�i�j<NB'ˁͨ�Mݓ��>�~�~H�E�g�-��>�������r

�!o�W&#��?P�����T�B�~}��yR�!��c\�%r��Ҷ;>IGՇ�Ox<��wzÄ�����#O��i�t��D��,N�a��t��j���X27@('��0�Y�j��S�,i.;�����(�G�/W��yb���5���cot��;��n�r�S�-$�/��wc9`S���\Y���/�� ͈g>ӫ��H�>�zf�(��7nȣ��:!c���ʣ�7	�H��1K�3�-Bw�3`��dv�b7��("3�efH8oZd�v��#2Ǜkx7Y�(8J]2xZ@&5e����C���;���@(��2/�@�-�J��_EG_z�K�v�Ž{U_��rH$��"?Rū
_�I(��9Bʐjz*���!-j|��~�O)rY&�/a��)���̢�XK�V_��~?���3���ob�r����5�[2�׷���A ���Ik�7v��1��	�c��h�W���J�Fy�.mҿ�}��ܠ��
>�� �����c��,G ��>h[�Ŏ��D�����`�x�5��� �\����+ڢX/��L���9z7�	mD �ȩ+��C!�ۢ�}�j�K��N>����D�b��9F3�>$cfTPxs7���iKRZ���}q�S��!א%�4n}�W��cA� m^�]x*�e*�k&��[S\��m"��H"W<y?2�qUZ�w��XF����]�8���qs=��)n,�P]o���j���PP}" E�+͚߅��{�#,5:kOr(�3���h��e�Г�Q���I�bD��F��9Q��6|�t}�u��`�D5=٩�0O��s��3Q�	�[�r׬l�����s��]K�UI�"��lο�j�6q|��}�l+�wC�!�-����?0�)�8'̲c�A�����Dt��^9�n0f�{B�n�N��VXF�9�M_u���v�ݟ��:�b���?�A%�,R���Ȭ<��NY�'��s�S�mA�c$���	&�����k��#��"�o����qB�mقb�T���;��G���A�ƅ�F��_��Ӛ���<���}�q��`�9��N��������K�6S�Q:U��J�.��^�Y�o�J	���>��FHi׍���8~�4�f�.H3���^[\��\Uv1�+z:��.�pb=T8`�w����ls.zr�;Czke܀��ǿ �@1���.y��uU�9U�2�:�6�������������=�v���0��p�T��žy����)l4ī�!H
�������i��A��������v�5����5�Ժc�iy�,6����0��1�L�dG@�aQx�{ԙ�h'�J����<�\CHO�d�RY<����]� vk���b|B(]9�w4�x����5�Pi^x��K�R�TK�u��j�C��Vx2��(�ŏ����� �#Ñ��P��-���H�
/����l��5>��_rQ�5ȶo�i�����Ms�ƶ;�t���m�4�xilX�?H���6.�7�@�bqbq�m��e�?�v�ei���S�ԩx�y�ˎ���&��*��C�X�_�!M�i[�x`��zGl<wƙc�N�%Y޿��`���E�Գ�8k�K6[�N�C�:<�5�m��G	L[[ʲK�z�:�rWnM�/�!dl��Q��2��(�\^d�~��������4j4�Z�S�8]��\�C��B��rp��Y�.pT��>Mc�l"P���ڞ=-p?�;}]�7�HN��.L�����vߪ�c��9/��%p���	��]��m` 7f�`��m�G&@.k�M*��6�l�Cf�2���"�ę%(Wlb+lA��)�{rn�4m��"���Vg���@S�fo�J�㐌��{��+�,��<@��M��(;������<zi�Di���io��W��.OtH��D͹�9k@w�-�d��V#8�FYۖBAN����d��ϛ~�P�_I�VTSje�Yި�X�e*��P�ҍjj��%��c=��<��^y���[�'��@gLW2a�"5S�3���龢�?��{$��h�L��p�\�(EՌ���p
-��z�u�wnQ\_⮋����	|8����E����ϝ���j�n�V�)��?I���{��+�1��e_�����O�A���M��"Ҳ�s�ߴgrʍ>�4�ܧh���ś�-m`�YfU��[�¼�k��}6�.U-��zg!����L"A��CU�d��<�'�]��L<>�.E	z�j��P�X��<�k����݈�
�D<у��6軷����]�� ����N�ib(v����l(��b!�n�"�T�/_�A�����i�%����L�bY���п����GH|u�]</�u_`�V/WF�97F�R��(z�،a�����h�*P�eiOL��ukJ�l/��5]lA��h�M�.�5�爵���	��R7߳ p�Xy�s>dgy*���t��騝��I��"�Ϟ4x���)0л8�oV��̞�f���4�d?�p(�<� �?��|�l-���X��j������Z1_���K�iO��<`�WND�,b����$����R�1<�-��ɱG_ƦNا<���r|:����x�-�%��	BZv[�T�%�Y��{;C�e׉�pȡ�Z%�Tgs��J�����c�A�u��O1���}2G���[�l��|�����$$0���W���"���lv��CΛ�~-$楉<Nm�����I_'ra����䒍��$�!=8��̹��_ �U9�7Q�)�@�R�2���a�/��Iz�,�[�H�2$��P�ԗ�:�D2���.ʹ�[�<�k=�DB��"��c�Tf���-H�E�L��}��M�ByB���B�Rꖭ�VLW �+�obf�@��7�[=޺0�+��_:
Y��qĽ-Sc�\f�I(Y���'�6=\�bs��������G&p�]���cY̱����71M��;0����b��4K�����\�G.��O���f���) `�f�����J,�!�;�脺~�W�S��	R��z�<�Ӵl-Ѭ���U��(��A��ۘ}��Z��}mw�H=@�|r%"x�Mׇ�7��`bN����{�uz]7����B"*��l��>�4�r uP���GN���9Ha�z�J˱���YBD�j��*�w'ͳs_v*z0��y��w9�~+HĢ��)�%bp�!w~r_�UO�[��g��`߱���4�o/�g�dP��Z�iN5�s>k������X��ɲ�I9;M ^�xo5O >L�В�jG�� hÈ�l��8(O�e?B!���q+�"��91BW�[.��&jf����t)�M��B�԰��y�/��&�� ʑ4��
�u��[���C>c�S�����~���7���;_�ʐ��w��zk��X�<wqp����,��yE8��~j8\������P#�HO�X.����p ��� q�Kew��ƿ�����΀����O-̞��i0��1:��R1�Q��w��:�t��_�.�	��-h\P��u�T�������w�Y"(��RQ���3���$s�]�kh�R�yz��D�򱥅���H�CM �*�s�:��UwP������vE�Ъ��=c�`�M^a�[����Z]��t��W�#(�{��3P��le*?���9D��/�F�|U{��Uk��=�m�dvo;=�t9�+�\f��+��2HU�uZ!H0�s��B;���)��YcT��酷��"��
��H-~P� M:QٌbUTu�e�E���7_�ls���X��ق��,��0@cB^9��K���<`�����U��t��knu��x�рm���_$I���V=�Q����-��.n��!�y�Cp�����Ul<�z�C=���=�C/�=�Ϭ[�G0�޻���:pume+���Q�>�Qn��lN���{�G9e'��v�tB�+�v)�ZΞ�Zӑ*U��8�row��t�7�t�^*#�� ®��� �Y )�"D}��-���n��;ЛLs�ݽ��ç��`CaY@{� ������R��F���t��E%��7��ܴ8�?q)'�]L��a�򔾏�|�T!0��0(cA�#����$��[�j���v�GfԶ���q�ry���u�!�c�EDáx���5���,xEZG�I=}r�)���&��s�4��#��J��Q~����H�6��ޗߍ����ɜty'"�^��1)��(��!PW�	'V[����L���g��w�"G�	h�Ce�i�]��GΖF�j;�����I�8��]J��R�`��W�gw/�z���UQ�ލ�����˭V�}\�[y���B'�:*���i%[�k�o*ʻ�Y�7���ƾ�7�4�}�h{z���o�*�c�ф�b���UY�\�	~4<��$�>�u[�U/> ��M��Ζ�^noc*��b*�S:��^w�ݖQb�FC&ο�C�3gP��	[����Y���0��~�-,���|#��+W����r@�f<��Ԗ:�%݂roW�g:*���TC<��Ѵ�b���F�
��P)/��B�&݈J�_ܹ��h���XL	��8��G��t(5���GBt,�p�_pTZ"a���������g;t`�{���M�ѧ������j�`n�4���'EG�8$�����Hm��K��`�_���6��Kv		�-n�4#Q��^^x�7��A����H>��+̱��9u"�\=ҹ�H�PG B��A��$$Q�4�rZ�ۧ	Ҝ^��3�N�#w63YkE^��+������ѡ��'�)�I=(K���7�Vկ�
��s��6B�cF}��τO+\m� �!n��u��-�Ѡ�v�;�/6;+��*�����}oЕr�ҳ���g�C6v�
��B������nw�T�U<�A�X�f럐�wi�%�eft��cA`��{?��ߥ9಩�I';�_-Վ_G��y���UJ�ydz�	~��|�hE�R����v7�a�5�׀���\�,��D���-J4�5��r�3X�{��H�KG���3)���uUd�qb�O+���F�鰯��9w�ܷ�G�z������G��W0@j���MIE�,Z�t�"�_���r6v��f�<�P=��?:r�����ضD���,Y~�S|\�|RUkg5��D�3EFÓ.�&�A��B��z���{w�L\M��>�J�i�e8��h�켠���H{>z0D�osxm�bx��N��>�Y��hI�w�9�.�o2��f:^��V�W�����ϫ���,Z��jC�	�6SA�����xB�<�MFT?�O��[��ٸ�{ޜI���&������ҏ����w!jX|?N�a/*i��*%���#�v���*�'H:X�=W�Ct��jwE�gSGs��ͨ �Ig'�5��m�-��lZ����>�O�?HE���
vj��	���<�>.vYC��J�[Ef������s�e���V�13beL�ngl�����z����@�:��["��ķP���b�:�V��V��{�7�2����r�:'�k�,B�u��Y̆�Z��!p�f�-��>���|ͫk���x
{8f���`ޔ�N�Fe��:_�*WTF�\��(Z��틦Q�|��H�pK���y�`�!+���W�� �;�aH@偀lý �:3�q��D�uq�.�_��.����\WcF����B�>����&��݉<hs��[���ӎ�]^2`���`:��|n�=�$71�l´�a�R(@���*搱ԹT�9-�­%
������^��ݸ����7ѣI��;Y��̔0��n2�Ql�o~��v/J"�L��Hi�e3,M����r��*P Q�	���������s���,�N�
l�L-�幄�~	z;`��6����#2ZV��K��Q�Qc��������V7� G(M�	�#C�~�� F�C�J���5��r6�ţ���@��a�7�30�J����S-	�޹�������f�ܰ܇���Kwؘ3�<����e�)#���֪ҧ��+� ��p�q�E��*��_~|=$�͑=�������]$����;t]���N�]_�o	㤟�J�W�z}��{�3Ϳ�ſJظ�s!W���{Ԡ��9����P��,Rpܘ�xN��[9�?��11W8)�����m�G��d�� f���4�iFh�is����� ���z,��݋�d�ssǩ�ս��G�/l{O��F�_����,�*��E=��2�YV�� �t Gw��@ɪ�!d��N2��Q!Ҙ7+O�"�X������F__�|�h��
v�N7ku��J{�~�
ٷ����;X*\3��x��X�P� W(\>���*� 7�4n�����׫8ofF8���!v�Q�	q�[� ����T?�l���d���58�M夁z�_=�~I(lXPKK#@�j�="���)�44ߵBz0
�c������?���d�]�Xى���K��7 ��*����]���m�:l�h�w��=!'�'fPˬ�G��[?� �o��Z[=AA����0����~C�5rGIVe+�fG=m�L��Qx�I�^¨������\�P�e���r�
�ϋ ���K����$�+ X�0��{Gf)����P��6��,��l��r�O�ρ�k��ۭ$�oR�ϙi�0�e-�<GN��ث�香���A]�<�yP{�Uh�������\CDļgc{jqy�8{Ӡ3��ۢ|�ڤsb�I0��������R?z֏^r��11�{��l357ϋt�%αj��\iV7�k�����������m:xO�#���D⥌���iXe�u ��(�4�m�q�l��W���C�*�iB�K_�JֶȻ�X~0��[�����a� ���9C�xt��Z��T�����Uc���@�шc>�4�@�1	;$� JL&ejN5�d�	�Dk�Z�oN����"�*���T����j+ዃ��Tr�$t��q<��Nא�f�����W(v1Cj�#��~F�<h����X1�P�[^5����ɮ9KZ:��n�_��W��T�+֥�*�D�׻Kډ6aY=YuN!�4�տ�B-ZYQ�ˬ�+N?kA�bc�|pڝ��%�j.Ϟ|���y��-��]�2�~z��&��e��N��ä�VI��];�F%߫������l��;b���A2i��f�NF���ka�����gO��n�ľC,�:b*'sO��j��s"��˯�z�
�2q�)5���'j���ƔŽG��v5! ������u 46�A^��ߥ�iz�����N��l(���m�/POQ����RZ�>C�
LG<��5┗9��&ɶe`?��i�3)��(�f4�^�!�ؑ��(�͘�o{���{X��KU�9֪�����;��ˊ/�������z�!v��D�S4��@7c�N�|��G�5��6���ԕc �P{E����1�p��y���>�mS�%h���HS��{���X3�Js}6��p�Y��-K�S�p^4߱x>��|�+�m�ݾ�g؜]!t Yڂw�u/f�+����f��0�vh���^dz<~�ƶ#��eKğ��_�?UW�]���峼�$z�}����H�u���(ve@����7�u��Vʶ��{�ʴr����3���f��]֌K���oo���biA��/>��R��]kç�Pä9���,��\Wr#i|?U��+w�w��X ���m���o*��q �vP��"O�}ɞ�k�xf�C��F"��L�;�\%�3� 0ނ�GL]�<o�,���C���B�l�G�Nq������`q�+��u,��Q��EY`�NLۏ���N2u:�(�k������J�߃����T�9I�di�.Vd� ]���"�!]���k��`�!r�*���H�0�#���A�Ī9A��ͥ�2b���r�.�W� @ٙcub���!yť��HF�SM����ĊJ<j߂=��:�@�$�Eݤ� a�A�����������I�I't��r]	(h4�8��O�2��b#ak�6�����偩pcc���S@9����s����[w�@3�ZG�SF*���hѭ�[6	6?	lV����}&�q�i<Y�K��@�	kh�d��
 ������o�a�d�'J���H��h �,�-���`���9�6*{��E�������|�ES�����+��h�/�/8(}��!���&��Ԛ�U���iP�,��c�;2�ǘ��f�=)g�������_��,Q�H�*�Q�� �*�
�y�����KBx����n�j�zF�GyR��W�j�B#&v�����M:�O`�����`�$Ei��
��$V�f�]r�˳ ��fr���^cG�Ɓ����L��!s̴�f<n)\;������P�
!D�ESo��#�hE+�D6O�� ��f�������I���6JY+��x)=�vUF[
��R����_�,"����k��Iܵi�"V_�6�x�(��q��`�sB+��dpfC��/���9O;�Q��%��@ȉ���t���N�^53w� �f�V��T~���`��r�L�Ӕ�������tSC?u}�}�4���G���o��4���n;C[�ţ��0��T��O�������4��.��n�`~E���Bk�f�����	~�9n�I}o#�����x��2w�z�@����
���/,�K��&��;	����%�_p��w5����dwb�h-Z&� �ɞ^�H�uS~y�ݨ�F��T%�v��LQ]!,}$z'ң��o-�6k�'x
�2dC��{��@|�$��ɣ[�g/Z��-�؛8=8�x�h쀎�Z�k�k�m1�ؐ��jvnQ�Fσ���֥3)BZ��^q޷�Sf��:SH���R�Ν�8��Ĩ���ly�l���]�.;'wj��F���.��$�U�K��A}E��cb���V1�^��E����qa�-�gJ:��$�rds-�}��YIw+:��k�L�[{}�١�G�f��h1z �z�?�hxp���ѻ	����QNy��Q�h���q��<��#�ʉ�����s�����n�:O�����f�����V�{�@u}]p��н<��_���A ���}��������������U��h�G�*4�Qॲ|W+���_g��;���K��]����m��h��Mz嫮��M�N��}_bz����F?:059���G��=7�	�\H�-��0�WO�T(�;U;8���8b�k����Ɂ	�~1��@��K�q���0+��_��L1��l�~�v��v�Q��nU��Ft\���.0
Z�U��k���U(*w>d�,�Lw��y�.O�<6μ���
I�jb9������sX0Y��B`1�MQw��shi1}S�ݷnb�,�q�����J�Oݸ� _e�[��`:ͽU�XTT~�:ڣ�!5>T��^����I�9Ҧ=k��B1�1�)�`������w��[��#��5�$��.[��e!L���"����y��FG��)#���׎��|��ju-'�.��
��*[�[�y]$j��Oa8��'�7����!�����A����w��wS����"��CY�^��$I'#²�L�qA�-�%J���;���}PV*1��SnY�]��`ӛ뫽/���5 >���;~������e�?�C9�ğ��9�5j(�J�1�������9�R�������3�I�� 4A�����@��,�{���b�"�&�ҼJ�%���z{N�?�)�ۆxy�+�|8�������F���ek5ҕ8b�p7�&���lk����fH#�������:y��n9�Ƃ���p�O�b��BӰC�]+��7�X����� I�X8��X�U&�IO�c�É�t��(P��p�xԕd�YǙ_�&�����`(	rСk��u����Wlz*��BU�B�2v@���� 5�:�U�d���x��9'
�I^ͫ0V���_�9c�C%��{=�<��)"�k6_��Q�w����˭���ؘM'
��d�c�d��/G���E���]S�6��*�f���%�uE�a�p(��s�6iJ�:�t��i�ܙc���'��X�]H��}�j�Ӡ>��!kD���8��8���L�[�f9L�e}>�O�\(Y ��:����c���ev��c`��!�@k#��JM�_�Y�B�c�0}�#y�T��CZ����g��"=�]R��Ƙ)��C��Ӏ�`���r�&a#�4��ohfӮ�e@B���]˳���I��t� c��mT���0�� Lj^����!͚��^<��0s�w�99é�� pJb�p�6�`qLS#�_*�ʌ `�X��6��ʺ"��;@g�a�{MX�q�7/�E_� ���d��Hѩ��r��bi;;BBK����ڏ�3Aw:��P�8����(�A��T&�`���,2@�yʭ����H�� Hh��;)�!�>`����^q9��AAL�LG҅S���	(��Ƒ1��]�fћl�W�B��-��)��c�����WK����
Cj�Y�j�F1����?o�U�f�,�� �AKx�g��J!���	=R]�-�r����V݌���a�]~���2�Sc5�'�(|�i���ޛnl
���6�X��Q�N~!D�/�&{�E56�3z
�����@~AU!k��z�V��7r"��3���iFonp�ѓ�s�c����S�`y�Q^+�~r �����+BTK⠝ɾ�q�HW�%AGU����NR��陰�B�:5 %���-%S���ō�Ԋ�ٗ�$�X�I��ʮ��@������W��m�&.�	'��W���Kj��%���8N����4(���ۼ�毻Y�8w!�`qv���l/��;��H�'lcI\r:��`&�Q�� 27ȯSF��m)}�넎�!�RP�C�(�g�/J�4o-�DD�4��@{��PO؁+�<�W�����~��nYA�S�I=�:�� x�2���Tp�Z)R��;$H�8��S��A�����,	��PfT^u���őWJ��5�q�c��R�RG�iR5��66K$�>yR}���y�8��?��NN����Z��ހ�K��0o@��S�6NP3KV�9ӷ1P��\O��s���j�I�e0�!����i�(8)��	��% D���OR��1�#[�WH��R��x���~������z��%|�^u�#�>XL��`��Q��-�_�}��ݐG]�Ӊ���&h�?�&{�:ȼg-�\�,��qإ��f�l���
*v�\T��M�0ٰz�&��K�un�ƪ-ב�:�O�Q'B��6���\�|i�)���6�}F�Q�w�Fb嶛��[v5�i	��bqM�0M��|j`�Kb�4w���&��\2��Óֱ���;�^�䗢���"-��G���H�@&�ʹ�H[����?v����{���\����� ƕ>�N��a�t�~��EH,�L:��^嚟�T����C�r$ğ�ڔ�+��Gs��͎�#�et(�hQ��n��Qm|/߽������_�I�W�_����Hl�Ur5s��7z��OӁI
�7@Z�lW3�6�gј�^؜����g�P�]X����g���г[d��L�W B<D@�l�\D,��}�����q���ǊJ��o
�9u�t�刊�Rk�i�a�O"EC`�dh�7A�*Mԃڗ|�8{/8b .7w;�Sg�\��ӃG"���P �ސg`v��ce�u�|Xȳ��R�[���H�c�>ȋ�@�C�p�|���gFvgK�����C�p�w*,Nܤ�Ӵ�j��7���|�G��G��o@-�]l�/�h1*�kl�F�e�z0�%|�M����5���(��[�#�����c�/Uꂣ�p%��04p%j�=�����mRoM�8n�)���d���<�iu�y:%�u�#.���t��a����)  ?pBK�Qrڻ�[
j;�	����
�l��a�ʡ���H�݊%S}N�AY���ɪ�
q[�8�c�8�$ s����%��A}^IU5n����$>O�3����I�P������rT&]�g����1T#�^�_Za�R-�����Sq�$#DI�<Y祟?�`-%jT����t.���]ͺH�:�:�I�A7K��q}�G��Ξ��ز���zE iY��"�,=��K��#���&� B���,�I�BӀ%���`Ѡ4 y�\��]��_&�z�Ij��7f������LEՊ,3��0��<�>���S4�N�)�]�v��.��v=�=�@�'��M��MY�nujȿZ$L�W�;r #�}Aaߦ$��%�&�Z62�`���zw[ۣ��Ob0�s�	II��q�+�����CN\nP����N�ҏCN(K���z7�	��fN	�[.�w���3����|kf��ﭭ�Fs�d��G�	�s�㱳��=�VW���*�X�`��.��v�W�� �w6��+?����ǿ_پ���KA)h~�}��������5&`�F�?@��8>����@u�TW����r��<�;�(��l��)�!�4�r]_��aN��SA�#��k�7��s��f���;�����/���Ű8n�J��#T������}f) Jh �H`o!U4:X��Y�(Q�����pך�B�gKzl�9⎱Y��k����d�#KY������[c����å��L����%�TҨ0��P�[�����w�E7{�ϖ�U��_����?�q5eF�k3`j���5�.S�2�d��7������;^&xk�X��,Ϭ-vC`�K�\
�SG3R�}��t�!�p���)`uM�tx �=%�V�"�<q-Ky��N��r���d��y�B�)ߤ������ Yb�Wi���̝�T�窸��ﲙH'k9gz�Wbf�TjU���i|�=�7EB�p�1�ύ���AP� ��)@��{��7&pbyI��/ �5�+��A���	�9l�@�K��o?�x?2k��>'�6�D��2�^���� ��VǐjH,& [�K�22�����Q��cZ!�ƶKx�����w�O�6����}�c�� �0�aLK�UE7�����C���MP�|X`ˋ2��X��b��̂Q����(>��&Ho�������a���6)N�8�����QϿ#Vr��m�b��1���+��r�2�{�e��hQ�,��e�>!R�����?�=��ixBC-��#��Rߠ@Ar�L*͐<0�������OP@���� v���9@�{�ļ=J_���N�bQ�:��*E�Ǉ���d�7��u���������m��[�{�qHD�L_�ui\hN����h����z=v�AZg$lW�8����n\8ƗIK����.[Je�S�~�?�O��፹y��{J�8]ut�a�<�O��)����j�fr��I3-��uLM���ښT���v�<�+�d6y^{p��;ο�$�����_.�Ԝ���:*��6g�r���$��v�'�m��{bk1�y%η�ZnM%���ѡ�ӫ(U=�N0��]4�8wt��@�4�)�_B2��)��Uv6�N�<�;|�<xʯ߁�W$k	��ӭ�� �����m��J@,���#칳�yN�Q�ʼ-(L���E��L2V-aP�%�6���� ��B��d�����) �h�����(I�������+���s�ւ��K��ł�U����ۨ�=,��� ��+���� 9���ʳJ��"�bgP4ڐ�/6��0X]�_��so����22`���'�K�_, g�̩ 6�S��הү~�|�J"w��i�!�	�"u���� <����bt�m���DU�-������#�cӨ�*8A��θr���t��Bۜ�ż�ر{R!�^�D��"��;���>���N�<��V���3w0@�X�}�x���O�񷸓���� ��� %َ0��*QB����p�ξx�0�A�#�l��
g@bce	&,M��sp5�:�+H�r���o㇃�#�|����y$�g;�ӥ���&�s�Ѱ�C�eb7K�>�<}O�!����~7�=,����do�xI$+��x/�:Z���E�vzC���
��I�z9��V1�\�5�O���{�ࣔ1�W/����o(���
[Fu�tkԹ�{�V��S�d>���W���g�D������n����:W��e$C���P�.��)8G�9��Qq��F+y�ě��5_�a��z^5f���:���	�a��V�R�sBsh2��fæ�z���64������ؘi�ҹ1�F�@�	���$�ȉ���Et;ь�|L�$5s�F�p1���hu ���C7*��K㚸������=9rJ��Z�.ٌF@
�B�U�հ���[ ��˅�Eɥ�)�r� a{ ���pR+�&�#+��k��_��W�"���<4��1k=1�PQH���3ד�$ѫӢ�F�|g�g���WV�W#� 
U-�n���
�k���M��(��M�{^?ȲVN���x���h���6��Z*�,��:�w��w��K9>�����������ܨ`����F6�����Z����
�g�P��~���Q�2J�?�C�����2�JG"�S���Ѩ��x<.����s�^��x��7-n��]�RwIv �2OF\y>^Ȉ�4���z�:���6�	��f�x�A�T>
�p��	���r�w��w��F�v��$+B_<t»(��0��#�v^}�	t����q�gc`�~�F�՞0ADދ/�[�{�#�W��� 6L�ě6VW���|����L1�0��>~��CU!�����ǽ��r�\*W8��F&a�㣗8�+�`8�Yhn^u�G+h��YW��/���,e�a$&D�G�=�3$ܽ��mQ�M��[Xl@�/qh�`�{F��ƕ>�p�Z7��^�E��`�N��cd|ނ��A|Ϳs3g�ز4� -C�uA���}�����5�*M�]�F��|�!���
ԓ��t�6��h �?{sm�eI�<�~ I؁�.�b����20�IYV�sJ"������MM�$[��jE�EAK���4�ۿ%�]p���<(��)��,�,5��+�hjA��4��@�¯���1�i6S/���k�WGJ�l�����ieH�DU�2:_O٫�I������h{�؂�����|���o({�H������YXȃ[+��E}��_�P+%c��S�z�*f7oD���}3`�ު*��;tz�L�D��:��J�Q��+���w��	pŐ�4�+��8'TV�sx��K�}�z�9��K";PSdY�����rn��A�i�/���ʕq����L�w����I�BLqq�9a�6:�(1S�*��q�0\�uϴn�%�,\�����W�9��"��EO���똂tQ6X\#�da�y��yvޠ)�{�W��1���?�����b6��Iw_?�JF[���L���)"+ؔ����������Ġ��h5�_([7B�~�^�Ni�����	n�9�!�%-�n�g`�җ�*3K�z�KnJg|�;J�,`��t]u�W���.�asw�g���U�H�S܂ߜ�D+�݉��k�x�.�h	2o<+��:v��(髇�#Qۇ�0�4��x!���H8��e���0�=5�r$q���/
�����@�LnGV�yax�7����
u2�L�o9[Ɣ�ю��=�#���]<&�T�E����E��ն��H:��D��B���*'k�SQm�>�>P
�DQWʟƕz�O�ܟ�vMs��ݦ|�CnꖥOzj�o�Y�`�C�R��^g��5��)֡TUl�_'�R#FS8L+[���{��'L���\	��ن2N�'n��]�q\:����}�Kw;6w��F0� =��>e0��?������Ib*���Ċ��ݸ��UH�]����.�4�3� f�m�E�Z$�>RR�06����<�Kݨ:a_�%�*�{8OJ���f��9���?���f�D\&�؝�nO9}����xDG��F|��F�u��$ :�3�|����]�Z+���J��x�/��ّA��_S��aѳmeO� &&
��h�9'6��؇�����:V��]��[�/�zʉU	��q���O��|�A��X��u��,OXPg��ӟ5p��P�B��gK�܂f�R���{I?�&?q�g"��j�A�> #�M/���?��8�cpL${�8��
W"�9�;;�tX����j��3w�t�7U��M�;kQ{kYD���ř��W�I���sk'J���Qj�o�|���H�+a�C_�Ͷ���r��	$I6�E���O�X���nw7�AK���Dia{b#8�� �1���y��eo��O�]*�#H��>�k��%�P(z�S ��Uz>P	����jV^���O�Ϧm�_�5�?e�!�_�W۞�)3@)%� ��8&�ù�ϭQp&y��;��/�t��C]k� ���2c���50��\ ����_���Dn��1�n�J�j�:`~��l��B��Q1����.�S�eL�nSyk���������8By�|۵Ļb��鵬���m�>�"}vT:�v�2(�Br�c�Y�#(N�]ܦ=�|ɵA	����"k�0��B|��ۘgwk\c�_�����Sk�i�u'��3�D�r�{4�1Jo�m��-�P��~YE�{�g<$��O���U5�c(�/����nx%9O��l�>���%7���3�1%�-,�g���O�?TzEf�qe/�m��-K���2\+�ms�U�Gq�Bj4���#�U=dZ=(�Ջ��5��S���A�`��,Hrz̃���CK|6�������Ե�Kc�eӏ65�"�fT�
�n�{js̼��Z�n�e�����׎U�lo��mz�(o`�a{�P~���̃�3�������^�np-Ϻ �?7Pm^��Gn���pw*������װC�!����Vn�	��|��5�&����2�Raj��;�K���B.��6ЇO	�U0z[��v57����*�!��V���\��(���G3��W:�f��|��O��;�K��Υ����Y/������K�ѷ�EK8��_�r飪��:}�g�&KsK��e'�v�:�C:�a98DA�-�v��vC��m�TCR��2��ȶylO��P畍N��}X�x�$����W���Up��[\1�c>�!�=Zv@x>J�Yw�i���	�*���:�
�d���#��(���})�3o}�ݟ���;�>d&!��i"Ft-�b#�!�`v�1�$�i->�l"cw��o�e�N����	����G��YΨk�L|�L��� ���[wrX?"��7 �yΠ1� Y��t9
�ޏa󗎻T��Hх屟_�a��^�<��y����F{��>$�~����@#�w��4�7���a!#q2*;ܚZ�	���5,�M�]Pm><>��6�z���ICr�ߢs�
7mk�jDQH���+ �sX��P��}.�<Qښ7��p~0q���gU�U�DP��JWߊ��O�m���a�+O�e�����Ή-Fiy�G�JmU�/ɹ1 ��W��B��O_D�z��7D�)��W���!J\¢�F�>�*c�*�b$�Z�V]t%�����G��EY������"C1���vs�X��3��4��1d���Z
�� ��p�����%_ȴ�K\�&������r;�5��
�}���M�8�(Ψq��)�~)��I�������0�F�G�jz�@�(�=�S̥�����:��30��浬1o� x��2���I Qti{Z=�,�sq���n�G|b$��I��*��N~�O�҄N���u��,�w�Pdo8�cB���3�n iv��۳�e����9?K����j��G���o��jt���X�u����R��#�d9�����q�z3�,�������=�|��{��i+/F��1��
���Sy������g�G�ީ3���ߵj��Vb)p���<�q�`M#a���'��{�u�M2QO%T��w����5�U]��up3zjq�=r�=����"O@������]�"�j���?���OV�qSvt%�8��S \�9�������l}Tj!jp��hk`N<	��y�e��W ��9+'e��)���I0<#iM��Tؐ��E������)���'ΰ�p*G�w�]��n_=A�D|)詫���VL���$����@� �=�kHş��,�z�;�N�'��[ˀ��_|�������DiP�Iߤ��xM���Nں�v���fgD�cm�P�Ɍ�]��o��$*��z���ɋS�{�1�ʱ1���)��j)�1<��:���~�:�M�j ��jИ���I=���y�\��q%����ĉ<�!D�/$���4���~�:%=R9�pY��ހb����E�O�kn�1���)����,�ƀ��#y�E�x_t��Y洈mC�-βA��;]�d��[�љVMK+n6�3�W��Z�I �]o��u�(�;�Jq�c�Կ�HO(L���
z����~��
�"�,��->>��͇QdI�4�p6�.�Q���9i�n�r��o��@��0xqX�S؂`��Da~�$A��+P~���uw�x}�Bn@��Zd[` �c�n�޵���G���6�[�P�fWv3�?�����C�;��}A�ea�$½�3o)ھ���i$.�����=@c���B�W#����P{�w
�N�m�V�Ŷ�x�qw!�SF1���0/L�����7���܁��{5	��L,�Y�V�(<��C�.�»�ă�P	�:Y�ߔyQ���|��D���A̢ŉ�9��)�LT�^��4mW�@�c@�6�K�g��(a�ҝ*Bzt�2R�ϋD�;��{@��0ٱ1W㳜�m`'�{����M,� 07�[���,�p?��yG�c��(�Я�&�y��tS�M��F�g�e�i{Fw\���|�"���%�W�n�#�V���9yx��I�%o'��"���}ߩ��w|P}��}kS���5m`X�#�p(�B���F2z8��鳊4�Q�U��VW�LHk&�/�(�(p5[��)�՟��H��=H���Y/�\z�~�f�Xǌ3��_O?(��ѐ��jk��T��p�Ӂ]N�$�}>�����%M2af&�LX+�����T�)��_X�q�������}�m��Ŏ�[��N�^o��AE�c&�2Ɲ�@�(�Zqݯ�ࡉ���:�Ô�q�"�|�6:X]��?wS�{��E�d��oM;��;g���ކ���^�Pd?9�	ڔ_o$�Kʖ�C$E�s�p��3'��(�o[�������)p��X��k���[��崼�y��d��|8g��3�����D�����������ٴi��[�J�.;��i�r��$�^��M�Q�nY��r �Fw�E�'x�˾ҩuB��qŃ-f��2����@a�3E�����U̾өO�;�ֶ�
��0�ex�X#�?K��bF���#���m��;����g)����YfG�k֣w"g\�x��ð�`6}��E6R�h��[ \k̊5$0���*2C��;E��K�F%�"�H�׳o��3+���z]}؉��S?��2$̥��ߎCI��=]�� ����M1����.��듶f�W�u���]C�aqg7�-��r����\J0N;��#+����[F_{7xr���9w^��q��G�F���NHf���fQzx��r.iiZ/����7u��(���]1p��΅���Uk�B^��y�[$��~i/yj�o��E\B-�Yp��w(^twU���i4�֞=�]�X�+��	�&�5��bN�M���Í�u�ǧ8ZJȇ	����6�>9�J�5�T8�0�&m�;-�:��~̯�ķ�����YPt�?ngF��1�^\�Pc�̍�7t����7G|�~�=Dl��(Z�H��/h�Mj�n\A��)�i���Y>Kou�{�'`yO����
wnZO3�n��
�X�~��)�y�`|��S���WM!�+��$���gh%Ӵ]�r�1���^��@��(kLy�§~L��j���������I����x�B���,� ��%��i%8�M�	v�K�=a�8��B��]	^Hje�����8���y�P�����"�+�-�5F�ʨ�1
��덶���s-<����g	�2�d�#�<���\.	}��J$�,K?$��Q�az�Ǭ�݆�<�~8�9��H�&�,U���	�W+���C��¯�B�j�u|��5����Ʊ�f*դ�ǾՍ��)��ʑ@�#V��7(��ի0O�vG?��Wɥ'�{��~�{(F!!D��o�T�P�E�;�$��OKl9ϖ�=���Sa���N��6|z?��>Ѡ��H�&�#n���_B��Q@��[�S�N���[�,a`s�Qiс�ش�/ ��g�<�r�F������f�GCK�8�=U�c�Yf��O[[Q�d�����#���,�[��XX�h;�ާbʗx 5	7ʁ̳q���R��(~QU�A��G�ĶJR���v�n1|�߅Lp%q��Y�u��e�'���ϻ5��(�|�s�.H�U��I�ؔ�k�E?[d�z+#�?�Ȥ�f��K�0�:��<��t�ĉ�]/���ug�Zv��aI�Z}>D`��������3�Ȑ��Q�ȗ{��V�aq�����Sib�b������[S�_���"=w�5��K����tjh� p=���׫ɴ�n�.�����|����֫z��,�ϟ`�*�MDT�������,�U���(���5�%�ET�o����g�q� 
�qLjo[�BQ��H�3���S��
�\���ܮ�pJ�E��J�R3|hri�uv��<UAUy���~�x]̂��[��5�#Z� ȸ7��9�c���.���~��Ґn�F0V�M��wy,x�E�B)b�^P���v E�؛B~s�,�T9��	�1�X�F�[\p�*�$�5�>��BU}��«��N��M��Z�6�ft� *$A�n��2��yh�&:�nە��;�3m�����Іk-��zSh����vT�����'�-����vHvYg��O��7B��DS�<�[}'F70,忞�TK�+�$�;U�*����r4p�'J%o��ra�%?�x��R�R%ST=�&5F]kw�#�J�Y�S�^[�O���}�k�y+�k|�x&C�Ir����<�)P�j�|�T{���T�+Jr�a�bE*�k��<f�L��kk��j��.<q���^���gi#{'Q�G���C�$���c���s�]6 Wn��]���hX-M�j��A$ۓ5b�
�(�!������%�/���y�Pg����jY���Q���+_�OV���6P�9�#�؀^�4��M��*`���7�^�]٘_���p%�x9�(���P��!,��LK]z��'��Vɓ.)�,�jTd�+�m����>�)�ۈ��Ǉ��G]�t��:��g�h�������p/�����$ߑ�iV����v���G���{�E]SΡ#�=	p�~����i�v�Z��Dh����q�����{�<^�C�*xc�ڿ�������þt �H�w�gg�D5�h��P����dZ�8̀89�k;ugk!=ڣ��w\��x	��#�G��B�f����=��?��#�b���l�Ä$�P�R/�e$�p�.�h�TtȘ��>����)B�n����2��e%囔��Ba��?V��U�Z�|�n��I�I�F�ȵ��_V٠Z�XΚf��`#�7��������ʫ$#�L��=�N�r6�<��(>ǡ�d �9KrKm�k�P��8{;
\�Ĺz��Z��UJ����E$�~J��ue��+t�.�;|*����CP1w��	����ip�;!iI����@��j����*���My�جFA�b����"��h��mB1L��_���TVYZ���d�o��T�R{pt���y�Q��d@��8���/��.y�0�zP�!�3R$��;�
(GU��v��m�:���o6Q6I&���8G�c}�1m;�:�7A�V�<�cjs�(��6y�-��Ƈ�ail�w�ʀ:t��qe��c5��|J�Ao[���tO��-1;�ZN��]8��!Ɂ�Rx7z)?Z��_�`O��Y�y�WO\�2�z�QJr�;���("ـ6o��/ok!)|>�0���`KF(��+�V�s��} /]+lN���t�CM�fB�xp�������Xt@��;�m'pۿ��uS�(K�����/�M�!��K"8FgZ����V
|�i�j�G˸ſ�2q��@b���pRΫ��W���v��GA *��8���0M-7oRY7%�tQص��i�=�&%�V��`����,)'��]}z��\�t�y6G���s��Z.���V�����J��.*��i3�P8�~�OBsLY)����e��2���Cs�2��@����Q�+������u��C��C�ّ��V��������`�@5�Tm<M"/}ă�dxi.�WX��' �hY�O�;�)D~��r%�y�� �)��8��Aϐګ�#;=(�NG@c�њ&�z$���k��c2.��yn� �ޚ�2�`&��^�;M�޵���9}��/�c�}�_�hsV�@�b_%s`}�gM���[�3�@�Ū]�kz���){�c��UA�c&CA���<&�h��<�e"hd�͒���Ɠ<Ľ��7]�-�:6b������ޗw���j#ㅫU����S��֕��3����y�)؟����~��8V��ꨗ�pi|ܮ�CEEn�g��/ m����tH��~��� Ķ�����ˎ^��>٥W��n��0�|e�д�£�ذ�D���{��#��ʧ�t�Y�5�/���`�Fpv_uU���M����׵p���2��(��05�B�	��D�g���_���+�k�f��������}�^�5����I�������s����>d�ں^Fؚ]{Z� Z��J�'1�;����	\�0��	cʫJ���Q�pW����~�������$�P�<�r^��W��u�ӊe���M���᱔�ƌyd��R_|�WCێ�ST�<�F�(��Թum"-����I���P�9X�x��A.�AV��e*�����$�q��~����GΞpv�֜��������{�a���h��7��1����K#J�г	�Ҟ����$)�u��g <��ΐ[�^\;
`�È0B9�9	��J��,x�Y�3�uZ3l*��輵Xs(�XJq��?I�ktcm����\�Q��,l?�_����ن��"Jp���%P�6r~(���2�9c(�g��lFA[��I�<n����c+�0h2���xw�_�w�����|�reǽ�J��(����E���I�f2U<���'F����Kd�����8%B�!8�6�n�$g ���x����d
�q�覶C��X�����:�X�����A�Y��5��˥C%�q�x�!U�>�ŵl6��S�y�F�~tlOo��<�/.����YRl�����Ur�� פ"��M�ȯ��NpdCM8��C�4�}�4ް ��
Y�U�t9�5���m�BI�!�J���eO9�z�=ľ���m6H%�i�zR��������l��y�ɵ 8Q����9��c˙����!�k�O+[J�n��v�j:��`���ߺ�zP��a�'mL�ݗ�ݴsa2�Py�c�Z��䃯����芗i�<�L��Q��p/,#X���Kt�Uj�����I3�ƀ��m��(!Pl	��h�c���/���ڔ���$�FI�
z%p���w �H�y�Dw+��'���8{�!��H�!.���KX�OȐ^����p-F�ْ2��n��p���J����?<������>���i��g�x-J��E�������� ��P�9遂�Z��]mpM�Zv|�/P�/y���iV���c�vb령�����^�t��I��ߌI=��Dm��-��M�"��K�v��N�tR��a���^C>Rz�r^h�Ğ�q��hG�Q��j��L2��`��
W�1�kj2M�����j�ڃ|�"�C7�����e��#�[��\{x�?��we���嶣R������rKdu����3��7AJK�H��%�����8���]�F��qY��:�׿��K�Rg���7ָ �,[`�]��V����e�U�9G�����3�=y�C|���O�фHr��^Ĩ���B�x��jѓ߸;g!Ӝ�� 0콬�|���w��{Q�a3&�Jpm3bA����iQ�v'�p��}ee�*0O��.��nBH'�����^"3�]�z,�����"�?��V�F�:*�%�V��&B�Ϯe6�-@=p~�Jm�`n@��=�̑��)��G?���$	?%@&\p�c�����4%�@�VW+w�	���k���dzs�F�bW9Ȗ^�G���@h��p�ni�c,�Y=�ٖ%�U���r���>t{�yq�y�ſ�I{�|��������.�Gt���MK�,�-|Rc�eA8l���a863��x�zL0�U��-�e4�8[FYkuD��(�Y(�?*|���X#��#p�L�}�J=\����66���&���ۧ@�]��a�9��m;�(u�x������M׌�Sܑ���M��]��a%�+H����a���� ��tp��〛�VJ�$������"4���Ą�;�^Gg��4����V������M�{��LK�?�qOL�O����������m��٢&���S=.׷_�C3�qZ�@�����oW��bi�KfMBHڡ��
����J~�;�H\�V�@b��E��F�ܳ���kI�lͪ��=�Qt��}����U�nu[n
fY��jbQ�چ�\`U���B�ߋd]�c�Y���)�����Z{�r+���ݏV��s���0 �Ì݁{�nN3�cc_h+��/B~n��d	6ۍ`�w�:��"A�"|�*���f�X�HĹ䢆V|4x�m�i�Xª-L��NV����OM[���Oj�7���;v�l�m�uCL:�"�f}�Փ�=�2�s]�ra�#ҳHzf@Wҥ�^���-���a����'�{L�]������At'0�"N7m֦C���9���)���/�~R��lf��氞��/$�9��4�r4�?��>n������1,�_��j ��4���L�����b>���?#�@Gx��M!@�>�/@�q;����S����s�}���o0`́P?�L.ⶫOv�c�܉�L'("�����D��v�*�9�;��Q�a���N�} ��q[��]�n>ATt :�s3��d+��,�r$�<�[nφ��f$�?#����kau`K��N��S/�
��g�����L.�o|vaFCOo�ZM�t������|O3<N`�~(J��٨��L⭸N,��
8���X������$=�@�Y�:*�2�۽�9dpT���=?:.��"9���#��\��� �O��q�6�Q� ��փ x�H��WČ�J�m�)7�iU��;���:Fk��[��q���>��_/��!D�H���n@'�q�p4�jt�� �zwC�aWv+�ๅ�]��Gx�u���'���Sׯ�8��_ʟ�\J�xtn�)���`�O��d�]�N8P
�$Ug�`� �g3��<���U�� =��{���@�����Ũ���c��c\!�.7���HQV�*{�k׳��ŎQ���Xz6���=n���T�X��p=��Hfd�#0���50��ף��9+�
�J���7$�T������������ε��I��o:�e6���_�BKvݘ�C�]a�w,wgLˈ_��� ��z٫�ܷ$u�������]uW ������Ĕc�~�ar�j�+�;����'(r������'��)>봈�:"��6��%U�6��O�{nJ��8TMe~;,���u�pe`�!��Y/����Q�='�����ؓ�O�.:��ץ�ҟ���4�Z�ysk��*�1��S���NF'�8��A(1q�\�*F�AQx~�z�~b��#5E��������	q	���t�P���LJ���_I�Y�:6���ʁQ�q� &vM��s/�[n?��L`@;�ҏ��H�5O�L4>[w���יD��Ih	���&���'�O����6�N[����0��J�n*�k"�E�B+}��'E~a�yYQ�'����uۇ8!�of���wϮi�_ޡ��о%�.lm&'!�B%�����s���#�a�Ҕ�?�a'=��;�@�:A�L�'�	
�X�
�0[��VB�>؂��<\5:]t�\�g.��F恐*V���Qwt�������?(��]	��G{L�Cں����|���g�Q��%j�XQ��B<A�{4�yK�l���5\�!>��G}ճ�$J�� �@+b��F@��|I�U�8�U?-TA����P��;[������sY$�N�/�
��V� h֕�s�����@��M����F��6͋�y�o�2���ƣ����*��z�ڊ��;�F٣�:�X5�-3��'����ų�X���F���Qf̮=$�r�,���~!0<˚�"������v��9������vu���yĬw��ǋY���ƽxc�j*�8�c�3�Q9׎�R���ػ�8Q�y[mj��N���z���5^��kΩb:���E�tQ����x ��{H�~�;�i�� D���Y͆R�����#�����:�PA*Sg�͇' ³]k��šf8#G^e��$Te'�����u�'�2/h�5z�.���dZ���{�|F8 .-��){aP��g�r��v�ɃL���{��1����M������M���c`d`-e֒r0�Qz�)�oq��(��z��3vkNF��}P�jS|Mܔ�.�]l+ga��F�;k�5
P���e�.�+�O�j���Q]��ܙK����R��!�_��&�7�'	�7^e�:U��k�Ĥ���Y���db�]l��l)�:�i�T*FL���&�tH�#��>�[J=�a���{�PL��R�J�y�v� }u�A
�;K ߯�3*�d�ЫO��Bf�cD��V%c(����E
�q�1d��u"�u�*�^�uMu�uLj�� m^w��Ӳ�T�9~�	c�H�2���_\mJ��OŮ�r�C��:8�o�>�Y$�"�ێ�Dj��h 2H�i�$��@�x<	������U��=�`�6�A�[�9�G'9�d������EmK���ޥoM�Q�_�	�o�,�%�=�����������rq+�O�Їw�S/���o�e��&܌]�� ��=G�qw�|�t��Wɺ����*W�����$��}4��{��1�"�3AhHP�t,4��������%{�Q��,i���T	��|^��t��%������of�z�V��#�,5Ġ��������*I:�,�\�˭M�����h=ƒ�f#U���F�6�e���}�`M�?&oGh7i�)�_���nsyN:{�?U��6m�wBoՉ/KrVy��ܜ���\~�W<Į�&�����l�%���Ŝ&X�OJy�U�����3��ń�m��i����T]���=g�u�r�hN��k���TؚI�,�z	 D����X����s�_ea�^�����r##�ļ>�����B2!sO�43V�k��@ک+��U����|ZPuɛ )��ґ�L=yʭ�
��2��p���aC���ښy�E0I�N��)�c����)�U���'�?`��m%w6 ;k�#Y3��$�Z�%?�dv2�ixj0|����+�ׯ�H���X��(�
'F�܎�.�e�\�F_�
[RZm�!�^Bx��Q8tCA��R���ns �O*E~���4���8��{���C��_���c��X\�ڟi���[�-j���������VD!��Ca���&�G��?��4[Tg+�BW���z|����h�.��z�I�4�ìR�_f�b��Ԁ���$˯M��]�E9��d��4	�Q]�����%?xg9c=�ط��L���b�0����k�W��ע�?���s'��,;�ߚx ~�s��[1(�b;�I׮�8  �K��Z�/���[91�GU�Fe�d��{t���D�W�b��o+�!6J�"DE���Lf#��'�@gջQ�+Ew*!��R��&��j=�6�I�͸��6���,s��?9c�J��q,?#�6�h�{d�Fy�!���n�r��?�\χ	�n]����^:�:���{���}��*�Q]L��0g�Y�/�r��bB�cZ�q�
����d����V��η�I�������Sn��#.��z.!vf�J��Y��V��uH�=��U9��b�ߒ-�c5�3��;���!Y跦g����΅؅.	�dl��\5`z��ش�����Iɕ�J�tQ�qa�I��ȶF�L�.����,�?�s0���F�4����g�{��7�!֐�L9��|�V�M��󭪈E˷!*�l�H�O�(��*v��]��+���{Ś���R�J���Cش�,�}E7�O>"�Z�9hH��/ȃ�vu0 �Sv�Bk���l�-�����ӾϾջ�ίj����[�Ek��֭s��IygG��$0�U������I=�y�xK�^�F�����:^���� b"(�Y��2+�(^��<,��a0�%ñ#]�8:��5�4^���������������2�d�#�>��#\��٪[Y��2g�2S&�/�'2G(�����q5�ˊ� @�],�%�C�t"xc�U\�o�jl���� �$�8��z&g�5��w�f&).?�G��fZm�r�'�E�ӧ7 [,SA�"lNoޝ[���n[�f���7��=�4�	�/Xc�({+�M�/�;��P��G�Hc����QaU{ޫi���1��f"Gej�Ǹzd��^�����eU࿷�f8�vMI�(���i�P�Ĝ}��:�Ʃ�
���F�TI���¤���ڗ��8�$i�Jؗ��
�����s��f�oI��T�<���і�W%����P�;-{�HMfr3�{^i��L���I�������F?��F\\WF>�[g�I�lBs�4���ݶ�����s�ʹ�Y8%(T�ﵸOl�ԟ~����1�a�`Oh�|q��}���&F��R��Ef���9�A�B��GV	uTU����ڢ��8k	C�
��`(M�ޝ�:��K;�W�ӏ��B�1������r7��"��ԗcI�wU4��7A]T�Y��T]o�\��$���	o�e9;+��p�i)S�>j�_�7	����%�<<�[�B+Ɨ�6m9�G(:��������E¨�f�)d��C��pV��3���.��	���S�J��MIb0�9RGw���]��	9s鱖����d�~wC�,����b���wP5kPk.`x�}O�b�{�ǜ��92��\�:����7*�2�.���@�gs��ɑJ>9����sLt`z��3��Ĩ���CtO[��]��u(|m:��k�\��<gB\+��>z6,�k��r����O��	�܃���_��O��!]�ͯJ�Q!���ɞ~~4W�sTlȫ޿=��e�j)����y%B(��`*�ykn���������d�x���������W�Mm5��b�H0�I@�����8@�~1�L���M=�T��4	�{n�,��K����/�����Ò<��3�?���z����fl,�Pr�Fkp/�Q��*�͵�t�#[���W���P�qc��[�9 #v0�k�l��@�]	����9z2���_����������Ф'V��Uϭ9�~��6#5/�¦z��(QYm�]R�H�
��v�7/��
��;��/��vي�+6��(�H(w��؂��������b>�ґ-���<��R�켈F��̂׭u)�t�ps��H�ڪ�дGD<�si� <7t�;/Ϟ���%Y��q��Q��\`�
̊�I�˩��h��c�\�%�P��zy$�BT�'s������LL��L�&/�[ު��K���o�P�$#B}HŰ������Y����l����vX���F��h�s��(k��ac����6KZ�^q���V���2d�g/�pcΎ�r1[�ʾ&0��o�$��Yz�AQ��>�.k�DR\��,Pz�u8�n>�&p�Y^2y8�m�^0u�
'������	J��E�1̖�׌�WyS��g��q����7�h;��M��9��/́� ��Y"�6®a����5�=��p�_��y�HYKkM�^r�FUNI��?�U��͝�˙z�X�gD8T݇�yK��Q�]��mzA���r�j�t´,�v{w�!�I���i/�'��m)W�m���}�
��
��׳YJ���'�3�M��v�軬=�5:���Q�U�R��Q��A���(��[��s�M�	H=v{B �FW�w+t�۬�Rh�6*��z���	f��3�Wng*���Ym׬Q���#���|x��Δ�33�$�2yEk�t$t��ɡ���>���d��jZe#O��Y�"�\̺�4��o0�YQ�I�8��	c��� �`��.��K?��=�������œa�4���Q����嚪���������~�x��+}�nҮ�AI6�O�*�O��f]*��r�N��Mhy1�xA`��9i)$k��"7it�y�5�:�ЧgA?�{�k����B��m�:�![x�}j.o�V�mC[�pՑ��0y.�(��OuS��tO�Y�Gb(�(H 38�&k9
������*d�=^�(�� R��Z5�x4u�B�f�/MN��}�O�l]R6�Խ���^LSc`^P�r���w�o
��7�2�`��kG����#�VΙ��z�o��_��T3vD<f�p��5���k'�8�~�Ơ���i8wʥ�ps�+�3�J΋��ѩQ�z+�X�ԜA2�G��� q�p�ݯŧ��`�M��s5]�YÖ$�%h)�Nܿ�����J�.������Ml�)Z���n��s#n���3�V�V��� ��~1�M�\�.�9l)���Y�~'�hsA��A�������`�{ϫd]F!۶�^i��S$1*�$�&��9IC�����k���O�)l�H�͊QB	@�6D�� ^�N��6kS(�*�����h���g��V⑬�5��E��$@����ac>���-}K��=PN����楖�O�3s_�'���@ ������$���5�QzA��0�EZ�d6s(��9���Õ��W�*-�&<���)nO����W�jޓ�� ��"zMxJ��YW<��DN�ke�@���"& �>n�е���#���-cɖ� �|R��	���=�Y��ڿ&����WmĆ���j�ˑ`y���w)�F[�/#�n����]s5D�xA ��풯];"̃�lup��^�+�����=�)h�����2ew��-�Q��m��*S��e��n��-BO/�뾪E5�P��gQK���}��-#hH�
������2��jF	�K�h�
��t��� (W��G�Ԃ����Ǔ2�`��7e
%Bi����Y�NköqH�%����
�|y[q2�[��V�#]�^.���r��}���?����9<?/c���n4�U�͑�E8K��7i�����$O�m���N��p���)�e�I���K�0�S�'�P�\0M�9GدJM���k���ث̝J�e�����E�B�����ܻZY�Ӗ��*^��P>��UAb�����}\�R�d�v�u,�P���4���G��3�X��._0����,N�����Z��J�}ͺ�iÃ�㐎fN
p�3ށ��{�M�r$��+ $J� ���ͱ�D3��C3��]'M�������P6V�ދ|�0�<̡�ɉ wf2^�[��n�RD�.���=��儾���V�����
e����eP̙"���Z�!1����Wk��<XA�3]`+c���Z��t�3��>lփ�˱
��&1䛷�%�Rb\��<蕇����M�y�.r��l��b� ���B�*�S�a���N���&V!�܏�yT#���M��F�t�̇̒�E�+�+Q�J��z)��`��S�r�)��)�
�ʇ���H�KA�(���Z�rHz�O�r�Z����IK�����>��E��<x۪�9���������B���')��= g��^��{��d��"�n!	��"0C��L�K�T�%v1���̅�h͒Y���M���GJW�Y^o ��o�����oC/��e���
�ҘJ~��D��{��W����n~X������Zp�$�m�V��̢w�ʄķ�m�7�&�\)�/�ƛXC�W\7O�u�/-��|�%s���/i�r?���8k!�D�r���H�`�ya��)$c����������kG��c��1� ��?�;����l�gU큤�q���H�*4f�x^'ib������u^�G�)i��Pp�!�.���屰il��0�s\uI�������L�h ֗ r#]��2�LsuCۡ��gB��^��5��	8�Ƶ��*��}�)fMSq���лn�2����%�b�|X�uP1s�yM9��h4��.2B.�	�7����h��u�E����TB��C)Z`:Յ���Qslq�<^�E?s\�:���:}�נ���B�`Mk��]�4ܜ�#s� �Sν�!&q\�w��D_�
m�v��	u�=�}1���Z�M�����yj���2z?��h?����T �#���ކ�m+#��G� ��_W�ebXt{��w~�P�Lp�ԑ�����Y��xv�'y��6�0�N��I�W����s������ܠ܄ ��12�9g5�A���i���l�H�O����O^6�ʕ�7�ț3�a3�z頢mQ6J�v���y�!�Uc`?AmPZ5u���
3%g�IhrM���(uiB'i��$���9������9r�QQ���Ea�#�,7��J9@����s?-��R��S�[`��xq��dZ>��� aI�G�J���d����fDS����9��� �5m^~�B(�-�_�p��#QG�n�:��R����W5w�'��ь|���j����'-�Ք�����Q�������⓳4��g2ʆ��r�%<��������m��yнI�떩\iqg� ZiH$p�h�~��oQ�V�b(J$^$s�z8�S����.x��m�h ��5��VDrn�1��ixoӌ��Ǧ�����ԯ|
9�Tz����|������3���w��Bl��LN�뵘����ׇ�Ͼ�3�°V�FA�h�n
�5�[D�>�%�0c9Q����Oy��gS��Nt����T.�i�Oo{�պ	�1b~�a���j���/��M*��]��Sp�Sյ�F�F­��%]8���v��N�4�ې��~C�b1�ԝ�K	���4�	@q*�e�ڼvB*P��(	T'�6��R7��KyBӜM�Ehz$�1�����&����r�t�2g��n��Uiu�e�Z�}Ko#K�\����$7c��5��q�r'��4[D��u����G�"C�,i��gF�aMp'�&�S`'�a���>;x��[%�З?�L��(��4�L)�j���`�23D�����6�-�ˤ�A�y��=<h�N��,�Ҧ/n��A~�'Sï�=����,[Ķɱ�m 6�K�Xٞ  �K[�U�����r����$���y��-�V��:lIm�h�z�m�o֙�@#���C�2��j����O�%�xz ?�az��3Oݶ��
�q;\�Z�1mսU�j5���t��'�W����;�iM��ě�DTiI��#��}��3��Tٞ�_��*��G�Z辁�R�ľ�*�7��{��ߢ�������L���Vm�M0u1Å��u�8���3�D�#i��#�7�Gh���_e�����1�q�*�ykV=;�kO|�XFcՠt�N���֢t���Wc��h���2��dN��� $���\��b���ڛ��d0����$y�$t�������x:q��[S�ۛ)�/�l��D��d6>7S���~B	�K����"�"]uUà��$tI���k�W���{�����|k�B��������3�5R;F� ,���V)��?�hߧ�gH���0<O��Щ�H5��!��^ø��z.����˰�	v�P)���1�q��uGYJ�nȍ j7Z��s9�D>2��*�����Sگ䝙�֗<*��9s�\a�̟�I�V��"�Õ��s/�Z�U�>���A7��Ӄ��3S�%鑼�O[^Nx��+�Q@����,�_������ s�2GB*�Q�:���öueDl�:�,/D	����Av���VK�55�����_D�7&��c��^w��N���MQ�u�>��R���m:����p[�Z��!ߥt��!$��M\ȷ�t�<;a�>^Qi�y�IĤ|�q��`�zeκ8e9�����Z�*��Dep_��tҝE�;Sp&����"�/��sx��Z�}�r'��Xm��[�\���/wǤ���z+�j������e�:&ޮ��:��j_߈vr'6a-W�s&T 8��"��O��N�g������W��i��5{~0ܢ�4��E���KTb��RB�2��s�d.�qG�D��~��eHXve@5�Ty�̝�q65�ж2�`+�f��"rfR��W��<�޷!���u&�wI�2Ӗ�h|#��0O�҄���ե����?�����s׈��]�, 5�h�@�񤃼_�5�D-���ܯMŞ}��5PqT.����Nl{p^�N�ρ�+*]ߔ^�8��:D�8Ж���|�@4���s�\ߕ�Q(����i|�[zτ��A�/�O̾�nfb�k�k�\��5�3�̦���$��l��z�F`�t1�7�8��$��2|!C��p7`�č��;��fy��(h�ݭ�p3`��w��گ��G�dxM��(x<��8���yz�j��\+�jg�{~m<�2�M{�?�3�>%�9�9㳿���-zM��W��mI��sg|Ks�Bُ�&TX�)�9
�yU�` �»��N) F���G��0Um �i��Y���;�@���c�18�e?�۾0��Q?|Jg���"��y�9W]�����=���?=��[��-F\�j7�ɯR��PSď�
��!��������������Qś�X얕 �)��Ē@�-�!�]� ��4X�����5����/27{�ǳά�'�Ȏ׎_3.|H��S�����sN� �D&/��G��u��0U�fŻρ���h���vA����B�uV.J����4%���s��f����ƛ^�١e]uX��.�%��}��#y�;F�݅~���qx�{������3��b����6�)�.=��*����K�KoZ������c��04g��u$�n��s�5��XJ%�~�w*o֋L��3����j�[o'�W�o�P�?=��_�1���I��Adw�Z%��J����V5#T��F>Ѯ��<�g:����$�p}54%!�y$I�(}lnhG#y^�,����Pt�%�������G<��9���
����^�4��!:DR�2�Z����G�P���q�BGjrG�ϑJɦ�=�	֙�@\~
E�����*?<� ���s�"r7uXEt}r����������؆���DW�>@���f�`ig��NGj$El*�Ǉ7s��c��RP34[�롯c��<z�<
����-��s����!�꣰ɜGL������}Kz�zg�/��k��p��x��� {��/��zO�tV���{��o}׵��KΞ� ��i�	j���X��/3}�1fY*S}Ǜ�y��x�xbv���IBs"8�R>�bp^ms��JQ�r^q�Vo�h:���݁ /���Q��G|��zs�W��E�g��k���Hl���V�8��}�f��?Ų��Q��=�V,C�Vҗ���E��r�J_Z;���=��t��($T�I� 2�ٹ}��|����'��4��$#
�1EȀw R�+��4s���?�ib��l�I���Pm[E��	]1�,@�#/��9<D��@3��yx���%؍A-e4�[}�o��|������ez��z�ER1�x�IDv���>�Z�\44�-�S�4$�kT��D?U�i�r�8��|<�dT�;!~d�Ҥ���7mT�6g��*hD�|��ͻ��A���L�H�s��8}	�8��"�t/��;#Kl���nu^ͤ�-ks11Ԣ�%@���`:6��� ��v�{�D����\�\�s�'��E:�(�݇�Kģ}��G�1��c�{���5˺��R逦%ȵ��D�;~՝��3����P/��t7����?���-��Y�5�
-9C0��z��"�(�4�#X|�#��4���� �1�v� A�A�� .�M�c���
j�t���F�p
���}B���R5�{c�b�{�N5v��!|��*������4�=y4�Y������,��<(����"�kg�Z����g�.��5vm=Fk�>Wf����kC1_˽,xb��K�4�_�x�@���&@��A�}K]EX(\*a���yR���8����w�9u�t⳴m`8�gZZ�؃�9�Lމ]��Ar��8|.Sey��T��f
����a���&���N���.�Ƨ��tL09Tߟ'�����g��ug<�����FֺoH��5�A���;���F�lR�8�SU�}�9����@���t;�59�^�F����m{yTs�r����$��=�}2���ű��#���b�5e�p7���f%2Dz�/'�<1�Im �0NE·Y�M2�QH܈e`���L��s��u^��F�{4j�#=��wjLc	F)�JJZ��������:ۡ�:c�C]��J	��&�[e��@A�h=xb��Oq�ԅrj�dh~}��\��Ƅ��郇��`����g��1]��~��T��'ɍW�fˑ�-&SEl���@� פ���F�>i���e7���9���F�&n��9�F��m�H�#�4���? _Ҕ��T�3+��^�?-������INwx1�$���y���H�?v��3����ҽs��m����̺͎[���������������u��>S����R�j9!��zµ�=��*�C�}^��uC+�I��d+�)&�$NC(i#>*Ӧm��k��d�Y'��,*����9�0K!�����'�b&Y������7p�X�Q��Y2vcL�߹�\Y�	9��b��6��v�ڮ+�Z�E�ft�U��3{�V+��P�L�L��ƖMʖ�o�)�H�Sj��%Ux��\O�!+nI��9�c�A5�������\-�n?��̴�+�w�-n�dx
(i[�������WE;�Yљ�1�����\L��T��D`���E�f�5T\�\�Se�)�iTcU��L�����$�J�v���%����Z�!�D�./ՑG�L��axR�m����W���v�,z�݊v��J���zfn'�a��o|/��}�^Wkb�)��b������ж����|��:�@���-�4b�����MVX2�SP�<������E˪��OP�##^�9禎4���h���k�|U�A�v�"�]�x��h��d�3	�iB��F�K�3m�^�0{h��A�%���\.Lm�,�*��2�x���|�S�;v[:e���o�sk�\�Dk�j_��V���x�`�7-;�rWl#�C���]�=Q�E���h�6��	PA���F�����՛��o-�@p =���)+��2`����N�7���)��F��Է�����hSND�hPy��|ˁH���C���MБ���d���R�������9����!������\���?mΧ�n"s/��)�����xg8�X8��<���p,?~(`�e�vΌt�N��Tm�ح���(��0E�ЬD��c��Z��m���M�4ˌ$L��k�>o�|��"m?�3"���w����ǥteЖ+e�6��;���Cƥ!��G��G叒U�M:�(!�'�6�5�bm0�v�6Ҝ����#��2�yZ�,rv�Al��H#<g[���o�"��^���S!��oCl4��|v�N uX\'�o���7#ʉ���%�fB`󎟉�?��|��_�8�Y�������-u�}R\���:k�Q$��`�ϋ�((+��"���2�FHQ>�+Y��Xr�z�9����9��\�]�Mw��- �bn=����i.�"�/S��U7���"���Ԟd���7SE��
o�R'S��&��	ފ=kHo����	�2��-t�c�5���Z��k�m�	/�ȝ$�E1n���K�U0̠P�s�	m�3�0�x§�L�7�b���V��?�߽X��&����#jK#_HT~�I���.�w&�Ą�! ݫ��5��������b;�ی"B@��q��t����HD�iU�/i;�hsL�!R˙�n��
�Z����Ӆ�q|����о�p�z�	5���QH�￰䉘���L�T��juFi*���)S�FE�ns,N���+�>�q���~��cO���b������&J�o�O�)舜#��$�Ѝ��c0��?�m�Jw��t�|�.C0��|:�����(��8m�綶�yB�@��9L��0d�H�`��C<�oi
mz	U�r[��T!#��PP�Em�l
y퀍W����mI�p��f�ui�f��Svۡq��q��n������h�)����i�6;{��ϧEP�]#)�0)F�_�����c�:���g|H��%nP�Q�??���mc41������{VT��,�[��V5�AP�����O/K�����Rw!^�_6�fJ%�ϕ��h���̷B�v�E���c�����P息�R%�_�_��o�6or�A�z?�n�s��˯QVo�Nn�R�V�h�,L�RS�[U7ڃ<��c�Go���fW\6��ɪ���/xM|�0��py�<�,�8��~��2��(ܞC]�P3���FO3 �����Z�X�/̴�����0|9�h(�ѕ��eФy�S�21 W`$.�fj�~*�n���\�o̼gC^��)t���Zs��T	)ð��,�LZ�#��ts�٥@�Ti���t�Mj�ч�V���e���5?��\�؍�]�|��Cø�K*�ٛ�$��]�`���`��@�2j?5�ץ�q����:������i%��1������a���{�t����}&�^Zp��4�gp!#z*0c�Ǚ��[�>@�ޡ�oKL��b��@c1)O�����nO7*=A��a���&#���_Lt�<�.<o�S��*)k�T����-�P����1�3��o�U�G���zı	���{@)�>F���EM�wR��&(jƃF�c�� �H��G����HbmLW��dbrjr���X�=�eɃh�������d��Q���ϊ�~��`�هJ��4��+��<̨d	q0K#-K�y�k݆Y/���d���~�(w��1I����ӛ���y}�Wy$��U�oPWk�^0b�=-q4�#�g����ޟ���kEX���V=�y�D�S�Px ���dR�A���*vP�4�Vc��M�}V��/��"��<Ы����O��c��/Ƹ��m5A����
>�%ח#�dFK�j��ҳ Yd���m�H���6`īZ�l�wF-1|x��Zm��_�|<[X=W	_
�|�~�)yy�WHΖ�����7am��7	�[�����׆�y2��X�]�<�
VO�^���O%�04�; @�J�rXL�4a�m�[Z9-�S�Iɝ�n�.H�AJ��Ħa�߿��b�jt�xʛ�eJ�6hgϴn��g���Ӯ��NB$��=�f+2옡 �E�}l=4�М�QX�;!�P`8���1���l�p��aO!d������ E5���Z�~�1㫫@��	�^u���)�x>��y9���t�=�b6���{��/�g�w̨|��&�Dߜ�s�B߇Ws]߁�D������芤ՙ�����/��Me�s_N�٫�rV��ݢ>�ViG�����	�|m ��[�|Rv���Ԡ��<A�.3oǒz��%}�?`���EF�|mw��D�%mm��ߐ]o3EC�L�`�q�z��r��gӿ¼�!s���1:6���U��w��9�z��"�\���A�m�F��&�f��O����k�?�8|���n��H���B�D>t���	��v��3����U�[�UX�%g��� t9Z6�&K6�ò��/�|�.��z1=qq�2n�Y<�����$N�{�d�ĵ���Q �����)�'�s�B�FF6��?{빬~�*��	��.��
#�e�F�fEf'����|�8���+�]�R0|���n��p�XDt��.]O��k+�A�I[�-���<vI�����ҏ��݈742�JC2:�Ͻ���6��-�����[��}�K��N�,��MjA�A5'�e�c�S)7��t�%@��t�3�U¦/y���?ye�iO�3#y�W������$�u��q2��Hy"A,���`<�W,Ypʝ�Ax��)�n�����iM�۾y�Vf��֮wʷ�=��\�"����Rj�ٰZ�C@B�pX3�kM�Ou�7�і�����u��~�
Q�]��e֐�i �@�H=H���u���5Yd�He��CĎ]5K]���X��Q�����\I<�9g��Q�cT���D�Z��>�}�� >�E0�FȝTZA�zy��L�3�,���g�L�X���袝ՐR��h=�"p|���` ��~}��><t�}t�7\U?ڳ��P�l���Xi� Oj���,�L=J�&�I+4n��~]jV�\�6�*$�Q߃bFF3?gEn�m� :�f�0��c���E!А3m����z�*R���Y����A1G�7?1��ofF����C?�Ij,�p��M�fr7���ո�a]���M�?)�oX0S���8K53��3���އ�b&�X�1�����;��*� T���ΟKX�x=�*'��qO,������6��X������u	��ri�t�Љ��
��{��敄��AUI;��w�x���o�3�M��?Qpuأ��I��lzC�kH)ӣk/#��=*F��� X��ظ���4���rݢ��3�U/R9ZN*�O��צ�kv2gA-W�_�4�ʣ=y�}��_M���Z'_P���C�Y_IYl'��Yp������zlފW����mN��滀m/��v���<S�
�B]FGp�t��l{\�8���r�{��km�������K{� ɭ5K p
�o��TJ~���{���A��t/��@����q *�����?Z2�9I�-��g�6���)�1����
bY�.y�����Q��&4)�U�4d�E����W�8`��BF�/�넂c=p[�&�/�!��feK�� �6�C��P�\�O�NB�R��ݡ�����K��]��/���l�4�CO;dq��DR��j?M��By�`������l���Ӈ�C�wF	mO�X4�F<6���v!E���&R6��}�����\��~�F����hJ呙Xish�F����;�hgyA) �7�80Y@�����c/�[�-dn|�)��](�r�`�]J�n8�Gm�K�5U�\:��Bp��jH���2��=�Ԑ�f��Q�N2�[����:���pƿf	+0_�2 �c
��r�\�X�m`���:LN�����4��ե���{��h��Q�����e.�����}:N�s4��do��@鵟bW���P�����C�ՈpV	_������2WT�(�K�a�5�I��X���V|�+�{|dd���Y��j�,�����#��ZC�훮X=���oWG��x��f�Nk"����<�c�&��6�8�K[�D�Oh�3�4Q��6k��k��h�9OkA��eM��֠i�Z��BQ)�����/��c���y܃Ӛ�7�m^�����ڡ !�K㋎Y��!�3�	�O"JU%�ҋ�~	vp�s�E�ڱt�)�X�<"*�Xf�M���L'��d��: Ā���1�eq������>���tGJ��Ϣu�xhђ��;�vf��0��:�}�n�g%\L�6:�@˭K�@n�C��o�\Z�9�K��u'��9�e+dj#��7��jnJ�}��S�]NU�~&�����l��0~�IO|7��{�'��V����!�oY�<f��FL���f}FB����_�Ϳ9��J�E���`����V�� Խ�SJ���+�����������b)$�@� n��Ԕ��1v�`^D���)��f�j�W����WRL�!0w���a�9P3���Y�a7+a��)�|c'���^T��� ���w�J@RƼv	x�����F�������~܅.�uc�S,Se�I��&d��SVA��M#/�$#�K�yMEG�m�������,jM�xnem��JX��	L׉H/��h���f�o���#��m�{g�P_����N�� ��ۭ��~���9�A9�kbVh��U�3��^����fJ>�5�n�j���a����Ӿ-w�I����Í�v�Qg�s�ț�Ͼi	s���G:��F�]Y�%���9�'�H yN~�l-��ו���cx�������Y���Haڟ� N���:)Q�R�y4u�CМs��>_�e��F��k�b�sA�9�9ٌ�w�|A��|d�u�y�Դ�V�r�o'm�,�,Ss|��C{'�ѯ�{��+h�2�,�,�Ri�wk��",h��Y�S�:ro��:k�#��^��C���D�NbR�9x�{�w��{�#��|B�����ĵ��@YO�q(�n6䨠o�ޗ{6a�'�n���,ק��1=\^	 h����0Brh ����;H�
Q]���HЙ��շ)�P�j���{��=�P>�_��h�J���Ѫ�AzRw��e�"R��Z��l<�=�	�I#� mZ�D�h[�{���n�#�?�9"�N>�J2������e��NEtET�VܿRF�#nt�#&�q�Y�2{-U�hcZƶ �-I%��w�����j^�̺+7E�o���]A�$���pdҒ�D;Kur���M�� ���l��񼷡���Q�P΀^�ু9������}�,�48�pT���K~0:Q������Kۻ�E��vi�&O*}
��-7���}�PU_�yO��N?�k�`�S��	bnN,�T�Y C�z�>��Cc,Og�s����,����������C����S�u�a�9
�-�L��xօ�\����*Q a����'H)���V~j��R�t����Z��m�9��Q'f7�d'�#3����w�FdT֬(�_`w\��K��rq��ץ���/)��<�s)*���!���{-�1ƭ]���s1i^
�E3b�y�<���$� ��{���ǝ7f�|إ��Sh���!��"��Sj�o*Ӱ� O�-q�0��պBZw̘�JO����6�p�nUN�}w�ȧ�\���R����U����Һ��ǔ�����Ř�m���Z��ex	i3Â�a-ϔ�7���� +��*���?:�B�����V}�۸�W��Xa�mT� \��7��@��'���d�8�ve�����VC��%�1�ACƙ��ȚWg���u쪖���D
ǰM�ө��zB<�z�hW��j֝a����:J�kzO�bS�it����XQ�ZN>�ϐ��Cו3�f<'���n�RclK\���J�(��Q��xB�޲���_��ЙN�|�!��S� ƶ�[z  �K#��i(����p~�@��9�<��K$<r�T�&>�
�tK/�u������M��b��\�v|�|���݉n��ڇ��=mQ�7���j,A?�p[j�u8<h����1ȔH2Q	�F�>����+3Β�%�ۢ��*n�3�щin-/Y0�Q"�ũ;�U��ɕ�j.��������4�F�_d�K�rڛ���S)�N��%��Ȗ�0%V0��ö(�3l���	��*Pp1�,an���WpI�nFy��A��a ��\��7�}M7_ɝѲ��r�t���n���>�C�C;�r���EΞA���7R�܍��(J�#x�ky�򌡅��JgT�>���z�`�K��ÙwV�R�w�Z;�8�v^�R3�5i	U|�`b��?�)l��Y�1�
�I�
��^�h�Σ�yB퉦��d�����S�G�Y��/�t!m�����$�y�S�Έ�Bg�
��� ���$0���Z��IG�/C �z����J{k~4c&��.7mImz� C�5\JgM���o�q������{8�y@	�ۯ��kM��=����y�:N�X���M�Z`�I�R��i���̠SK����Q��#qU����$A����^�lG��D�4�8�ٻO���X��W��K�,���tڝi�~eO��}7�������E�_K�lb஧��_?�U����F��'����U��)�?�͝����Z��,i>��Kqͫ�s^p��7�4�QEK���`�g��N`֫" �d�� �v�|��C%�TG�X�I�*0�w�~sŇ.]f���r7��eih�Hrx�/�)X�I����X�+Z6I����� �zN�B�R�AH&ʴ��E)>m�]�:��$#6�qg#A�kZI3:��'�v�i���~�j��o
���dA��-�C@���H���������ޘ�e4���h�l�<���p]ւۯu���A\8��s.��������/b��l_�Za9n�훡5��K��7]�)�Ó�8\�ͯ�����a��j��].�
��s��"���%��G��n�`V{̞���-nX�L�;i�U�|ay��!�ذld����c��]գEg�j�֣�s���q�\�mФ�Y`ʟ)UAp��t���I�a��{���5��\#@�d�������\����}��|x�ʆ��ˣY�D�c+�R�w�)M���Mkʌ2F���qM�#ő&���JR���5�w�tHi�?O*�~��b)�/��5������no^���u��*er�۰tlSw`+����l�_u=V+ rYŘw2isZ�l��D������*�T���R[�,F}���C��}�o�hCմ�G'�2S�XvO\u����k��6�9w�3�z��q ���;�1vi�ȋ����� �P2�;Uh6s¢�Ρެ�2299��?��m�]X�*U��T�a3)9B�����/�BJ�h�Y(�i-��E9ϰ^OIr9|�]�fޢz�?񾵈UT�+4���~U�>��b;m�z�l[����̃ium(���N�4>�J<:4>�ټ��ea_��2B�	�Kk
@�iD��'�r�U�����.ڔS��>}5���NBT)�������wy� M��A�J�6,��h�'],T��ձĔBB��9�X�*g���*��1͢ҁ�bg)�}ȥk���A��d.^s`��%�>�mBR;����u:�.EףE���_��u��X�3<ܗݡ���|�����#/�}�w/Yc�/��>^\)11r��H?E�zSV�$�ALi�x�к:�g�ږ���U�5ֿ�p4�wQ:�pS<[p�.%),��Lm�>�L;�X�*�^�_$��/��J���¶�I?WU��s /C9b����:�N���c�u�(lbi.�� ��hl3ɲ�_�&�jő,qZ&�Q������Q���Ş��2Ɣս�k���x�����)"����;N�ϲ�+��?%�Q1d�+dB��p�J�� �2���������)��G�t�&"_��Ik�ož�����r:'�[2blǧ�H&?��nH)��E4[��±I���U�~�ف$7�5�Xg�-
�iC�`�G�S�%!e�Ȏ��?��4"���gT���A��Z`؅����(��8r�b`ye������nƵ�s���w6��5r�(ه��� �qn�"	|
�k������H�����6{jވ:�B��D��7Y0�� �����}�U�F�@�F=2-��rѷ����j�5{��Q���r$3�<l˩XM`*Cۈ�4$�G�~8E�ET��<�8�`N_T��Tk5Y�NN�<5��f|���o_�C`r�g��"�J���n0wtþ�eO��� �E¬�ˀn�|H�y$��+XCê�whQ�tB���9���e�<��ͱ���)�.��� ~�� �Cw�TAHa�����pY�-�k("�`�m��=.�������aXY����^@D�v���7���=����a~,����H��5��� ��71.UW^���(�Z�$�.��!d��凫��=X֞��@ư��ðF� +"�,��?ֹoM�M3�"������^�=�ݛl�B9�eo��3���(<����,�4���6e��sfP<s������Pxu ��2��Ew�=���)[��]�.���<�Wkp�@C����^.t0�~�E���5���~�ȴ%~F�p7<��g�{;d86���D4 ��!�u��|P��{d.��5?a�9ٹ��Leێ�I����rVO$�Lm�N�' �9�v�#� �����|y$	d���r�P������P���d�C�;ܪW ޴X�|�3UB�\�� ���O��ƬA��7BŁ�T
>Y=�w����ː�H���5�K9dE�<���Rf�B�A69�Y�.K�s�T��x�ό��{�Nw��'&�w>2A�#��Y� �Hi	_�9Wz#G��?`UMy��km˦o���z�nY9���Y�����`J\���v�-x>c=�o�D'�Ģ���6<�zF�����u�n4,zVU��X.�)��q�j���;���>�EL"N$Nj�&�6E�.��{���6��/����aP��;�<�*����Њg'�5j����5�M��S<D:�٢��k� �s<̦C"����&�dS:���:��F�Z3���ݸ�h^ Ow�^+}(6���#�CCρ�����z�'k?F[ň�+��>�O/�}dA�6h���3I�c�� ��e��0�|�p���C�*�A��-K��I��@�?Μ�4�bD�Gl�I����eM}��:p�7�L�����WRsU����;��� �G�������Г��V�Gzk��-W�������y�j-�q��z=N=���Tu��b�����ƓJ��*z$D��aykS[�Vo��Rb<�"ɾC�����1}����V��=Lq���:�4�)��ֆWj 
�_0Z}���fD���?�g�}�5�q�]7[{�����F�sI�c��ĆC#:�şPϲ�g�(J�)�Yܔ��2y��"xbq=68�!~�*n�{ɐB����K�ַ�ݏx���b��=h=n�J��e}�+�o�˒&͈�W{?h1~�
��djj�1��X���v1w��k3$�1�㭰�'�Q炐W��~���
j� zY���ޢ�7JA��`����փ�K���dG��jz���g��8���N��pCXꙉ��pi�5S2���Y�� ��^fU�_�.�C��?���n��\)���Ē���2�J�D���"�td/?%n�JS��h�pSx���~2��0�g 7tG�ٙo�S X�X㥛7
�܅tT�5N��&��h�����������W�l6Bv�d)�s�gk܊�5��VaJ膞 x��DYk1�B� y�/G����>��"D_֚[��І'�v�x$p��p�c�7ċT����7�ė��2eEAB�B�y�$�9#9x�i�(b�t���D}}�{u���a�Xx� �$�-r���.2���@1#s�0Q���Z���"�g':-�}Z��*^��s�w���cD)ܢ�턶�V���,�o���V�MQ	0���N���s�����H(i#\;8t��j��L>Y0�-޾N��ʎ�
���dg�P��z�z���on\�a�z���v�.��h~X�L���F�v�;�����$�W߭f}�>cv�ﳠ~bvS��N��D�����@ͮ��b6��G��B�1_4��
��_-,�P\�`K����?A�)��|�oOv��K]��H��n��_�<y���m/Vv�9L1�b90y�sL8��S /_M�I4���T� ����#��Z2�<�|��CcQ�_��C�z(���lhݶ��ѕȋ����o�I�hHI6�k�9�-��)h���6Z'R���Y��Z�����jxήU�� ���5����D����T��3������i���Z `�5��9�����i��>]Ռ�Ȣ�l��y
��hc�p�,�s�܄����6�v+����d��1dN�VV퐾�~_��]\krM�Ȇ=��6��NU�d����,&� �٬)��'�8VV'��##߀��� 6�����������J�m�~�l	>�P�t��4
����<��{�46?ۄFw�z:N�_�M踱�Y����{�ZK{�n�[�+��,(��.��hqh ���.7��BgB30��~��d����}ۊ?�幃�r'��J��Ha�5B0_ȅ�ɛ�ύk� �%���`��̥i�Xr��~\g�/s��\��jy�
�f�ɴk<T��[�)V�'5NAE炘I�.k,������X�r5o�,,-�,2�i� L
;��f�Q�}��1᪌mƵ&Q_�6�ߔ�3�o��(F�E�j����UF��* ��8�B(�FqmZU�?~�~JU@9���;|���^�	�*���(:R=�H���D4���_�Q�Y`��''6������ ��A��ܨOls�3
�����Rߢ���C�Ӯ7��fk^����`��C�*3�%gRvV�s����@���7m5w�P���d�';�Ä�&,O��.4�Z԰�i��o�u�_$C/yl$@N<OBj�����U �$�t�K3�Wp%�1)�Q����<Sc���~vl�=��7����$�
�ߓ3����v�&Ǻ�N�o�&Ft���-�[@GNh���C��QH�JBF)�� >�����n,��'Z��G�k��Ӟ�&�`jQ��X�l��O�&�{�_�2�L��*ה�е�`�i� �td
��ƨP]�)�BD&�Ok��_��v�,'�܁1��dH��U&ѵ��:dc/���j�q�;�z�[|����J�x���*���EaqA�����X4��摀2��%~��Ƿf$/�6���^�d��Ið)FV�p��2��rA�ǩ�wy����Q)o�I�Mv)�+g>��i֋�tJ2�f0�jV_Y��D!����*A���ʡ���Aɣj �bn,)�&�n�^� >2�{N��!�x�Q�g��j�����)�"��e)� ���q	W��fd����E�]��^�$�5st0�T�ގx�����֨�\5(�[��l�\�`���oR���=P�A�(i�����X7ƫ���O���t)1W#bf�P���k��M��T�у��擟�����V+uF��C|Q�'�����ݦ@��a[�$�:��0S^�oumZc�7�����r�^^1Bu���/���P�JH��N3b~ɉ�`�Q��>�|��1�}p
c$UWߍ��A�H�h��w{O�F������8=�>$�L��]��X��]�ƋE�KA��]F��%u,�4w�}�з��;���V)��@�o-���V�I�@5?���@HY���m�/��mǉ�C�����(�'䕛
��VB�����ٽJ6Θ��Y��S�R=���W}��8{�}��nuC-[�	�y9.�������52P7ַ�<ü����<����l/е�����ST�L����U�`?%�|^��k�*�l�/�ܶ�g5�ܑ[��k�.�#���AcJ��iex����d��)@�l�i-��y��`�.�֧H>��<�G�S�RM��5�>�r�(�@���w�3϶� IL�g�<qw�t�j��Qv![݅�y����<��u�[8.d�NǤ#:�M^;aׁ[�	���^t�T�yNz����Zs�h�e(��涶��#�=u.5��W�E�V��k:y{�h$�I��/uN6��;Nk�Os��qQ�G�\~���2�刋�o��*ɂ�6�Qg�Tj�gw�$�	�7_���i1t2��oj����� ���br0nN	?��/������T��|��̦�D�JG�����3�]�:�S4�g��"Sbu�s������8mY��k���%o�//�5P�q-���k�X�v�s=�p��!;��$}�� 4v��2I�����*/��7lO
t����2�&a��b�6�R�'ǫY,q!>��	N:*�VA�W���L_�g���y朒�?�D>)����X�Ll��'���G4�r� ��i;��س�M�u{�0�?���Q������lꇥߡǸ��I�u�m���1�a��%8��InF�"I%����Ι��Mu"����ER��L��p���Rާ��0��(@�^��o� cc�%{�Aw(l8��a>�4���)cвe�Bgg�I�6�rI��}퍂��ek��uN���+��x�K�d�f���AKs[ ��E�����$�	�
Ȩ?�kyR��2��k��L��rm���w������uX��L-r�Q�*LS.U2������؀O��y�S^�Q�2c�k��V�e���	���EG[�w�Lg׈� �P�PdR��gʍp >_�.���~�!Kº-��E��8�|��j�7%�� �W0�Iݙ�E���A��ؠ�K]�ɩT{|��}���B5�������!�9b�<���d��4�(�g枯�!
E�۰�0������� S��W��J���
X�POD,��/G�nj��}�t�Ns��ֻ�w��N�Dp)�3��I�A&��7��sp�Lk��I����TB *Z�+����f��S��I<4��Cf�I����Ww����0]~	w۟��� �D��.���6���޺V6�M�?�]oU���o���6M�r�LcR��ּhv��t�U2��@8�^9��9t����ʥ��a?2p�
�ʎ�gH�D����}�	6\������ֽ�;|d	�)�Twf4����5�(�޸�;I__��]}��~����,f��;Atq���q��V�Ƌ ��),'i P�3m�H(�E�W.���4�HiȈ-�	��_�j�vB.7���^�!�q�ba��Gs����0j���̸������ek��8T��fC���~���\ ���P6^<��@�f=�)�U�#� �e�GP�ն}p���%�Y������<��<��`V��r� ����K���
�3-dUg�w�Ҽ��"{�������a6_!r_�u����V�Fj����3?���ҡ��k~���@��Xd�iyf��9:���2�]����p��O������#�����1�g�Q��Tjs�,�bȟ����G�T���f(�n(f0�p%r�ȗ0��d}E�2�z����L��e���i���WM��㧺2-��p����'u���c|Q�*y�C��Cx츢�,��P����}l?(��j�V�!��?(!?}I %����ԇ�����	/n�Gܬ~��E������j?��8�/���<�tWZ�L%��9�*+0oQ�-nr�H����an{Y+�>k���D�m<4��7X~b���L?�nA,�F��1�gV������� �6��ޏu������ΫLp�^	����%���./�M�����W�_T���I26r����h��d3~�>������������ԢZ
�/QCd�j)_��"��At������5]m���"���GF�33�rrwT��ʍ�a6 ��MmC����l�Ӿ\�ӛc饧A�]��흞]<��͊t�o�4������3aA����jv��j����ė�p����*<��T�]Cv���2��y��1�۩07�n��yEjbwf�4q��P��]fH_1;,yb�3m�Xj�>�8����a}ܞ���˞�
ӛ{�V;�3�uA�.�r7�q-����-�D8���8Q��=v�YY��~q��{��%p�a��� �U
:��Iv{����Bt�L���1��)X�]�V����'늆�k�Y��>�Hµfj�'�m0���t�B���z���n�X9L�>���� �mu���5�"kh�,��&�%7�WD�Y�j1�M����󕋤,�XF<jw����{������j`/f8ؒ�f�B�l���7L4}-!�zi�S�e���²�9_�Hp�a��I��潦��sǻ��L�0G`F<�����ߣ�Sb$������|���zAEM;����8���G#�����Qa�
?��OF+�c�žc5|����~8ͼ���
�V�� ��6Dܢ.DO�^�����BBr،��j=�$��`_&�D�Y ��3�	�J6��vcd���e�8Y�ED�^5խ�a��G�Q�Ӄhć�l��O���������ol+��(��zZ7�g���9lO)-��؍�i��L)��s�Q��.%���%�z����0�*�,��q�ڛ���aA����H�}S�b����G+�#'���Ԃ�m�o�,B(�	�:5a�l�0���5 j7}9�}Û�UV �k�I�#��q�t�|NQs
Z�}Jj��!B)c:��7�����Ӯq*����'��^�#���b�DYh?RG۽�'�~�P�l�֩ �����]��c���>"�1�~Pd�!c�(���Bw��s�:D����d�},�h��ԔE��]P��)_xC5[1�EBnʍ��䐊럱'���0Q�/c��RFH�##�? f�~�gn���}^"��f�����_�SiX�KT�\c��v�oəUN��-�� *�eJv|��*�(N�>{��H��c�]��8%f���^M�����������=�%t-�q�-�a�O��9)!+ �N�I�>�L�"�!'a/T����ڀ�8�I$��I�8����/���I-�y�!l(;�F�I�]O�l@s��}:��}>����Ìw6}6�~��f�km���=q�����f����&Ƒ�^�m����?{
5��d�jR����[���� P�/�������@7�dl{e�C����OT�9�X<�O�x1���`-ਅ��2�!C� ��\h������ �L1�^�@l`Q�䈪�OG���3)?�(��V#��	S]cR�C�|rOF�L���5�*B:�W��r\ã�Bnk*9��	XϻΚ�����)��si���ҭB�2����<����7�qT#����?$f�T̙3&��>M��t��&Ы6�d����OV<qh�1���X©_�P�a<	qtv?&n�,8i6���œ�Qf�����3��143��O_�� ���Iߓnh��#ޝ!�?�kA~��m�2��4U��\��1��T#��Q W���)�y�#̈́Q���N%[�x�UE�h�aCaT�~�d;�j�u����2���v>F KE�t�6_3r���aF�V5�hqc��#Ǽ,�L�-������,`X��Lx9({r-~�&E䀭� ��������K	ҳڂ��Ơ����qvG����I�G\ �8v[Lo�ˤ�j����#Z �5����^�B�=�A����	��ŝJ�W-�-=ALR�?���j�|�/~�����?�H�#��X6T�h��vRL�u��@�a��=�G`�Ύ�}�#��{W rzj�
��er*�G�+��wޔ��e�K\��!�
)�!��L�t�1��Ƥ^��H?{1�Jޔ&���{��:��ֶ(�O_7:��/|�t��v 'M���[O�F�&���|����?5C��J1��85���3?Q��9 (3�������4U���7?:�� �cUD�Q^֮�tY��>b<7@2Xu��?�QhT[�o{X*i����`�����p�?CJ��X���/�LTf:9*��C�|vH��Z,~,H��MQe(�!�$�;8�[S�����֯	�3?�����l1�d����Yiq@�-�COa�5f}OÍ�=���X�6�8Re�?��������`آ����~���E��!b>]n���-y\���Ԛ���C�[H.n<)æ���8����Y���������NO�t8D�9�ߑ�F��<ŋ��������U(��=�}Lڈ� pz$����c ��<ȑ��`��2i�'�8�l}��偝��h1�8D���[&���8�'��Ɏ�N��|�OwO���>}.��V���l}�]\H7v_�Av�KkS�s�bu4�Hؔ�m3<敠C2[������n�����v~C4.q u?�u��=�[�/�O��8훼�}:�e���yR��ň3��RZGY��鿡�b��B�HPx���Q���iR��R��8�j��^E�m�"pŜ�³��u���F3����vժ{u�G�to3�v(���s�D�:V�b���4XR�=q��Z/����U+��w�Q`���\�U��4<0=դ����9*��,��p���\���5�>)�D�U�\��"PZAJ|�A���B�`��"�	��[;�
(�߁?�S:G�|R]3�ϜU�W6�
&���.�_�x��1`
4�3���]�� �����f3�5p����������8s��4�}�R1=���Sw�c@L4W���CRN'�y怦n��{`|̗�_y�a�FE�(XG���05���4�����d���ϴ�
wl%[A��M��h*G-;P,.����y�>���� �J����Bm�Ar���e��/�N���������(���GD|.�#�j�y�\ai7�umV[��9�빬�/ )ᮠ���f���K�~2Ї��^XN>��.�>	�V�Z�?3YM��0YԨj�w�E�#�M�^�P�D��b��\�$�
���oL��K`�OP
=���狭��(�9_�y?�k�|e)�=�&\�K\$��E$�{I:�D�8�K�k8�K[
�`���p����uҔ#��!���%��)r֦l���>�`=5
S�A,�+q�Xhl%�#�9�l����@j$��8+[��	M�����[��U���ۻ:-ǺyXҺ0��޿A����*�J�a|��U>���xF�I=Y��_;l*�'ed��fm��L��s	V�N����r�3b�(f]0�Kچ]��������`0|x1YHv��v��@M��화k�$O���m���	�Mn���� Pdd&��v�~�jּ���lz���u�~�h�{a�~�/�Bo�͏ �%;���V�!��y���9?�l9��`3*\���'s�(�M�$W�K����PdU��isG3��`aS��3�@Fu%20A�WA@��xc2h0���������y�/R`-�}�#Dz6��x��^�k�[���Q���w$�Bױ�*ZH�(����䍧p;��}/��͟j8�3�vk�V��.h�E"ҧ�@��h��uCBU�2u� b�`�/��i q$�pi���}�CF�m�H�%����Fu���s�ul[b9�hϐ�gU�O��L��]yG�k:�:x�� In#?�_]�G}���e�=�şvR�)�7P3'��ݰ+�x�U0.�	�՗�/����1�5`�dE���گ�N�s���E����ֹ��� �=5����L��9|9Y��k�v��=��e���`�4n�7>��%�y�� g��v�Z�-�[�M����9T	�Bt���[�?�>��)�Y����RF�c0p��D1{�R���A���\\?C��fu[K��q�%�IW9�`�'�M�?��菁S���8k�,���#,Ճ�J�Q{Z�rL��3G�}��՜l�O%��c擶�x�yS��a����8v�"E��1EJ?�̡
���4��*^�X�%.�"�(�`\QIy�b8I ���r�~l�L+��ҨŪ iN�\Ru�5��xG��-�"(�
�@�qhB���
��R�1y?#����7T�|rĝ}��ޏ!��>&@��.l�q�B�gj���q��� u��O�z�`�	9u�dQ��f����$�_6K0����K{�G{��,�@

2IB�ۍs�_��U�]}l5"�g��=���C��$cT�Wzi����14@�e��z>4���\|�H�Z��~�C��qz��5ځR�šM�i��R?oe��jyr�fI���Ѿ����UF�~V�*��XQ�1�k$��@�Xs�*�S3��H�n���
��a����ަƌ��KG��o"�u�1�`b; b�ш���!(b���F�){椤s2R��p��7�X 9L��*}2dʒu �ټL�l���)䇶����nt�oq�H|�l�=����A-���`K��6I!%����Y�.;� -�zttsdl�]k��}�6I�=�1��cOQ���r�gf�D�N�ۦ�ҭ����QG�Ѐ��憈M�&v�ړj�@�D4T�Tj�����ʿ;�[����G#���6VI��N�p��X�����X�vn��6�/f�e��i��ͷ~�BE�_��?�s��ݪ��~hx*Z�䶾�=�O�
�+�B�w=ݪaJ�0B�`����
�xv��]~���-�'Z��˥r����ٲ�؆De�J.T) w��b��6m�g���a�>��G�gO�m��g_p�dYL�S���a%c��&4|��s>�Qd3�C��A��Vj;/�l�2��2�W���u��I�}��K�k��	wƖ����QdR�ŴPo����_r��o������%u����Z-v�P��v�s�7����כ�y���x�Z���]ާ���
�*�T/F�ί:�?�c_���p�*��Y3ܣ�a��0,]s!nlFH��.�*.���j���ٽx���6к�VxO�L��ٵԠYR!4�F��jN*,z�k��Q�6hYVAy׻�x!�D�0�(�!���w��ҖnӲ��i%Ή�0���ϧ�s��#��������(�v�fU�](���e����t�[���7��8�^x�����H�T8Fn�:C
�}_D�{OCBL��n�gW�t���$��@�߹EgG���ҍ����v��\d[��2�K�fv��/zg��2'D
\��r3���hf���Ḽ�pV��fO�����٢�~���{���H)����S�M�!K��20��-�Ħ���o�X�l"�I��*�^3;j<��x�6�,
�d���!O�)w�b��.ly���4,�c��l��Z�9Y��t�Hk!g�U,~16�E_�f���+��,�&��Dt�Pd��Mk6�;�?��QD�)�=�C@Cp���'��'��;y��'�0����u���MYՔ�,΢FZp7+G�=3m%��D��sˠ��V�C\w{����e�ekW���u��{ `Z��t9���	!����-���nj$z
*��p�d�+�K����}T��/����6
lr�/�,�NM }���s,���%����u�b���v��
^yl�e��x�

埾{��WBu���e�k�Pu����{[Е&b�9=\�ڈ�m|�=��h��:݌P��]�$�%Y�����3��:v�s�/�ar����cr|������^���x��H��R����[�Ի�z妄����E��h��D�2,'��-@�U���J�M�T7�4��+@���9D�T�ߢ���5�[v��D�MRA{�}���
3I^:��F�A�ؤ��R��>��qy�Нe�:e���}�5�э����xH~�>S���<k��〮��G���ټ�,&0��P3��#Ik(J��I�|K�)AC_��
5��@�A�/?��Q@!7{��sx��
Jq�gD��� �R���&�/�|�6 ��+u�ە0�S_�+&s�U�)�G��ŋ�,~���1i'9H!��B{�>�Ⱦ_5X�r��L)�W �+��8+Fs�̒p�1�s�@��:��|˷�
i+hA�� �!����s����m>�8��'t��%�r�x��L��H�W�E�K��7��'#R��m�������Xa`�w!�t~쀩L��c�m�0T��?Z��`�Y ��3���y{{`���.;���y@����3���F�Z/Z{���V����9q+\�xL*^P$��_x�Zc#���ڟf1�λ���f�f0;���Tԥ\��J�?
�K�oMne���蛭��>�9�e�}��7��̕���&b=��7m#��Y-b���DrJUFx�u	��]^>��R����fR <�X�����k(\k�{��\�p����^Zb��p��!I� UN��"'K�b�6_�m�6�?Q������+���oV!���\p�}nDj>�<���q�W؃���o�q�Y����S�W§��ȼ,�M̎�N�w����U���U�o~�1xgAfu�>*���8��%e�3P���
�:`d�ǃ%�	_�MF�N������q"���T*�� JE�P��}�l�D>A���������Cb��>-��!�N�3qx�]a��mɘ���ic�F�}��!�e7j�/��;{V�jy���+�m�Ѳ_L4�9���Z1��ؼl���oѺ+�߻#�'[6� ����e�����t�A�H�5m�K,�o�k��y��S�+�
M�A�.�r�ҍJ��Wĸ�8E<On�a��G�hj�&��x�O�|Ͼ�������*~r8���$���Ρ�-ͺ{�c�c����v��.��G ya����j9��B���Q k��퍡Fl���r��~�'J�)�n�o��UBI�������˿�R���C�z�s:cp�e5�F��D��pi"��Pmv�N�_�P�`w�;�=:�tO��[��"/!9�#j�8c0�D��J�H�K��6Eg.���)I��"B57��чw��JM��ȉ,-v2ͰBJ���$D��6p��b�z��-_X����jw�-S�j�P�h
���-$��"�G�<y'�5�m��*(���Z�5x�#���M��j������iۋ�_�QWs{�u�]~!��6Y|��2��ȁpM�^�K��h�)��Jl�&NN�@��f��%��1��~M��N��c��h4�?���/
=�)�H&S@P����X�����/+ʄ~2^_Dn����o9���6A���J�C��q��k�/�1i1R9Yb�y��޲�N�B� ��u:u�\���5��L�߼!��O<����m[�ޱ����R$	���02%�M�/�G��dc�`}Fl% [�%���2�D�S��Y�,::6����Ѯ�[��I� \����5;�|]�J�����i�q�-�]q5d .������sc^���5�(�x�?]�/u�ߘ3�t��{���-��o�=��M��g�ӷ���+hН����G��?����>���rÖn��~ �7��]��+�Zzuu��c' � �N���l=Ʒ*�]��m�W�(�������E%1�"_����5��?��P=t��c����VԽ^���t��2~�zw�c�����L�w;a;��'B0�t�x��]��d��1�����ajѾ	��	����^������1��Z������,�+j���}�@Va��&��ۊ) ��3���<��k秾�yk���ь%�4��>Yi���(2�U����R�@&���Z�K�������J�1"�T���p-�?k��=�k�($R����vXC����f��N,OXEu��X� '*b{!���֯.%��d�q���WPu@�T���|������f�.���'�q�JtH�N�\UT`?�2V:s9����^i��'��	>��6���I���u����״!��y@����1�S��T?���M�TM?=�DcT�8�z�|�x�0��Y"0N��'����Ж�C�y�nN�?�M�hHz�E��e�Ob�v�]K�F��r�z��($&J�Oؔ�ӃPah!Ie��͢U�_�T�W�O���-�0�#O
��7Fr���f��R�H�Fx+�m�H�<sޜx�s��Sr�nif�vj�Y	�'�rJk/A��p۶_�ן�kk�Er�ic�ޞ���6���0*��k��D@���Zݵ��P��\;G�6�X���FO����F���G����ŀ+jm�5�w��n���$Y�"F��%��>L�^p��������\`�g�c�{Ĵ�c~��^��{��~i>�Q��*!�t<�E]�W��ˑ]�-?�h��h��q��Z���\��dD`�6�¦��0���K֞z�u���>��n<���v߸P�멡����΂�ၶ G�Sn_'�.8�مy��!u(. Q2̜$�k�G�U-�C��רB�K����M���ܺ?��m�����`����U����:��XL8IE�a�U��"C�N��_��R/��S��x�U؋�֙���������mбBV�=���(ڐ�e��ƥ�u�T�1�)4؎3�\ �8./<��$ ���{�	5���� ���,Nd
�BLi"_y�Yg�� ���'�B2�������ψ�H �2�����y@V�C�ki�ψr��d<�����ǜT�oR`�{NT�ݤ�ۮZa�������3�Or�L�{�ʉzj�,{e�-PoP-�:�J@5uY>�y��4Fݾī�4�
�A��A���Q�ן11z���c�%p�,�n��Qf��H �1`�\G�kԗXs{K�2c�A�ϡF�� ~	E`CZ	��w&���$�+�3�!�PwSIլPi<�xN�T��i�AQ��������ѷ	�X؏����YaQe����-\�J�.zȉx"~��9�d&ϩ�2L}�]zb���]a������R��嵅n�b�x�kR��]xjx�x�i7^�un�r:*N7%�VK���4\2v��wJ�D�i����h���g+��nQ�y��-F�#�-�s!đP�2��3S?d���s��5��ʈ����h�k&�R��W��58s]wc>J����+���ق.g:m�$��p�}�l��;�͸�1FE� �J���8O����*�zZ<)�S�.��-�G�O��,/*09pm�|��q H�(>Z��~+���,D�Ԩ�`(K �*��ѧ#F5�	w�CTR�+-��t�&Б��< [h�mҝ5C^ś���D��f#�ǻK�g��U_��_�t!dc�ԩ�O� ������K�E���&N����x:1ń{�*5Qb�u��|V��l ]ʀ��-�}��h���E�u���
����^�4<�@���BZ^ 摎-:����x3���Ɩ�~t�c�[e�;�D�4{��z������D���3>N���2un�4�)OK�~/�x���9#yYU?i+Q�fM�ye9O�:[�6�_.@�`�w:iw�m�JXQ����D�
��^b�san4�HM���pHKi*��]V��bf�s�Bzga�R]i��E����Ӹ�3�[&𨜺�
�oC����y���˧�����%%]�O�{B���h�$e&��k�Jn�_�c���5�5��\���-�GH_hF�t���֞�<�����B�`�.=� ~����̾���=�DvS� �J�=�js8e�PWAڀ�͚�w,F2� ҧ�oInd�)�o�c,�U �M������%�'`��ޕ(pB'����3��a���%��U����Ԗbj@h��r(��Ʉ�P44��F�$ n��"�.";�0%2��'BND��J��>��j�<N(���"cty�u�E����_�ixPc��F��m���p�M�BH�2f�P�
�ͥ�Պq�H��pQ^�[��rmS��,�[0T�EP_���N�_���᩶�p�I�z�D2��(����>͹�\j�m�˦�
;+�)2l�w� �}�1��U$����1Ƞ�z��/�}�v��b8h����̹&\@
O��hC����F�d
?Q�\�`U���*}���N�=QWt�H�3�)�[<�����Z�K�儞�3�m��Y���N����6��c:�cړ�$(���'��(������Q�>A����P�����UQ
�($ ���&;#�Wm����
]b���Y�ʹ��r�}�
�I�f1��yS�+� �!��F��`�[-{{O��vkF/Q�3��Am�tu��j<��ê��T2$�Zs5G&{�8/N6{���~�-@�7b�W{�:꩸
X�g/a�N��@F.�EW�r�<��Ђ�>��2]>�Y�~���vg���;��xE,!���sA(����u$ť� y�c�FL���
����!<������}�	���*vr�#��etx�ޏ/E�}n�A����<�FR�	���.̳�ˇ ^P~�X��t:����(�_琢������sͫ�g\���'����X���#�R�BR0AR
ï6
�����t�}&��s���;��r�e�5?��n�V<K���ҰO1d�����T�Lt���H�X�r{���U�}&+�9L�-.����_������3^1���of�� cb�)�joG��$��ᮗ4^`�3
���b��vF0���� �R��8FNT����ζ�Tj��͹ꂢPYi'��|�e%ߺ"Y�8���n?<3& Ƥȥ\�7��c	�
�؊œ�Ug��{��J5ʦ�r�����R��a��Ss�e��m�{Ȗ,{I�C�7c\�3�d��oA�I�'0��q�UH~���"�Fg��VP�֍�p,���W��³N����RkW\7���(X����G9Ek5]6R���:;;��;��GǇn�����Ա��R�d�.C���`�6Nϳ���<��}�jp`B7��nT�������HWr���d���ά]9o�V�f�ճʎr�q��?��RR��sZԍzR/]y���Uf�ퟣ�@��L�B�3q5���L��L��P����m����A|��kD���s,='F��T]�L��G��Y��u�W1z1&4�骀���b�0�����ѵӷ�d�Q�y�t�&8���y$qU��֛Az���䘟��<<NF�u.#�o�m���&Lچ��h�OoM���b�����-ܜFr; �dS�b��"��Xer`�Y���N���Q�I���H�'��ՑR� ��;^�`ճ����B�>���&�&3��TG�z��kȍ<�f.o�p�C�ZwҔ�CT�NE�F�a�m����b���Z{w��:'�8Y�h*�wk>0&:p�3>67�y����������Д����	�o��G8"�9�C����J9<D�ދ�^LN���;���yHR����o��Fy�⮆~ZgX1�f���	�<�o5������؜3�����$H��?�oУ��'=�P_c�&J:]�ŃZ����]eۏ&�oH�7�"a�\���}��CRz��y@`�rv�)��N���^��Mخ�쵛[�R{(�|a�.��j����)�r]���6Z�l����#�hiL�����U����jɤB!E�z"ܤ�G��}�cu���2��Y�OL���h��|�k�Y�L��b�{_CF��wr�\���2�Q�7�`�f�k�'�v[�"TУ;[�.���@�M��r]$\x�J0`��pV)�^/��V�tZK�9�=���W����,��Ui#L*X�:�5�d
���RwT�L���󻭶i��l�Z�X�)#G��Ops�MOJb��s&ε*B�pޢ+ȝD����f�E��%��B��R���O?�b�)Y����m=IQ,׏Izx��3��\dMe�W��6�V����2�v�l�N#)���4fg0vu>)@�e��uIn$W�C��V�Gˍ�J���\�a%�Y<��6��\��,�ʜ��:(��:�ؿ�k�1%�b�vW�~H��eZ1|۝��V?�� �0�����f�9��GQ4Ԥm���t{0��>��6���5�m��캽�x܃zީˌ O�;|*���0�����Ω��-B��,����h0����&���RSػ)�i�\���oڪ��vC��e^��	%�G�R�6KCm� 2t��`�D�^�	�_��N��R���&�$g��F��;$�����.���(����Ѷ�k�;萟�2�8�kb��FHS��Z���!�D3�=��t�QRr�F���H����GFs���>ty���I��hjY�ȉ:|��yn��Y�ca�8�j�9��J���Q�T�-M�����(�XlXz�=�X=Ί!ڈ��RZ�R�f�1Po�����?V�|~��]�8����h㕹6��8����<�:��wc���.�̋φ>Dr��K��p"-S�������`8���������!"­&��P�Ӆ�vŉs�;�<���0!8}����K�QX:v��-������ƭJ]j?MJ#W�U�`�$dIY�}�e�⣾�m���9#��[����q�(�������x��{*������>n
5�V�e��KO-�Em�[�����"��'�)r���AI٪p��s�cx�N��_�fj��x�#{�x���trOX����ЂE��,��GK@�/���=W�3x�L5�T��o�`'k�L/C���l��to�#��ya�A��Ɏ�Nh_�?��y��#�{��ʃ�8=�"v�Z����|9�M[^��	U��F`Zg�仏��3L)�Ѣ���L�^�c f����,>Si�/aTN@<z���s���;Ȉ��ǭ�ά��0�O��T��:8d��/��q������5�QX�E��|m��`��G}v¨^Z�d��ƒE�t��R�������`�L�h��^w�ߤ++gc``'�./�l�E�IQ{c�d�	ސ������X����MŃ��P���.Ѽ�OgJf�⁧ǃ�u�!E�-8���zE��|�"�Z}ʪU��k,�l�#D�2XCpC��~�� \��Sp̡�-�it"�_ �6�Rn���Pޑ����_i���v*�!���6���+z�kB�?��r�AW�BZz.��3�l���șg����;E�||�Ą1ly�'��"��^�T�*���ɗ* �ڤd�����K��Z��ӈ���φ"�]�����d�}z���|���~ɾN��PP��N�Y� ��bs���6j�o�pznDY�C����Zaح��{�'���	�\&��܌ū�mG��[߽�;�~R�t�x鿨�}u~�,&ބ�P]�	���K����/�)������N�Gk:�RX�ig-���k.4{�%r>L�)54�zw�nj~��y�)����}�H���Vc�^H����[��_��_�mgwa"F����S�@�ٝ't��TB�5h�O%�C��WJ�ϵX8����K�S��ʯ�G D��xՉ���*��Ruc=�x��|f�{�!/L1���$�;�������:�:�^����ܒ�k�TM�3�?Ѐ��ul�C�'DuS�D�VYb"�,���c���oF���q�G:_��I㡠�3�U���U��ٖ-�W3Z�W�@��z�P��֖+��_��jf�8j*3r:�h�{&ϣu�[�&�����8nY(���4�E��D�gZ���M�-X��a�n}�xg���O��[�YL����. �������kD���gB�?�Im����O�A�%�+�dPL�wyAG�ɴ�L�p�� �;p��Ƴ�9 ��py��Y�&G���Y��R�%�o��r��3�f��[���-��OS;�B{;/s������7�W���P�75�b�'��V��uwf3D$`j��m�# �ko�*�C��?n��9�S��y�u5��rEJ@��z(~�0BV�q}E�~�>?f���`�iƌ��� i�PW$w���A����l/�ɧ�Cf��Fz�]_���pS%�3Cw�c�#��J���x�\&[�� Q�6`��,?S��x���<��a6�ȩ��&g�mG�%�խD���^�����2U�*6w"��7�_��hw�<7�)HF}�g� ��p>A��� �2������C�L�u����)ż�RG��ёv�9e�L��2�!O�����h=�?D������S���.ڠ=����vp��I�o9 �N�c��ǖ1��>Fu��p(u=�Xm���?�̈́
��0&�=�=�l�@�	�k�����^���|;��{nN�j������3��^��G�W���ڂ�U��ӵ#�B�g����ռa`��es��ʮ�����l�ez �&�C�Y�2�A��i�U�<1T	N�X�oI\Oͣ讂 ʿv>�9��"w�x�|�Q��EL������{]���Ww���Oh9SITRa�\M2/)�� 8K���֫��q,}��H_��pk�.�F��tj퍳�q��dOwزn�u`2�ٕD#�Lx��i�����hk�.�
�H#7ڑL��s�w�~$�ҁ�Ҝ�8^��F�O�ETǪ�~�c �!�`�n���z�-��G����{�W���ݒ� �bBk����z==�́"Z�ߞԣ#�Etx�i��o1Pu;�y�>	ڥ������wL\�5�c(j,1%���	��~�_���E��褠v3
y��LR[ڐ�&> [��*]'{6�Ƚe�P�L��1vH���yi��{ӄ�$��Cϛ�v���U.mr�O��� �%SR��� <�r��?ߒ l�`�v؁�丯��Nl�S�7���ڵ���6�`ʜ�AdJyֻ�l�T�]o>�l���k%��΃�ǣ|����լ�h��Ĺ��op׮��̡������ ��X-��	j����?�D�K�HU�AT�7z& a���_�!�һ���<:ۡ������+�xA �t���n���������;�@I�Y���s���~����J�@Lś�9���
JE87��{�{�&�rXD?�4#���G'�o�	���[���6>Uw�#�>%w�%��sK�Ƽ�<��yWr��E^>���}���ntk�}%fM���l���+��B�b�B{Q�~����79�R2!�kV�)~�)�O�̪�Fx��$v��|ȭG�ˢ$�ǻ�K���&�d�F#Hm-�]$�@N�Y+���I�&1bR.�l���bǝ-�f�#�f0��X��k�Ǌ#��h��~#R_<EW������f�j�S�����LT�FD�a=�a�"?�X	���Ĉ9|^�����N�+��~*?u�q4
S-�k�$e&�V�
T�a�G���B���ُ��&���w � G��*ˀ�p$!]�]�z�ƃ�2�ǯ��و��b���WS+ �0��i	���yW,Z�C���U|u�1��h� ��}SkaB�@����l��c�Q�	�D �9.��OQ��H�Ѻ��������J�����/��h� �;�0\�Or����AECT��a�D.TDN:
�ݣa��F��Bfx�8z�@�r�&-2���!O�Ӫ\**�,��y$,�5��W�y�U�3u�G�RG �u�SQ�R9S��I�������QTB.Hp�B��ȷ#zm�9����yA=�~��-��M=
bsq��@�����z�C���W=bm{��7������%�q����b;��B�a��V_v��r�<��V�sN���&�r������O���f�؃��M���F��!��Ԩ�ɳ�5䜵��i�-B���Ed�.+��gPD�)߇a�����1SM�R�{�C�S&�v��r0��������❻M��:_;����Z;F�<(4MY'$�EFp��K}r�`ip�q<���mm+,
u�3���t�&7�rq��1�Ab��u���X�/��q���FV~LP,GD�t���)��
��/y=	��1��T�ԫnH���oⳒ]D�>�*��7$���}Y!����ޚ0�u���Ԇ�����1���;��A���TY<�9���M�(d���N�$as�`���o��HG�Y�������-
a�sh��ٓF�dv#���:�S�Z@P&<=,S���%��M0(������H���Bvk���2nuѭ!��˗s;4c�zm G�UI��o��6c�pN5h����3�9�����']F/TbD�����c�l�ʟ����%I�;E��6d%D����"��jW�S����tM��4�X;��z�����v	s����<'�j�G��C��-�Z �4�߈Bah0�����9�K�f�]�_�V���U�p;�D�y�Jъ����^Mk��ӹ<뚑/I�7G[���c�nE���������^9����I?�""�����LE�M�i�+�ҹ��UxL�/@�{���.q��_)+�A�|�ko0�Y�{e���T��rI�j�/� WX�&��i}C��%� �F߬N_̶����_]��ۊ@���� vb�z�j%ރ  =EPd]{�v��X�vQ�T@��BV���wi}y2%^JL����U2����AV>�lX�Z���0H��<��S��oo�N�y�/�Y�)Sc���?!ըЩ��d;Q\�oO�D�̦�8�N�H��w�X�/SyX��il�" ȊA]��&��}؞ �Di|h7W��ֽu�uGPuD�+̟`�N��g���-z�i�U�����b6�HV��|����)l���ME֍�\u�gH��Z�{��3�uN��#�J��>��mǉY��}�s��:��&K��3[_<��Z@����6��qϥ:q��9TQJl�]�n�"�v�Wr���V!a'�M��L!7-xRKRoNІw ��6��t`��F�^�OԈa.e�kc�"D��Ci�0B�hR!�����Øo6�/��qN*R�<��uw_ujb�4�Q�����e�A���\�������
�f�7��X�~��}n��GlQ�q�M�&���od��` �����{�H1
��m���t'����Mj3j�ͥt�Y-�uI`���DDʨ�8l�ϰx1�h��O�\�T���;ؘ�X����E�3�-c��������*�t=�\(�d�8B��1�/��p*�(����¹x�%[����?��@I�l����G�^�{�*Ƴ,�W����[A���*�ɜ^Ѥ�g���9�o� =�G�`a:��qH�2r:NOT��C��U)θ�U�׵�	���)� s�K�6W����˼��c�(E^\jи��m�<Z��.b<du�a0�_'*�q���l9��A��C ����D��pѧ8��6�r�3LPz���*�BO������z�����Y�[�I�{�D���2��.b[�������k�����9����J��I%b��+�K_�$����-��G�༸�{�茝�ߚ������l�ʇ-mͻ�I	U2��S�g��YO���MUf��d�a�A�Z_2�$Í<%��,�G��2�����g�M"�vf�D.gi���T�&��ٞ��H\��$�/�R��e�$�����u^}�R����(���k�z���ʭzJ���cҳ�qi{n޻`��:�u-h%����#&H��{L�&&�������*��!^��Pԣ��s�x;�=<!�N�Y��߿:^��?L���k�@�%�Q)���Bz�T�n��٩�>A'�^}��#D�܍�[�\�8�V���	J@��l�C�RW�.�^C�tg�����W�1V�<��سQ:���ܲ��~Й?#^@f��6��0HxS�T?�K��W�J�Ǌ�}�A�NDY�H�K�?I�pV^5Z�h�C4��|S�h����H���L��ar'�S��u�����l�jmґUܴ��[Dj2,���y]&��0a���T�I����\���ϟ��J`���<�9%l��kc�x�����[��� \W"f�프`����5��������]_{�ܙ�<
ג�h׈?�4A��nC��u3{�����=�l���\� ��3���}�WY�P��:`7�PlКo�k�?�ؒ2nP���D��R�$6�#.�r��>@^ny��{�a_���!t��]�����y�C߯�:D��9��a6E���d~����.�D�b�;��=]�u;跺�%�k.�(�['�Ej�����%���>� gz}7z��:����Ҙ�DR�7�oD��DqHy�p`�b��~��Ƌ�|�LZ}h���>���3�v��� Ԭ�;��Z���̻;���v��&���c��~ ���IM���3s����/C^8�]x���j�Ǝ�8E�vԩ�8���t1�%����_ �I��A�C��!H*�	�D_A�	}��\Å��d��9����Z�%@���"�a<��~Te����jW�s7w��v�.Ǽ���#U���zRp	�:	έs�I(^�TbG���N����7hg ��b�F�@��^֏��CԐ.D��p���#`��)�6L>����� ���M�o���	�W
İe��,�:Y��RR��w���&�^����:j,��Qj~=7�d���cuۗ����h5˼tYV��	-#}�I��YO��Ͱ̗����$�@y�5��� ޔٿWJ_�6�U3��"b��ԯ���TxӋo�JJ��eԌԞg�����÷�:rva�E��Q��t��{�����G�D{O�\�Sr�2��`Bz�}�d�Q���k�H����~�2$-z^?�����k�>��u��=��2�����o����ZU%-�تa���|��tJj�����1NQG�ߏ��I���\g=�-T`�2w�jx�Ua���߀#�4���"�y���Y^��&.�S�(�|����ćb��윶�_~O��h�i��e��/�sug�Q�:���Gu3���џyF�>2��x��8�%�>��N�$�OP����*�L��9$�F'�iG+�U�i�z`*��߻�U�c��Hg��"���w���[�(�`�,z��!V�g��j�P��\S��Jz��~��/:4�$� 5��<��
	���Q<���PϰK{VM�^D�Lf~]J���𞵞��l�	�.V�n��6��g����7Y���
 <|E�Q<���)T���6s��*�jMJ�Ӻt|Y�I�C�2K��
��0�X��?km �ea��D�_�����'����s-��e�����!�m{�N����M��&FhL"�� ��9ƶJ�yg����}�92�UD[X��BD�je�o���15�a)���D99�B�8➓���ukD�TֺbT���`�+`GG𻐁I��uk��]ǜI�;i���
 �5D�����P!�VX�5s�<���C��-��q���B�R��5ߓ!]a#�@�o��̐�+��E�Q���1�q�(��v�s��$��������b�� IE��/�P���w�3�p�8>��̕h~�l���3*cZ�_����/��tSi���s�feA� �	�����b
nd��YS3e����_������k���i�__^A���Rv�9��� j��҃�бs��A6�0_Nx#����'�+���f����a����i	/kH�2�Il�FŰ�~��Jo?>���ITWO��턦��{�,7����79�&AA����^���J�FD���vY��Z����2z���@+�5���GԤbUJw��J�X�=O�pc����k��/HR��M;�M.	�������5�vit����3��3�(��)�g�D����cV+GS?[�CP^Q[�[r���$��6x�&��j����%��� J�[�+���U
^E<�/�V�H���2��õ������+�c�
��'f���uM�Yl�F��h��C��"��Q�V]|�_ ��~�3ZK%�<MD��M"N+�@'z����̌@U��i#������07M��Ρ����u��@Xv�o<���^�H�g���E�5 �`UC#M�����~__l����il=�b�-r]ý�{%M���+�3�+	��{��ڗ�`z����u�)S�D��:�@9>&Mi[�H�L/��g%]�U�s��YyhC�r4�<�%Loe$G1:˗��ը����2�[��E�b#C��/ޮ�����@͋� �H��!8	�Gx��7���FI`^C��m�W)̮t�FXʑr�b���0@���f�F(3#I�Pn�a���A�����&ZJg�;k�#zGA�bM/ ��l0r��`�sXF)�\��۽��3pّ/oD�G���A�H�x�p�����R�D���/�/+��
43��� ~����"���HC��[��ּFA�D�	�Mǐ����Mt����3��0�NT��2{�z	�dR�J'ԁ�@� 5� Q
[���g��}.�q{'���k x�7;r�X�7/è��2c�R�`�˕���1�J�f��[x�-�v6�ⳡz�kA̙�=%T���yq�ӫu��sz�]�v3�:�)�pWp/i�/8�I�"cU8�U��-5o������Ewc��K\Q<)��4�� �|l����
��x����X]]&s�)(���Es`B��������h!	�HB��"��~���d7�ݠl>	�t���R�P�`b�#N������Q���w��R.]I	��)I.��J�&���@C7:k��w�*۔ܤE�g�3�� �4A��X��)��asSo��M�^��i�>%l�'X!��h�n ��8����r��(���˜t\}	H�	s��n�?ޞ~�����ޔ��m���S}|�<�p��e�l��T7�)����g&D�dPr�3W���|I	����U�ܮ����~�9�Y��T�#������Zsb/�C�h�l
T��n:\/�N:0c��޴i4^�_���N5]R9�����SZ�������;{V�b�C[�.���o`ҫw�$GOn�<��oYC�K�"5b�9}��� ��%0�����-�̬�J�(X���^��dO��Ɯ�i_jPu�ԕx"1C��Q�#hMd�F�U(M	[�p�x̀r�j�-�=R�e�cc>���G��U$@(�ڵ�{5�.L8�p��v|�TLr����%����U�7�p&�`O����/Ĳ�|������X<
����-
���/�)M[:�43/:c1\r6�g[�d ��mb[Ϥ��[�|i�]�����x���Sm@����v�/R]-��5|��'���L���2�n�ۙ$!#��;�����&QK��qy�c��kj���菹�d�>�	�͆F�ZxD���~n��ې�O�T�<���g"�MJ��mQ���]���5�*���3�6.<j�De���hU����Z�dT�+��U�����ɚ|(]W���vM�/<y�[WC�OK�y�`�����m=��AK )�Ě�	첔�8��%�A����
���#k�JO�̼�s�n9�1�Z�\;E`��	g�h1,��'7��\����W�K�r�1�������p��<_~�Ȑ��>^5��gg�c��4�����	��k�r;���x������)K<�u2��"��}���"I�@�����+<�ﳯ�߾���
~�}���:�\���I��/��h��}�t����I������z*��LvF�ϣ��ƃ��8n� ��C�*��-�hM���x�}^)���:���
u%��@��8���V���\_J�:\�@�gqim����N��b��YF ��Xp���)��$�m������Č����#�_]��Tā茒�F���E�@0�
�ʥ�gJ���=���!������5Ŵ�g�4k��ۖ(��K����W��h��>hvi��Vյc8�frn���Xl���y���*DH��(�:�K)��b&d�T>\�4q�kYO8��$�ѩ1��'�N�-�OV�}y�����H��Rmֺ�W��������t�:�^GK-����d������k�/��t(�ܠI��൳V^�7j"�`_Yy(h@��Lp��%�ϺF��/��e���H�j�ˏ"3%C ��V|l*�y��3D��DY���C=y%�ڽ���v*<�cUs$*�M�c���<�Z���'k���|��iY*Y�&#�f��ZF�|���9�-�OT��᳢7H��@wOz��͑
|�˂�a��~pz���<���C��m&�Ê3ë�Y�t��/$?^17�#[Y���R��tNA��Y��7�;�$@�8x̫$�wY�0ӌ۞v\�cs�Lj�#��.��c4d��i�U��pM�r�8*�I�]����l��&�x��tBjt����P�N߹���Hp�)U��{��AG����V;I�􁏂2F�8E�W�� 6�����%�����d����\��q�;�.�}�,�������V�D�u̥'�Py�ҥwEب���>��f���u�&B�TN�b��uI�����ê�/J;w��	�/)P7���/���t!��M�{CH�>]�auG�mn��f��?ˏi0�2hfm��2�5#%K�U1�C�!Bv��w`LI�'�� hc'0�p��~o��HOy��w4�>3�9O���P�hhc����E��ײ�����\�*: �U�Ճ^�>Y���v�Qj]G�@��]��G�����w؎4��|����H��|�.�z�Gӣ
���]f�tl� ��3�v
?&:e�P�����ۤ�������o�O�46����b�^td]6Ͼ0���ǾT��w�U�Wk>@m�<��Rd
�^ϸe�m���|���mw�
�4�ґ�6�����O����8�(�K��e���c͒
+�zOM�R	]��%�����%�����=�Y��M`a��5�s<`{i�ԡ��~���N��A�碇e`�Ny�¾����2F2 k��&�J���J��<��l� ��#j�������;�u�<"aTb����>�����a��9C�X�>�E7����F�7'��������1�b��h%((ƨ��L{�r������u�D{1�B�+ ��6K;���a�6��K��\�)i�~�dὮF�L y\�g��6?�?W�`󴨗�%aq?�̠�QسS�ĠU�4-]��=�+J(!���:l����o
�c��1=/~�gV"�7X1ڦ����渔 �;�Nr
��6J�ݬ`H��:��>a&�(B��eY���@1�f[.���RQj8���Tu4�Sm��&ɥ |k�c����@�,�i����r��[j�R�MJJ�~V����kg��|r�q��ݭW0�ct��%މ@��|R�@H§��^}0Еe!����!�*wS�2v�_m��]��N�t�(=�薶�"����D	{�<T;�`�� �xT o���5��0SL�0*������g�P�Mwr�����������I�H�����t�$0<OW�W!�ҧ��mN�l	�c�����ua�Ep"�^7KEp3�_��"�m�f9V]�����W�|j(!��4q�[ݻ��ʝ}1\�	Bi�����~S�m��YņJÖ��gZ�?�	W�S@>su����'r%�>r�� ��ğ�A��_e�B�|�'g�>�Bj�O��u�\�C�r ٱ�o-�9��Ȝt�.�H����إ���LgNc�	!��� ]��4��jWQ��j�%���}�U�\Yϭ�ɗ���?�<E򨆅�k̂g����ƀڕs�06�$�ܦ�<�E�/��x'H���炣BcN;�kDW�Ѧ���!�6��j3���@��a��Kͤ�ts^D�dY:r�5�ք��e�d�)\
�X�	I� ���p5@�t���"J×x�S���������rk&��z^��FK?7��iJ5P�Ӡ����z�N�����wƱ���� .a��{�w3)-ؚeZ��z�Z���z�ɶ�a�`�Z�Yi�4)I������˧��s q�E��K�N�.����j����
$���7�(����0 <�����w��%�p�=�}��3L��]����K��Z�n-'���+�� zN��#�wks�Cl�lc?yz�<�g�b"�z�|����H��w1R;��C0?�ۚ`z��]���pKZ��x����~��Ɛ��s`IaL��r��e���;�|=@	�|1x�h����ӟ��]��=c5��i���7�V�x�q@�>�Q0r���
<�N"&^����5�:a�	����c�ӚbU	?����.�6���]zE�i)L#�F�h�2�VC��! X��YVX��n?r�o��@O���0�ui���.�}C:���(�ZD���h/�t< 5��.�0�`�o����W�% Λ�I[8�^U�Ys�@���|��#��4�쪳d؝e��M�{S/��E�����01X�z
����s��������k�t>��a�C+�������+����9Ҧ]�7ٚ�2�8R�l<�!��L���Uz72�U���KY�3�+�#Y��O��%��@C��C���~�gE�v/,^�>>���0��x^"W6-�0!�T[L��C�S:�y�E��5�]���Q�����.�@f�YVkx����y̰t���C�KH[z���;�8~�qvu_�;?��k@d�<�0m?!v����(@�O�5*{��Vh���c(��=�9[]��Wbii	Hnw�����Y����l�Y���%�k�켛݃����B�Dp�b/�8:_���M� r�g-���g���U�n~N�"�J�N���]��a2���h�DQ;�^����p��P/Hȧ@440���*�P�t;���÷Y"����?W[���׽���ƒ��Q��?PLKk���Z�Wn��1)dRZl�v�u��B����W�**�:���>�s^�'��
�@!5��,Jte�A�vY���7�q��5��>l��Bol��3�uS��'�p�p�;�.����q)P L�.�E���{"%�j��U�I׳�������������33���1��n�N1x�c��#g�3�Bz���$_�!M.��.�Hg�P�Gk�xB��eMwĮ��B�rؾ�� 2�9�S��!��W�O��9�<���<�߸P�\�a �֌��;>a��݉�7�7s�i_�io>�fX\8�F�X���=toI���M��i#t&jR�lG��b��e���|�9��FmZ4����N?��a_�AX#�v݉wFK��<�ۮ�'ㄮ������_��uE��*�o�W��n�OԤ4R
]y����B���/�fϔ઩�>	�c~�7?%99޴jEtm���sx@'@�<cy��h�A-�)��r����mȷ3[����۫���<I�|D��Ũ8s��H�h';݆��+"<����n�)�6ό�C�Bm���
Z�	|���+���w}f~��g�X����,{ɃlAQD��獒�#�M(m��+����Ӎ��v��,�q���V�&?皉ʧ;!���Ó����l]ڗoD�$-�}
���aT��n��-�)��vA2w%���G�8�,����S �����P2�s4Hg���4�d~�oB�r��ܯ�0�����I�l�XH|õ�E�?���\�p��!�n`�lDv;L�9�B�1hZxI�0��/1� �M�,�6PC~-SA:߷�K
'��Z&367$#T�ͻ]N-cN�Ke��PLՀo�j�:���
�9T���^5�壵{�B�X�u��{"?� ��r�C�����<�<b>�@�]���i��ХH�m}�E�/�-����/�R�}&���1����~F0�y����e@�ӈ��!��=�R"P��O���mm�a��E,�Bn{��R������u��1y�/�6��Uk�P����D����4f.s
�`r�+�e>)K�<�J�ϙ`�0�_ڍ_��YJi��?�����b�6Y����zs�8�d��\�ᦊ�mpu����>e^~���y�^��+�k�� ]�T��H�Q-��?���cX#��M-��X�x�5m��R��WН����/b��F7�&C��S|��~�����q�]5�c	s0=���c��3���̬F;��f ��9����~sn^���?�r��i��qv_V�A�]����*#����Ҋ��\xXy7�/�,��y��G%�9�l� �O�dӵ��na��n��I��<0Uxpop,��������#ۇ�so�P��B]�~�����3�2����a�o��/T��wO����E r*�ˣ;9��kZ�K%_�ۈ�~!�u��3k��}�JD9�89�����G�_�5��E��w��R��G������\h��j�
8۾�2�	??�$�ൄ�F���U�,݀�><Ŋ|!G��,;��d���M��+L$j}��Q���˲X���Ĥkw���i8���rt��)��j��?�^{N�k4��E
g�=J��Fqf�w���TT�d���.Z�t\��E1��7����ʦ,�F�������Yk�[@{K��@����a�-���8��%��Q��/~�s*qʹZ����9t:�i=e�a�*���AYU�c��Ĉ+|N.�S9)���g�����ϱ4��o{�9)bf�e7�7�J��8���+�0�_��\�0��:�B˶4Q���d*S͗��	�d��o�T�݊Eq������[��@V��/��N��iC�@E��m��~	�=�eZ��}jɧ?p�<A����D3"Q�z�nئ|�L��Z�
z�^¸���ߑc�F�u<�l3怘I��v�^�A3�����I�⇭���ޢه�G9�7z�\��
R�O�)��J�e*n�i�Rž����KZ���pЄ�9���I�ܕ�����=�� �f�܆��H��(���4���e�a�!��V"q�6�
3��r���mzO�����
�;>�����+c����q��,B�͔Y�gl�J��p����!�*�2����!�hb�qW�/�Z�(] � ��i �\� �o~�[��9=u��Zd���L�
�|����y!��<�t�w�ۤ�E�).�[$�2F����zi����|���}���'����#�qjÇغ[$L�R�� ~l5E:�����Wͧ.[�;�h#�	{�HZ�w���x�v�"d� [x��e-f8X}�U�4��жu�H��M-�#��D�ɚ� td�yÒ��6��cV��s��q^���}���-R��y7{i�x9A��R&R�>oL��_di�a�ߚ��������<H��! =%[�Yh:"������	��1���A�W�t��&�G�(}������U��&�_�(#(����?`@�d���p���sƣ������QƑ,�R�Q�eOz���9����|�b�"��2�r�� :�\�ǰ6y|��ۆ/~�U؋��rx�ܙ�3�=E�X�ۓ���Y�mM*��*R%��?�EUr?b=�rE�JR���п^7��z� ])a��P?����'��߁m����l�Em�Z񲉏�[in����wo楄��y�X$�b�3�Z���~��� ����C!ԣֻ�����X%Q�u�6w�_2Ay�2г��M6�� �'`Ҳ�2	DE�x����-(���.�B���_n|QE������x�w#�[�@3O3P��"�p��y/sr�O�n����*��p��U�J��q9Z�Uÿ�|���
��x�W�W� u.�A��7!y	��6c��K2ֻ���bs�;�r�ߨ��2��7Rl7}�K�lY)J��Ì��������1s�~�ܵ�Y�Y*�����&���{�@xn�������6d�_�q�����Yt�`[3�,@r �Z��pY; m�+�q���I,�N�&,?4)E�&�x.�v�")�����Ҕ�PX���u��h~aI\�>�]R�;�����O�z3��-tw/��!����.d�'븉�Ѻ�������[�E����W�	t=��m�R�#î�����,L)�5վi�Vh�v��D�}��4#�3����n��4�=�ҭ�&�e�9����('�(�5�G�j�������P�`]�&1��ﰘ3����\���J1H�(�"�`���˸�Ya����<�N�9�]o枌y�`��=��?����H��}	C�-Tٓv:�Ͷ��_��E�3�Tz�-�\x����Ga;=�����d|���$c�3
piII��5�n}7�r�3���f���K��a�1�Qpr����mQ�}y�X!����[��E&��m�+�g�B̋��a\�iAޤ�Y�zo�ONY�l�ֻ9y#� �(;H�<�`@�K�Z�&�a#�yh|�O��X��Ht�Gpߌ�5���ą�J��<j�ϗL�x{D��䃋������:P��fWǆ���x��&���"��3K�s�v~���K���U�K�GaN��h��[�3`�j�G���"���,}��LZ���p;��� ����QX@�5�la��k�k4��՝��eEp+���<�9��j��%߆9�0a��o��UW��H�|7�;��c�K:���47p�#��?��g��[)T�yH��yw��Z&��x����u5���v�'�Q�I�n(Xu����$p����ǡY���6��������2��&7�^�3��v7 -GO>�g��0�u�0!O��@�R��Qm���˥FŴ�����X��Iڿ��R�����g.0J�K�m�-���B$+�uA��������l�d~'���u)2��J����2�m�/۪�E2v{�NRp\���`C��F�j ���i��ܶ��8�~���d�^�ә�P͗L�y?��=p��ԃK�9�_�� �FO7���p��}�Vj� Ne8�1@�n��2i��vvO�뀻����Y�$R�Hr���Xe�}���P@�}�Y_N'��?̙�3q( �\W�'~Z������=�1�k]�!2�A�+8D�R]Q ��̟��%F6u
��Ni|xk�c�\��<.vBr��6��1ꮨ$�PţlWS���i=]��
�ty�Z�O�J�<R%˒� {9q1Q��2�j(T�ñ�
7�5�M/�H�4T�466~v�r��v�B�ۏS���x
��{���9�%�+��!L�X����-�i��cxX �nE2J�xd�V����6��������*`5���24�x��8��3�_��_�U�P�����%@�^�#ژ�|'8���a��nd�������\���M}��V�˖K�4ػXZ�]���P�6hr<�0�y3u.,m}q�G����5i�a�r� 8���[#4�P�NI=QK��8J���7v�O�He����&��J�$��}��w]R��-0c�?5.�|��~��Lc�9�9�	����R��ܤ:������˛oLP��yQ��+����q��5�%Ʋ�=������/�@�:�"s�����o�2,Ϛ�ר�\�90������?7#��9q>��}���p�E"��q��s��"�w�p����QK˭�����MR�|����d����ɾ
���}K!����TXM��/�VG��"������"t^�1��+=k�j[��P�Uʹ�(��������y�r���z�u��JX.���5�3
��X24G�4k���H8����/|�����ϝ�$��i��!����N�o����Ye�o�e����(n��rB��9�tO��M� c�>˒�NU�-�mt�C'A.����V�#�os^7?�@�т{bc�Í(B ��6`��'�<�vJ;�"���ky�0Q|z>�iG$�p�b	�GZM�:YR�eB�p�@���͂�4�96<&nGL��$�{}~1���]H�Ǒ�G.�$iS���I�x�g{y��#�5@|M���ND-��3(f]Gr�s�A����.ߒ��&+Ek	�\�]��K�;� r
*�L���\�^DyP�8�r�0�O �J�cM�F�3Q7�=�O2#�݀��F�z��@dZ��>�!� ���O�����h?Z�c>~`��}�v�����9��,.f��A3�m�aT�֨4�P�ۢ��T�D�x�~/�~A�.�3c3�W�qٍ ��N�����jNŠ!�UV^?�S���V�����\X�<U�|W����庍S"�,�����d����n�F�M^h���9����
U4�,�0)o��['uf�����ٱ����;��������L&v��X�)o��_A��+B,�f	Xy[��4S��H��Dꈧs��s���r[��2*� l��ه5�
S>@.��nCc*�)��u�ʦ�����<�?�Y�+Ṻ�E�S2�*�(A/f��w��7��R��W��xs�A��J�H5)�)��x"�bԁ���G�Y����D,K���?�	`��+e�+Q>r[��Pz���fP2y�Cw�0������,��V��+��֥v;�s��$L^`Lrך��,l9~�o�F
(g�:V�b�P�VQd�2�S�j�����KG�&�)�}.����O�Qqf��� �Ga�P�~��$iF���F5��qP+�9U��*M�?���D~f���ō��%sޢf�<�[-�q��#]���5��ұ��|��n�8�r]�l�}�����zH��,r-� �A�����>A������� �l��ʕ&�5��D(6n4\��X��o3ͭaV��C[�n�{�����M��� l�D�^%^�b��y�s'�H��`����?��순�:y��4}�|&Hp=8��󀲌���M��~& �H�Z��[IG�P��0-{Z����������xs@��k$�H)�����Q�r�f- �4�< S8���רc?H3���AD�v#�HpK2,�5�QLV��#���@Cت����NX�0���dg��'^_'��T�e�@�Ecj̰x:k������!���Ĕ��gFK����o��8/�ы0���/��U#�+�c�m�������+Em�B�O����a�/V�圸`�4��H>R�ʐӾH!�.v��+�]�C�ζ���'G���2K~��s��PxJ~I�d��Dc�C�Q�E�h��V"�o���%���z�����ˉ�{f7�r1J�5�%
���[�Z��*6���g�Ӥ�u���N�jQlc�^�����[�t^R�G��Z�O��!W���ncK��/�i\��--��C'�TL�*+ND�n�Պ�:"(Iq�Tp�O|\eD���xځ�R`@۰��E֧2E�r�qߡ16g�4lh�^�k��'����m� mVL��ns�+U8@�hM���3�(��pړW��`�̅�-/�2����&�\gO����u4,�u0�w����lGd`Ǳ��ر,F�f����˩lc�P�_.
��雪i 
� ɻ��#�Q����l�z�E/��U�����]*�����q��3��4S@��/�����Ln����'������[��P�z�_�v����!!9�YSˍ^�m3���;2��G3	�T��k�{
����sѲ��5�>]� Y�=v�&)��9��� �<%	�g'ݧ�^�X)8����Z�@���M�.F����&�u�/�y�E�N��?����t� �#L��S�\}(�AV�
�H�T�!y��}״$��n�����imc�屳&�(�76�D.�����À��#NQ�;�P!�R��q�-9-P�.��`q��Qs���![DM�:��Yj��J��=m\��H�M4B�r�&�v�ޘ���&�����u~P�gy$�!a�wQ�t�~Q�o�D��C`@��(�O��	�m,�; w�n�$7&j(���I�&��S�[���ќٚ���9�JZfT,����>��x��%��|2��	��E;���4tP�Э�ޔ`U�˵P����W�ࡈ#�����r�ױ3d=����1~<��/wy �}�,d�2kB�xD%��cL#+O��&��A����n��K:=τr2���#~iy*���Wp�#�p�)2=��+ ����O�o����0T_��U3����\R.�|/���He��]ڀ�9=4���i�����q�����qLK҃%�yc�����Gzp<4Yy��\q[��|���g*/�����:��<��5�Rp44�O��#C@� �.�o�"��(3�};�Պh��y.&���� w�ԃ��Y�����9X1�	��I��\��-
G����������=��՚��Z�\��l⋭=�ҐG.ځ�=|Q��\:����%7�,0��hwm;�EyYJ��~�9L�&G��/�0]�k�����V���k�X�T�e6X������0x)���i븚=ްF���:�u	>G*���&qmcڀ��Rq���P���jm�K�?q.f����:El��,Wy�7bV�P:�<y)|�U7ؔ��,�"jN��z�c�Qv����^���!���99��ڝ�����ޛ�D}��W.�`Ba�z�l����x���x2_C>¼k�<���:Қ���,��@Yf�ķN� ����� R����Y�����J'��������� &�����9��.�)n�,W Fl�O}��4N��å��G8��&n�w��iC�����K�qd�xT�S]�~�J�[��Ů�?�j��#x�Η�v�|+�tU/��iIkH9o���oB}ʊ�S�]�C��f=\~'��o�ao��z\s#��	R��L��\�7o?�@��y��U� �~W�x�<_�&"L��?3��ѐ�]��:����hʬم���i0Id��Z�]�(��� �4j!(z� ���	n��J�`��Ū���(?mH:�29�������W�/�a�@KaQ�e�]��^L�[�*:��赅T��i�-�B��Een�SG)��b$��CT�-��\�V���4,�M�q���d����O��p�H�����>n�v�~��b��baf�|�FO��H7+O�zr�j6�TvH+T�3��>�vK����E�?����^w�k��=�}��t�N@_���1u�k3g�<�lG(�������n��Η�K�M��6�����8Q��i'�lTj|;ٿ��D+W�¯i��	�����kء�Lсcj�	��/�6z�K������d�$��r3��NCI��Z���g7�+�B���Є���ٵ'v�UT�R���1�o쓿�Z��xp��a�Qz���>fo7�Q��&�����1�`��x8ˤ-�}�'on1,�Y{ &�mk� �Z��7ٿ���5y����X�f�t�ǭ����~6���e�^��?��HlOz+a/&_�~;D*�
��R&1���9�c�D�q�8�A{/UP�Ѯ؛	�|.���w��s;�ȹ�O8��v���/��$2�3$M̈�b߁Un�H�u?��:�d���|��K$$�o�c���������g��Q��m�HNzw=�uC^֡��C�{�i�϶��wܫ��mR�̰�^FLa�B�����T8r<�>a��lz�;~w6t�Z E��_�"6�xdM���t)r����8AG%���(�!wK,cMDt��q�/c���2�_C�t����b�|��ͽ�j�N�Ջa}ͨ�<���'�*�k�|��V�õK�Z�u�X��D�������[���ͤ�WY�ҳF���ؐ�H9̶��c���Gl��"�\��N��V?ᆹ*T�GYv��?:�=��X�����cb�Ec��a���.�- �r ����m���#�,�OG��V��M��p�e���6��؃�Gce?�1��Vi8Oa��FH�2y���#�܏5�"��_S��M���.��
m1}n�ja�G8&L�q�F�E������+�D�y5����c��I�\p�`'����t�e� �pzh�_+}`55�.��t��gTI��<j��n�MV�1����=������1�-b���򘕡ۅ�K���C�G[�<j��x颖0��<��_s�1Y:^O�@��NɁ���HU)'Eh�-%}f5�W~�8�v�p����Z�ύ�G���I���s�T��"�KO*����o���/��į�Wj�Q��c�嚇T�/(�R�	<7�4��&(�Jﲛb�rW�< q'&��b�H��`�m‒��}��j4f�<�i���6-`nɖX@>6|	���y�̎E1��Yr�F��������~�j���%�����D����TIaSZ���F
p�k�����f�O�v9��HG�`���9�NbBF�3y���u�u�ˢ���D̽ڃ �7�tث���l����W���)�0��"��IO(���HN��Ƹ&��vq�9Ծ�T�����TꩍL%%��I����~�,J�9	��U
c�����������P5�6��-}���m[�����˵U�C�K�Gy�ՠ��7��4��CKy�.��E��P�.�6j=��8�)4s/�H�7·���	����/m���"r>5�o8�B��J�rm��
�<�-���>~�ZD��ۚ��xQ�ِZ�H�<R�W�H�6�`겺�T<?M�S��B���l%������x�a&�v�j�\]x�+��}i�26ܥ��J����\�j1(�i�A=�Ќx�e�E���Z9�)��4L���q�s�t	�۷��Z�Y�����eԙ�u�*�����bH��b�ӑ�(�_5fk{�-�-�sN =F� �M�n�?�ڮ�q.E�M���]�h�t#�'����ph�dJ��,�ʄ�7�d�n�ű�Q|��8`�~g��`�S��<w�Z�ީ,�Nƞ��a��my��8Ҭx*���w���嫋`�ش�a��r'7��_(�1���즞^���v��@�w�L �+E�c���$%���i�7n�8!�y�s7z5N���fJ����;�L%�r�@�-�����ݴ��m�H�(uZ�SK�@�dp�:�����ul��o\k/W�p��=�v��A'@T����{����7o6|�$( 3յz��էv֛�pb���Ӭ��TVL��*4F��Cը��W����0�g�"��&�����E��O��X��Ǿ9'v	���TB���"����EA�G=�1Qc�cA�*Y�� ��t���Ah�m����~ �%��Gap�Όn������_����5=��; �S�	R�?;�V���o�j��Z��w�"�	;�x�b/�(zj�gV��eQ��.�x~��^\ L�_����n�Gɐ=�%�O�vi�;���Ʃ2���ߪ0"�/yh�w�@���=�y��l�ݏ9U�&@���St��kH�HqG�ˬ�`D�{�mI���#������*���	)2��y~%��{����h�A���%��rt��*]2��U;|y�KI.�����3a�;ٸ���p��g�1[�M��FtFp��-�X������B�� q�*�UTO�?Bq7��<jɣQԯ�E]tR��x� &=^w=/�U�h����r�Nь$PH`���v)�d����'3M6��{K�k.ջ�n5y��=h_�a[�!�·�C�s8W�Ȝ���"�o�A� a1M;��_�9��Rs���᧪`|jJ�mY��0f[�����B�WX�di�*�m�bN��wy��^,����RX��n�@8�?z�tq�#I*M��3`8�b�/�Y�a�V��W귺C��YOA�Mtҋ��V��te`����tB�yu��?#��P ����|�`@Nqf
)J�$F��E�O�����W�r��U~��s��������l�E��8�Ѩ��y�� ��nǤ�A-����	�b�`��=�O�׏}q�!���Q�-雠5��������TJ��A��E�H��x���-����,k��<f��b-�g��غtꛎX����t
��~�8��&�ΔӀ�9���L�v��*�r�J�Xh��}�D���[g����gwc4җS/_��`��"�GI95gҧ��y�٦<�#��叟S�b.^��[1�����x1K��j�j1�Sj�/�H�nK�hA�kx��%d�6
��-Z�YJJ<0@i$�#���mT�����#1*B[S-��Ie�#5��2=�Hɗ�q�Bc�����*�`�j ���BSv�o"<T�;(vZ|)3���p�z� �ظc�ز!]+�Ε������"o97>(hW@�rH$��#��9���i�ַ�) M,���NK����zWh>�f�,�%�����3}"O�Y?l��ܨ/���5ͤ�F��,�&����˩F6�,N7��L��Y+g���ے�s�L�Uɓ�7zv�@['��i9Q��c�{��Y�0�Ϣ�X/�%)ԕ�-x����!�sa�"3B]��y˪�S�"��O�:6xo���s�d$�..��\[���k[
�ܺќ����HKUQȈ���l�$��:<i�<	����ђ�$D��;ƒ��,�\8=�*"֔#8��V�6�&;S��QN�s��?{�iطfǀq�G��F~:�~�b������O�������Ʈ���!\&tCN���7O���I��H�m���D5PΆ*��I��S��n�!}gk��t����e>���)�q4|&�'�!u���5�֚�߂�uP������{`��<��x "du`�ciAN�ITW ��]`��Yc���aԂ.Y飝�H+Fa�iۊ���3s�-�#�	���@-���� �kar�L9$�h��N�ݽp���P���*��B�]0���t;�P�9(�w��,�k�%�d�" />Y����RLls#�6���L��_Oq]�����I%�//����+p3�\��s4�y
2m)3�kڄ��
#���cΩ|�.|��b�	�*�z(�ߛ,�S/!��"N��AWN������Y8dG�!�����ŗvY���=]���Ig�TgY#�IM�Mx�L~��ސB�Q�{X;:c�E��+|�B`�?I�#�5�ݢ�c�i##�l"���M�����'_�Xz/kfim���Q�bЇb� 2,0�~T0�X\�\Eo����_L$%�ۓ#��b�LtF	������s�����Q�9���+O��x3x;H�;QWЏoU����]�BO*����Ȝ ���Z��Ⱥ�g�(1�k䬖�^XF ^��|�ԓ,��p�iø�bk��n�*����ߥ��LBP���]e��mz�fڟ}�d�-8M��h�W�C�H\�R�7�A<)�D�s�V��<ǽ�co|a�5ruBb������<h�����)kFz�6�X�6u��<��,t"D��2Ct����՚�DPĤ����4��%�~ܼ�\�,=:�+Nh�&s�NR᫵g�'Pp;��74�ۧ�?�]��O��3*x�"G��E�Z.�m���m��B��;|�(��F�yeN�R�b�a@��[AmO���U��l�Vh�ēt � }�9�v+I��@,Vrb��P����o1��|�����,I�l7�;Ma�3���U]�N�Ȭ�V[��;�&l(�$]1O��������ʹv:����Nq5���VZE�b�Ȱ}T�E�a�	BH̀sz�D�|�M"�T�(�&��(��Z�*��H�*Q&�����>�� ;�Y�&`;y�Ǌ�m8�w�i�iT3���f�z�pI�'�u�:E�m��o�Ni�p{�Q��~��M�ʎ�_�ۯY)\C�1Ǹ�I.T��Ɛ5� �0K��(��
W��G>���Z��oi�t��	��'4udo��p(��f��]naz�z�T�!��q��ey���z;e��{ݭZ�q�r��G��m�]�g++�'MQ�A���=��V�8V��Иɥ�(b}!9UPa�Ξ��z*k�����>>{���r�~�\���nhi�� ���iDo�O9��=w�)�R�7s�ѾR�A*C�ʲ}gٵ�����4��zl�J��a&;��Zs��n���oZ���/���K
Fm~��LA�D~x���?�%$�:ŋ+f�A�x�+�%�`�:�1��^�5�+��l����4�|)��;�\��yp��E���[�p0LO	�71``����8'N�O�8;*	X�l#-]�.6g��L�I4�߹�;���d���mŏ����;����� �#1����.��*���^&���Y#z/�HƳ0�a����wU}���F�we0_���@9�����O�J�I���2V\�b�W(��{=�C��[*֣���DC���.Т�y�{�Yװ|�	"�G/��긡��q�\����fʜ�G[������;�:QJx�_�cs�r
���G�����u��5�'-�0C"��-c�Cq����
�SL����U��xR�F
p�l�UO���?�)����L@*,���k߰)9�x]_bR�"<G-��S�n����X�a��&�V��g�g��Lr�ڤ����R|.��XO)��p������ ��[{�bO��A����.Ԯ�G�6�P̺`w*��;|`��?q��7�A�OF���B����v��Zjf����'/ճk��M�5��D�E.�	�'g0L�Cf-����p�:\���ub^a�2���fU��s�q
�Ⱆ�t��q��l�',�PJFRhQ������P��2�����j�����e�!�G�(�+��t1�;jkY��m�wH��،�.�&�3����[��PYe���G��� ��p�Q���N��u:�쬖����.'gec`n���"&�#��?׈0�=��fX�����P35��C�X���\���ct<[��^�P�8	�';1X��T��}x��+�NYۋ��,�ߴ�4�
X�ʭ���=�l�X����qQ?Uqq��JGԯ>������/#�'$tCEn��t�#E�͡�ں����UT:���{����zbT�w+�k�W�f_n�,cK�`Вoro ����w����	S�͝-���Xg%���>Ѻ\�$bgL���ل�g�߱����-F�7/��NWU�JA 2�F.�$	]n\ ���ߕ�P @�}�ɋ��e�2�vP��+Ɗo�RiΫ���%E�n�ۈjG�����MQ_)�X�%�"�܋������R�9��]���4.�-�&ilI�I��hi(Č�V��"��'�>��-��1?�xZ�A~��d�s����������{�"l�`RW�N��Y�j%hcI���Dr�ۦ?�r��Ƨ���+]�*�%c��[h����W�B�?������~��ԁ�+�q�Ӎ�|�е&P��(��f%�\S�Xs�iH:��]Nh1���'�o|��o�52�6g�}��1=�]���eӴ��5b�jx؄����.)4]�-r�S"υ���$�E�f���g ���l��*�W2*N��;�.-�P��M�nx:�`�0���R��Ѥ�H$�=��@���`@�{a�6Kӧ���%f�����+�,`�A��᷻U��ZD���n�p=�M�)��ϟ����16��o'g���.� g�=8���]�r��(ZĚǰ��Ȋ�#��Èt��r ���;�돉׹�$ٷ.�bS�<�u2�5O��9W�ؖ���I� �U	��歨�박���?z�_��7TB�)�P�O�f�w��cJv�F>�/��]�4&�M�Q�r�%�8ہ�PU$��ap�1O@ǾS/�
��z�������O2b��[YxFe� 6N{)�Qb����	���v.��d��x��[d�T��I �">�NTFyG���lfwfR�qK�w�z�
Ӳ�0J�+�c&����/�3$�:_�<�J�"�w�֒��%�[��"_`EC��0T�c��:��Ϛ�𳌳����Sy�&�?�YeJF�Ϊnu�kʕCSjT�[J3�)Ǔ矻u;��{^�`� zb��'XÂ�i!�����r�Yԩ`f�Z�C�f#yv���P�
�~;� _EΞU7D=���d���m5���2\8W.P��X9i��߮`��-ڥ��깾,��ǝ�����xi-=��`�8q�׿��Q���K�t8C�c��F�^�B9ؔg:u1��d<��B��O�͹j�^�E�a!����3����/$��t�_\�w����2ʼcg�yP8X��nl[mQ��j,�ec�8���9"�[�!���57Zx}�NѬT����975�3hXP��2��Cs��NA���&t,�e���}I��
]�H��j��5��?��^7(�Z�HC<������o����D�0,⋃�ԛ=#���g޹*�VB��!D�!7�}p���]{�]4�PU՘�&�j�5�aiyy6j�Z��e� �>��gu��V��(p�D���D�^	E�I�y���L��Oqё�^�A«<J����B��W##���N/���l7W�k!�\X���edw��DHr���U��6��`�K�d�XZe%�#�|�M��ҖX��1I_�J���g��B�7h��?}�w�q����J�!M> ��;z�[~�#6�s(�-��K��������m0i������OvQ�K���_MhgP TL�2���M��A��8���&�Z:�SIkK�J?	+�>��H�k�'-���8l�y��X�2*�ŋL�>�v�mTF�c�Gh1p��\�:3��阢�-��GY:;m�Ď��\�5���l���δbS'�4T���?�K�W�S�L���zU�e�𷽕 ���N*$��t�CxiK�qY5|4�|:��L�SgDv����B�J~��,�.���ՕV­i2��bs����F��L�:�����"K�Q	��q�ƅפ��Y���5����jJ��ǦKp��~+f�`�V�&���.T!j���;�W�2p���&F���<e4 ��	C|�?�kO�a	]ˌ�ǨQm�m�di�X�?i�\�)�{?��M��Su�!>�<"��zW�^�'�!�k2�~0x�S<k�C�K0�pW�����3����7�6ͤc�gFܨ��9a��~O4T���wCk樨�m� ��2웆�q�,�Q\�����|Іrs@!n�:��%� ?���BO`Jz)���*x�������Q�<���Zp��B���=	��$���B�Ͼ���v��u����\9V��E1�	�n�oVo��{�79T�woH7�;F}!��TA�m@-�
\��GOp�|��M�Xx����|��#ձ�D�����G��ZM4$�`��{�b�p�+�u�A��(��&B'�����
�@&�<�W�:�ը� �� �4r��O�g�"�_-I~��FnnyF�`u|E\O`�	K�&�c�pU�<]�K%��Ol)k:(�I���x��i�
�.h��:&B\�ߡ�b���[�|2��'}t`�'c��nMtF��?��gKPRk�A[���y�'��A��m��E�ܶ����z�|�������ˉf��e(�����6Vۋ��|(�������&�ӎ6d�R��cX�=e��i�t��\x9D���&s�G<��xcc������<K�T2 >�Xpp��A�͞��^Y`L%��ĺ���XV]����lX�Q;��A���a��xG\G�����T��q�h	H��J��?�ጵ����L}�	(U[�>�TkG�gM��L	+���n'��mf��½��X�ѱ�&��t��fw�����?D���'t�� �G����}�jY�>b�på�u|=��v(5�ь�x��÷�g�=��C�7Y���i8S��ikw�Cp�L��C��ν,���-���S�Mx����ز��es}�}WL�[� !-v��H�pjc��)U��0F�G��(�>��fNIM�岱F�c
��=�����&�Ou�^�X4~�6�s�}��.|��V'����]r�.a�jA�Վ�����;Ɇ�����\+WƑt��+���BU{�U�gS�S9�|w�,!�v�s�ml~�7sdlL���%&H��cЪ�Gqv�s:�(�W�C�D���+J:��#"��]�����N��!�ģ�\�X0�,��_�7<�$uC3s���IS��[��z�cZ���<X�U.Pei��ide�T�O\Q��G	K�f�I�ٸ����9�w����tա���Z����7�WI��+�4�� �����r2���[5޶�p3W��Ш�1{���'?��z#�8E��T�L����k g;��sż]T��5o�x'g�j����k#Qc�R`����*�(�)���F�7d��������t��	���C#�ǯ��HpK�m[!A��p���Jnw�_"�; |;��V���BE�����2dQ�J5��P�G��]�u�î��M�
/'�hx⼩	ץ��U�X�P�jF��f+ƥ�M~�H�薺�"�F8�X$#���E}YO�V/?n�`Y�I�Ja�����>�Y�o�߀SW�E�[-����3���& {�w�>��ְ�{Ac����U�˶������+�.+o��|=��߼�?P�N����i��OK�-��V!��Q�����:�`�/i7�6�/Q�ZõUz!��+��Ĕ F.Sm�3Ko�1�������05L����ISV��%T�Ƹ�te���U�4A�|i�U�b�.�,�J� a\��\S�[��~�~y�Uީf�0��	7�����#� �!q�tؙ��0��ړ���A��y� ���3V�s�(��`D�3�'�pu�BB�י@��E�E���:Ux��������%�����]��5(�Z��JR)�ݸո�d2[�/ZE,��S�$�H��!�<^����F�����>8-��6��t���p���������
~G眔�%?��){�\�����}�P��5��i sl��)W}�w�&WyS�8��WJ�����|�d1wH
�����E�'�.R��:�m��7����hqry��DVD�AfD�8�Om@�O@�(�G�h!L�8s�ہ~�������J������jk�t���=��t{T��U���8��jW�BUD�{0j�r2N6��F���e]q�f��-<�t��J�Q�/���gV���i�ҵ�<&0	Gv���h�M�X��\����wޗ��=�p��s3��z���)gK�V{6Ŭ0-\-���ϴv%w��e"Jj�W�BXװ,ΐg���d�u�w;C�=g�X8�LC@���D}:�8�ktb��5�+�I*OQA^�\���S�F1���%�D�+fkgJB��z�:�����j�DA@%�
���A���ʜ�}Bmz����^wǆ�b�E�'�U�WK�WiE�0l�TO�!V�8�~sD�~�ŀ�Q���J�l ���;>!��2f*����H�Ɓ�������7~�c���'S{RiX��!��/����v��M�PC�-g�i���#��cE��L�nnD>DM���!�c�z!`�uI��J���������
/d�����W+=��>^ooJ����&��rKR(�+��q�ab�mw����-�P�~0l��c� �.���c��Z,�����t�p��_p���ʒ�4͕4s��Xɺ�������>��󵶎8~��\`�U#��nTcH�\�yJ���-ߓ9��pՕ��ŧ0�
}��mҦ�,��!A��z�"a���g�c���� �n�LҪ(���Țw���>xT|���E�{(x��Fr�)WQ�'Αc<�5-*�]���H��9��u�D����j����a<N�MgZB��:X�`�_p5�7(^��m�/V�T��{@Z�޷��_;��;P�o����_)}��������HwnMk�g�a9L��
�6��6��/�Ҳ>tW���i�%��2��&4�o����sى^"�)�xN�6g2ǣWw��p���SZ�B�ǇfU��H�P���ɽ�ܵ"sʻ�5ǡ��}�N�VSN}�D
5k9���FF���}֑��B����έ�����L=�]�w(��}1*,�.��٧��zy�oh���n�)_�h��Cq��{[v	�}�u�)ns,*�8a�3&�K�pjN�nVo�����~m��9���w��_s�=2y������J�>f�����(����+q#�|��u�G?�5i�7���ӇT��m�-�T�'=�]��$I��ځNd�&B�2�"b���L8e7�nH��0
[$?m?4���du�(X�a@rY�� �����{� ���x����<��y��F��A�gĔ�=���z�;���ַ<���<�;�^���E DX�b.k燒�ǄRZ�fCI��߭��ˠ�!\ji���<בGz��g�LI$��(�sc΁�!Q��&Z�Th,|��/۹.EY�+)�PAӿ�P��GZ��L;�[ô�?�0lN��B����*rj��,E�	���e%}*iy�4��"���E㚅��'���`h�0m�ZAr�^7�n��6�i���O����L%��l2�j�[��p�k�^�?<21,�A\�TU�nІ�kG����>�L���_/5��C���������]��OǺ����U@ڴ��yW�O� �.��JL)�<��c]���T���������t6�e��$7xG��_?�=�]�\�B/(���<ب�����	7�5l�B��LE�/�t'N�1��\ �+�8��������ЗEj�4ʸ������
���l���%čCȾ��58���#B��K�od8�p� �j%������㟪�K��<��yz}��r�o�m9}[����ǿ��:�v�eɋ�Pf�]jL-���Ű�$���6�X��O���$2�tw���� �=C��xt�x�vѳ\�Ӎ!�i�H�R��}�@�/n��»���������:�Q����z�99V��V�tdͫ�pn:��C���I�>�f�H,C��O���_��i*1DG���&�$u�6ٺ�-��w�-���GK�1��E��_�b=��Ɔu8�o��Nr�̃ԭ�y����
_�ĔN���JJia����6�t`�_/����F!���J��ҁj�p ���]���N�m���6G�s��������X�k������͹���h��=z`���@��?f��,H�_�lPM��Y�5_��5O���|�3~�g��w	\���g�5��A��˫`!�w����`>J�/�uJ1t�v"?�]��D����Bd�8.����ڰ�L(��f�3I�&���AR���ƣ����b	�u��p��c����o'��&_��3��O�C)CC��D����tC�	U:�G�J�Ci� �"��a����$�Y��W��Q}P[m����� ��cN{��(�G��P��R��������f|�����6��Q3Z(f�_�\�_sY�΀e��=�~���O�Tf7�Q�H�%ʍ(jj������õt]dv�`�K���y����B�8T���-�$���AYݟ����W���ԏң>{[��;��S8~<
��k��|`�v�Qֵ����"j�-���7�Af�b�i6m#�1�5nＶ�	����^�Ҽ~��q}���u+P�[6��&w��.��YU:B���Lő΄ݿA�����8-��Oy!H����tg =kL���W'��q%U��[tk�Y��@z��H�2	,X������p"P�S���&��`��Urq�k2J��ȱ��RGVh����MN���;�4��+�WT��r�#?e{�˼`�^^Dc�[�g��5BZU��e�I����'�\?��PV��J�K�ހ~���k�$��S�Wg���/0����O��]Y�L�y�"(9��L��@�NɅ��!�)Ȱo�e4#Rg7U]���%�[<"@+��k ����4c��a��r��|�.�dKS���n�@���_[�M;��u5Twq��U�hӃjhq���|^ܲ�	4 G��o�A/��J@)�fԦ�-����/h�Y���e��̎Z�qk�m�n)kd�eb�R?��Q9���=a�� �7l%2�x>������pn lVsj��B[��]b�^��8�����n�y�ugMб	Ê�۔�tL����(��x�ۊ30ag`ٞR+\��9 _1Sn�8#��V�s_Ajӏ�9*L���K�����S{g��w�G�R�IoP��iUP���B�ٓ�\ +$����~����Y�d��k��cd&�{ iZ�jU�j;��}0�y���\��������ߞi����}���J��4+��+��F*2�3/!3|8#p�������ꦎ`Aq�ek.�_�F_zq0�COc��7W,q�R�p]edJNÌ����#�o'��QI�]���2xj`�sV/0Z� H�,��� pV�eC��+;�ُ���%���%��Q�>��8rPE^[��.��6�@�ڤ�X�)w��>sP���أK�mHY�JA�YP�f)@����јs+O��P�?�Ce�%{�]W�a~�3 ��P��/=$o��
���֔��F.���N��i]i�0��<��MÇ:5�ݥ���)q1F3��� �WW޽>WM�O���v2[�dȦ�.�t�@��#�S��@�T����=�Q
[˝1��v��أ���7S�V�!O��`E�eOL�;��L�*Bp\�?`�zT���|��0���RӬ�G'�$�d%b(V�$�b�c�~�y�cFh��ѓ�c��N T�E{Ì+q_��ca?#2ȉ�ধ{Zo)��f��I������	=�߆���|�ύ�Qi�;��'��]8�����|�ǵ����9>|��������J��o�w�h��H��<�z!�Y�$ �f�˲�=(b���+lϖFadO���R
Ň~r��{:��D�ǃX��f��`��oYb��]�������^��H>���W�{�r��WԦd��~�5�FK�����H���'%�E�B�㨝:��_��I!��q�0�32��A����^)Bv���g�O�0��Z��z��(���Aj0q�&�1���|�޼��Kf�.&����d�y��`B6�n��8�)i|�p��"�f�>lY����ȣ�����BY5�s��ѽ�<D�R�|�ʪ�*��JE9εz�ڸ¢p�=�Q��'P���~B�a[�f�̢�AM׎��bvf���Ͱ#�x� U�����J�Ȧ):����ݨ�G��l�x�cu���V�i�+׼<�J����:�r����舉y�s�Z<F+�Ef�	�y.}f����du������ܬ�-r1G7϶ex�0:��Y� MHԆMX*KY�C�G��V<n�t�zR�ᖇ������Onݯ\L�3b�E�0�ߒ\�?b�"R�l�Us�% ��g�����J�\���܌�`iR�AMП�-�.��������|�~�c:-�?n��Ԉ�yYw:�{���.E�����Ϯߐ1�Do.���xb#��X��6>��&��9's�O�Q�B �Pʮ!�t��T�����@k������8�a���o>8�6E�P�<���O�<��f�⽣��a�(-\WM�괖��cH�<�R�kQ�[����W����}TosQ��\5�
 ����#O�*@i:4J��t6��rjQ�`��5"���5���M�Z��'9'�2��9R<ȭʧ�` è�cpJg�a۴ ��aI��r��u����S�:73�rX�+f��Tq4�)v">�9+�"$�.�_�*1A4���S:6�q˒3A�Z\s�o]��2���
T��Zल+d��z�g�r:||$��.ܶ��IEJ{�H��1h�#�iL~65 ���˂�5�}8P�`C��R�ޮ��>y��D�3r�M"F�C8���43��!��s�~9!��r��k%��b2;*��`�3w$�����I³.nڢ-�֖d��G�H0��.4�?�J��+?���t^��ֹ���ㅗ���,j��z�&k�g�����욹뜋ݏ�e�v�����D��5�^�ؕ�7@���wH�ӵ5.\��=c���IWs�ؖz����x���V�;���~�
G_�~�:p��θ�z/W�:2�&��U���������R�����|~��z�'�C��z
D�ؚ��8\]��"촖��d��t�)�mn��.#q�ѩd�gڗH�O�K��	��f���92��|"�6+�3�9b��Q����_=-���[�F�?,�0���6��<2��T8Y�A�������^K���ܳ���T��"�3������%�苝xM %Q*_�杄�wD���D��k^ | .�Ɖ�o�l�"�9+�Ork��]���'�b($t/���<���0�+.��W��_�6��!��$T�+3��E����|+�t��=�L\�U/Wְ��]S�3$���{��zk��p8mB��b��#��~�v����(��_�s�cCب<Y���8͸%�Z_	�(�P����b��;4ˠ���K��!�W=��W6���h97s������Y%7�O����g���3��A��]b��Tn��Z<��.�4�s�"5�;Č?��yB��������*X,��G�5�{��2>�h�ʼ-*���7xP��؝Z����tqt͢�̡}RJ$Kb�����5g�{I��d� L���;����McU:jY��P�MF�;�Njl���,�`�D�opŌ��)��Y��A�'��UPL��c���- #�T�� ��#	 ɱjl>Y LJ��kޚh8����>�ܚ��K��k�9P���:��&d)�\Dv{G��$[���u�㫏����^�Ԧ�%�"UJy�T"�e�JPjFE^*��7wm5�8#f���i�.��i�F�
�a��dǒ�*� ����ȍD��<��6�?t��ӥ���d�M��9S��H.?�cv�!�Ŭ@����Ƅ3�`�'tl�m��;m[�r!fY���^$ԏ�[6�<������~�Y���z�B|�����J�����4eD��� �e��7�F\ʧ����Xxꁊ��\Y�`�]8���v ���؂Óa��^~k�an��� ��#�X؁��B��#�|T��-�\��v�CG���eع�Ê)E4��eeE;�(x;]o6��<��i�������z�u��'J�q��On�?E4� #�����Nq��$��#�Y�C(��]��j�O��pZ���*��l��ަ/ʔ��L��P�c�y����G��^_��<h�\�0�};�p2��p盋� v�t����Õ\�x|���<��u��H�/bd�O���[H\l����7�x�\m��t�%g�H��ꢩ:�,q��G�� �
�:^��Y5RF�0����>�۹�)鰍/�.@8#�s���+�M�<P��L�k���
��6�%�i[�܂��x����T�f�/�d�ďS�2DT���0����S�m�ո6P+�(�o�v�-�j]����p��RW��q�X�ń9U�f��9�����%�z*5��e.��`.76� �z��ss�JKs^�Y����ǢƠ�<�������=��K@m�PP��Խ��v�3S$�;���9Bi>B�ֻ�J���|7�=�)c�5�"����U�U�'�"��o����L��^�D�ؕb�4�p�����m�����uB8L쎀���z�X {=th�\��s�Q�w�&k�u� ��g�2��.� hC����Hp����\��z��Z��.�:^_Zߓ�"i�W	p)eZZ��m(D�S/�:���Q�t�� ��4��K�<:;���5���<qn����(e�vt~R4jFU��NHp@XÃYN�3�Vԕ�p��e���������Ӎa����MGS�0_q ެ���/nQ.�h��,�1�J�QH����T�0��_�Y�115Ί\[͙$.:r\~C��4S�E8�smYŴ�zlKY����B�qg�"������
P �_��V��A- "�����R�<>�yU�eM�i�G&"K#X���"T�"|s}�bFﵕN��t����o�Re��E-��0��p;���a�����ci�<���R���T��;�{�x��h��`�
�<���Y�ܢz�I�V{n�m�?-9�t�����ɞ}�}Ih@[�ׁm@��]"��j>�cY�,�����y�F�W=������+�s���64(��F�y�Ծqv��כ�.�d3⟨����0/��}�vF��RI��O\\"ۡYtT����Q������q�5,��_-Џ�B�j�
K���}%����̫�]���C����MaZ|�^���"jr�lSsi��b�QM?���'��Vk�ܘ����X~����g�"���$����a~o�����ȗ�� ��lZ�p}[?�A�b��bʳz� c/UA�߄wj���n���,v�Zc$#?�$��"���4
aUP���fK��Yb�]���Խ���-`�����Y�G]�6⤜���"`;�����qBI���d��OVc&�	�J����Ff�Wr2Y]::'z=(o|�
v�Z�5!R5BN�(nBJʚ�Z?[�k�!��Rh�쏁�UP���&Wj�v�Cu�Ɖ#�^�X^��[�B���3��_9%�N�Fv�S$ѐ���(珡NW��r����&M�>{�t���k!B�j�<{�Q̹��>�E���������_����� eZ]��f��i�0�C�jR��4�62���p�!��BƔ���"���Z�[Y�Ǥ)�J��(p���͝e v@��W��f�n�<ke���A颖��D��X=w�>����h����¦�΂��~=@U���菘�G�������Y�.j�ܪ��uAN6��4�a�Zޅ\��r1_��5�1�o��|E��B��[���N2,��;�	6^l������ɒ7
�4ys��]%�8!��H�\�0l�%�V�����-�
�Z���c�ȴwfO.:�7��:�-��Y�MRx�{p=������v�I�'FԷZ�,x�esړhE(G\�h���D����k���J:����y�!�]���n 9~<�i�B#0�U^T�����	f��5O�Y��mV�QCI�ۥr��C�2���G���A��tR�����oޠoӈ�E�F�c���qAIՇz�W6�tj=�G�lVVg~rd��Z|�\Q��GB�a5Ls�y2���С(�ݷk-}!m[��#�5F��)Y�j(����vp��w@D���鐒�'��[֓�02�Rp�V� ?�f&<�0�I��H'�׉3_S��:x)ޛ���S��"u+pR_���*@�1��J��;�o?h�#H��.ZOf�)�5�^���i�+�z�4�5�?�������hx�h����=˷a@{�r҂J2iȋ�������d-LI�l��-,�G^וp���GG㰏������X�Ƞ�'M���,P�~6���,��n=wj?v��Ѧ4d��Q�O����������s������l$��� ���M5ُ&;��.2a�4]��'�u���*N�Gx���:R<h!�"��7�D1�O������}?'�0҈Ы�<����M�E������(�* vc���)�o�!�{ȗ��R	[C�9�Ť-#��y�%��/�h�ր|��u�ΩF�=t�[�s�d�������M�m��5��]u������`����|��ʑnJC�*�7�r2ī�v��PZ�����%M���H�'܀���E]�	>j=��ѕSN�!�؜�Q2)�?���f>�̐��I��I����YO�[E�-��� H���S^'��븩�m�k�C����n+���g(�^���{���[��;o�)��'|ڥgx�o�p��BoѨ %��7����W�D3������9����+�h�1V�g��jT�xܐ-Z�����QۺWS��=�)���-��<�8�7ʂ�g'�g�����v���w2��I�T��ޫ�~�3dhۭN`d�<����UV� ȇL؆���"�)H���S��!�P�$�L�ǃ� �tOrls�8�_��gxc�<�$���3kD�W*����i-�gtk����ķl��QG�.�Dө�q䔜,�z.�w���{k W�8'��kҌ��}��#��&F0��`���pX�`턭x����}E\D���������tԖtnG
�Pb��N��i��1�G�����ؤK"��.�/�f7&�O~<�Y��3u�V��5�U�S������������*+-�t�b�ȡ�fЛ�z�c;>�پ�!������,2��K*�*f�<w����V�2�+sъ�����ք4��\�r�ݹ�EP�Ƒ^�P�,�6E2��c�Z���ċX����!C<`�/��{�U������Mm�6F�����Z�l�����6$�u����3��}0@9��k�u��{{�606Fҗ�{��^͏�z�6V�Y�5�s�� �B�����.
�n5f���%-�4SMW&����������<+������,V gC�X�v�����>g}�ll3\���΁6]+����m�7�Os�R���<�w�˰K�9��7��\�&��VbLہG7�d�.���Ɉ��~в��4�nJ�;`�{���� �5�x�N���D@ؑ� �^<�}�
��ly����[0���-��F�P��'�[	�n?5C�D�U �±GdpN��c$�z�e,�=m�aE�θu0�-�c�����&7�"j����EFL���v�q�r*x��ZO��?���,��J+�%�ȨI�k��d �,��������~��f\�z���*��y���MO4� ��}�xT�x�cz�h�pI��hm����|��)n�J���wY4�fND��؂�O���M?��zY�ֱc�<n��&|�é��$>����gѱ�h͍��qeS K-�'^�u��08&�!wfT��}*���F��P7ġ�:n�$�ϰ�/8�	����0l/���_J��9*!���
�]F]���%�p"�q����y�Rm/����t)�.�2�"^2�ܔ� �Z+���e�����s���gY��?D��gì�`>,�9I��`g7�E=�D���D�9"�A�Tv�Tg9G8�=�%|��F���rQ�<��~v�����Dǟs:���M���6��$j[ُ�`�+o�3���Y�lS�"�T��OP�xb�!άk�x6��rl��k���ӽ�@��w���ܶv��o���3B	��Pޭ��{q�l%� U�n���ڡ4��+N�+�e�Ɏv@��3!����`�JܰD`~wpH�m��@�����e�{�v�$a/ w5 ��Dy�Z�o7)]�$ۑ����;4�?,�ZP��20�KF.mFN�W̴m'1���'��b�q�?9�F�>޸}h�>��@�^7�����+��LI�U�n�?���@F��P�}\ȭ!����MS04w��ߊ|�w�70˼��֧n��	7z<��P:�8����7�
\}�R���1��.��]@�VF(@�e�w����X�����+�3�L�1Է�G��F��[f���Da���i(�k��>))/�"N�����Ӟ�-8��#��0�1K����%�1�{$�e������ιBkK����r�O<(� +b$TD�+�n�W1���Z�W���s�jtKz�G�r�f���0A01:ӒP@�,�qH�u�ج���b�FT�ڥ��;qՒ�W���\�T��^8�{S��Џ��&��|��a�r�����rh�~y�F�I��i>����Ѫ]؁�O�=���� AY%z���cE���9�#F�$��W�@�P�%B����孆�[���:�֡@�e%>�wV�"�.a�!������x�i�$,�F^)�W�Z[zK��u�].��c-���ήt�.�7.����R+8�H\�n8�����FiT�<(x4��cK,��l/�L����1'R�󬖘v4L�R
��kf}P����V"�>x�"�R�V�G��:6<�u����W��C?q\�T�8~��`Qn\*�^H�ak�</۬``��ںb��CJ�م|��)c#/����Y�Ԟ�/k���n�^���>�c�)Z7�anI&�i��±W�Wd(~lX�B�:`�sv�t\z�CZ���׶�*&�rH0~X�i�}���i��R"=4���V:QG���P�VXpޏ�B^��M٠�J�HA~��9��7[Q�Q&`���_c���l�:�j��OgҟN�����C�B�'�Ysq��՗��50�جqy����!)����Ă�Z8zA��A��@b�z��4{���.1}�}��v�Nⵢ�5�[�&�]���'W�۰�yj�j��r�'<N���뢪!JP�6^��۴e�����a��>#Uk�#x��E������W��,#�OA����,�Hk�w��π���.Iq��(�TR����{eB,1�&�y[��w��,��ݏ~��je������#E�k݇��1w.G}.϶&-�1����'x�Ae��l? f4��*��9��,�?��)��>df�c�<�e
�n�<#P�>���4Ҷ��<%f��̹�v<��Qw�<��O��5r	vd\�M�Gj���vif,6V�_L�n~ʐ�&xTNS�=வ?�w����o�Z|XVc����3����֐^�8VR2�-��[�m����ᛧ������:�E��%��-ϳ,��(�Fs@�_I��򎜂'�M��n���Η��p�\�5~�g}��f<�*n�{�}M����D�\���y|��e��
�F@O���T�QF����>��IPFI/����1xRDQY�5P��[ʸ���^6����q�J��A�Zl"T��>f7��_	6���sR�Ge\�D&�YjC��	�Fa��%��MG�_I�wP�q'h�pfw˟�*��U԰����Q�me܅�+5��2�&a:�29����'V�@\���DP�gֲ ����׃�(��*���_�!��B�.�w�=M�����4�o}�L�z���p;A��k�O�To������C��� �»}��스d� �ԈM#�m�6&�3}M .@jR��T�Չ|2�dI��r�(���u��
�8ޏ�v�ѷ�Y��e�)E�����컟fЈ[N�p5�5(��Hx;j�>���g�\TU�6.��6�A�����ZR��?}�B���_
����N?x�2|-���-TU鿳��j�~b������)�mCw�z���$�o�XIWc}Ʃ[����޽:�v���ϖ��c���7I�7����>>7f!���=��|�\)|��&��2�n����
\ H��~��^�ϫ#p�ː!�K�^��\��dz� 7�,v�q|���N��y(������^~�|3��[J&n�1sq\ g�h�l\��>@��ǣ��{�,�eHR�M@��;ÎG�MC��0�}I�[S.ն�u~YJ/Gf���_vTg�3�:	S!Dyѧi�K�!���	���z�o��#$-D�2]�m:H��5�~��(�;T��8<��Եj������0(��ʔR���ț8Q�G���/�p�bS�ՒZI!�T�����/u���#�| f�x_�����:E��>��1���}% �"��MR�.��;D&�_��̭��g�&ꤻH���ƫ����/�_@�����,o;,���G�/�	:F�ü�HC��$��m���Sh�g�r�4�>0m.�c�T����pD+��N,ȉxQ���؈|׷W!�#D]Qn�,�~< ��B�|N��F�ƙC# �̔@/0��v"�*%�5b��s�ߜ��'"ԙ����{��t�;
a�\Xo
K�o�d���0 ����D��O�i�!�3�{A��V	���f�Ku�1�"��u�`�{#���Z��Q������Vs�u��u��qޡ]�BIr�s/���M��6�����C���q*��Q�����l�߷��������;�V�9���Es}��n��Lo+�TG��-�W��_ͱ��]�i�Pn�`�����;X�_|3�k�2WCg�s���E��2ç=��e'C:!/��Af�Bȳ��L�\�W.�� Vh��b�	�����fу!3'&����K�gkZ����ℸO��؄Df>U��n������Ԇ��M���XbE�j{ʃQ]�WR�x̘�'���vK$��x)��[,�p�A 8�a,�)�����v���g|������+2}\�F���%��l��%����-�W���M�	�^���ސ�~�/v�A�����΄U�VeG���Q	Q�9�󙍆ۙ�!���Pmg�;�e�Q��m2��f�ŗ���@st@���k1�w�n�xk}&�e0��8e�f�u�)gKl�M�j�=�`�/!�gT=����Pq�'��ڥ����f�Xf��q�|�U^Ϣ��zle9Y8JF�n�"�U�B�a[*4:��uP����)J13����}7��
��qf��n[&������q�
5^��.;��s�n�����5W�Ʒ�W���mL�t��c����@��9��i<�wq\�����T`�	;�戡lSE3�_�.A���V�!@������Vs�X�=�0R>e���}�<�̯� Jg��(�Ʊ?>4}��]��W�83и����w_��J�ư�Y-�m~R�N�<�5��z�QS�|J[qH�rw� ����gY"��BE
Y�~�0�Ǫ��	��5�aCz���v�hh�r��&�=�7��uc������3'>����L��@�����4����f����E�Y�����d�����ⳜE@��6��1��0�v��x���s\�Z�$��%q�����d�r����#�QU ͗��\���J5t(LD��$���
h��n��:*����W`���v�!iEh�6҆:,�Z��g����n¯I�?�ڕ�����ՁqooU��(�ԙV�qG�9� ��<��da�L�����/5��.1껺Pl���L�ivz����[��������-LD���	�y%����0uG�#īb>l91���՝�E.D�J���M.E�"+���hktW+�a��:6��[^ ��>G�Շ5��Vl@CU�c�J��S�&l��=!Ѕ��>7U�/���:�R.`�x�D���93�yH�N�*��%����>��N���� �>4u�v�h�f�DX�����.�I@��l�dU�4| nB"����}�lB��N CDkvlpb<\pI����fo(� sf=~.���Sx7��M�x����7_�ZY�:5~����[��Y1��`+5�H-����o���<b?`�B٤ee�H��Ï9$x�K�9�8k�/p�V��֌���`�h&'Z@�6����B�̈�CB;�c�^ʭF�Qb"`|d9@�G�,R��#�c0�#[%l��n���E�
��(.XI�i�7VX��N9=/� I��{��L�e^S�{g�ݯHW0V>y�닿�q��
hP����]_UeG��5����$"��lM���DY��))���#�=S�*��_P���4�z��<]F�w��d\�z�Ȣ��*�Q!U�=�!��x�7�]d�ʠ	ht�o'��0�n�z+I�#b�p�)��m�jl����p��M��B�$b-�j�6�§g�!�Rz�a���P�ө�<p��O�����N���զ.����Q��	����Ի�l��ƣ�{�ȏ���-�`j=�����=[��6������n'R��}9E_�f3�9�BBtcmr�^�c8���Z]��e=����i����E*@�T>Wǎ����AX��
N��{C�_��H%�>��Bէ����?��ZG���؆�vt�j+%�oc���X��5�K$��,wcu��|������MHu�묨`��oW����&	C�0�ay���t��V���g���Bq8��6|�*��[
,����96�H"Gݧ2ZX�$Pޥк|rR����E2L�wi"fU� ��A�r
��w	�t��-�r���BC`N��"��[gkq!�}�:β�����6�S��`!�G�^����ؕA�:g46�0>X�d��J�:�t��zșLm�1%X�B����xQ{[8i)�k6O3*O�A�%4�g1c�A�hb=�x��(駔S`�h�ͅ0vh�*���D"�m0���\<�A�օq������#I��f��]y��6vxZ2͉Dխ����di�l�9ȗ�l�W��1\�xW|�+J�]��7;#�ф���E�}� ��\(��Ϋ���8�'�K\�[��=�o��&��;4��4�{}]�r�PD�`-J�q:�6�n-J�p���٘�M��9��u̲"L�߭5V��Y#lO<89�-�>��խ�K�C�z�/	L���5j��4s 	�'�B���� ����hR�R�����ݢ���%��z��uY8�MT�*<6;�.����+��;��η��9�}�i�Cr�fg(���aq����|1�c�O��j��%Ls�gc�8���)�k>&����FK{h+gn�Iiy�sȒ���p���h���K�q����N2~�?K�% Ѓn����<^�C��U3���;���'���U|8qe��382�/f���x���A`��%���T4^��BG��!��U��D`~�ݿK���'ic?��Ԭ�+��
��.ә�ʮ�£՘#ɌO�,�<]X�w!�9LT�R��&�;T�:Oo�
���������cdJ�F5NU�7�� �[�
���~�2\�H����d�	K�b�c�s>f\��5g��v�V�7�Z����~�V_��.���!��]k�4�Qׂ��TTv�{ܡ6��iE*���6����E�1�d����[�	�N����]�@6�U7�BB� �,�.BiA�O� s�RN=���g�d��f�h]��j��.Gj7 XP˺&G�Y'����^�'D���YQ�n>��ry"�:P��ωM�p`�s���ͭb�R"�2��G�����J����3�u�:�%AC������ǹp�7l���=�f���]�)�h3�b���ԫ�X�`�	Z�D��添!R/�DF~�&���
�F��x����Om�oݭ�N�ݬD��%��0d3˟3�H-�����V���t�V3�$پ�ۗQ�B�%[�|���̧�[>j�}������HY���V��Im��U��O�r7o�B]Cdcn�q�S�H(��Yj+�*s,CAQ�Mv�з�]��(�P]Ɵ�ַ�d��pR_�t�-�l�@L���0I��'	G�ұ�g�s��?�j �	L����:q�DL��bV�;gdB�$6"���Dd���q�@���r=� �`a�M5�m�M�<hѪ�t�l�� �.W�6f�Lm:$a�Фw͋��3��Ѿ��Qk�Sy�}�����4����P�x��!����O��\Ȇ�f^�Iq஦
]�Fh^T�]R|?֏�Q�LF
������4�E�P�0D&�s1;��j��L�s�#n��t֙:�U]kK�z{ ��Z"&
?b�x�OU�Z�^��%�FX�#K�I���
�G�њ|ڟ�����ӧ�נ�ZA���z�o��S
�B*b\M�Oc�`�����t��=66ȫg�8�ۯ���ө��3�Yq�
h7Ť�i�ۇʝK�}ޓ���X�& �$�:T�tR/�Gs�aZZ��!��R4������8�}7�\�UXĥ}�ӕǙ��|�M��=q\C��w��?q������΃l*S �)�l�Y�t�̽S��䒅�A�MK�#U�}TԔQ䲸�{&�y¿ηl��0~���`a9pd�y\s��%�t'���_���A-g��Uj�Bչ�e��ҊF��7��U4��ܝ������iV~1��v��e���?�2���*Zc/��(�SnuI�{�����C@�n�F�~31&W�5�<�D��?C����#���cﭾ	H!E�b�z\dM��2&�(G�y;�ͩ9#��H��G�*��V�v�L��	4���r4v_;��b��o�I]g	I7�&.	��ĐRI>�l�>Br�6���n֭��f��Z�����X�.J��!����>O7`JҠ]˸�>��W�U��/X%���Aŏ�3��SuR���P�UQfb�p��dmͫ�:�E����r�4Ep�8��A^p_��a�~&����i�
�n�N�|}���eF�٨���vB����5�#�m���}�Q�?���8=�n�d�����6+p*��Yw���r
-R�=#�sz�H;�N6��H�=o��c+QgYe��|>�.��aԥm��פ<��`�]�I��,AH��ո�&�g�WS2_´X�]�z`Ϥ}���]��Ov�rsՎQG����*��/n����2�;C-���TD�Oӫ����G�55�&B���k�1�_�LNv���*�լ��gEI5���6��muS�PB�N~�Vݵ6�$�����8�$�X�R��eRZ��H9Hă��R�OTfb�8����N����U�F�6n�;9d���:ū/~���t�5��X�iGRAi"����p��U��x�K����tV������r���� ��:Bu@�D�ws��X󎰋�y��Y���;�2��Cz����f����3��ܫ�)bHvbY��7>�N�:����W��9i)3�"**���� :��5�juD��Y|I~ϹG�d��	��sR�F�%� "Y���7<��^���s�v�w9������1lx�~����%�퓍ZFkP�ZLe��D�A�ЦY8بQ����xH�3��v{��GY�lhøAy�8�B��O�����'�K	����=ՔJ@���p�6��K��N���g�h_��g��'3�nɍ��^�>o�Esӯ@��YϏ���zg�p�����
�&��E��,����KU�T>q��m>K|��'�M���%_C$:��
������a'�d�Dö�5�"��	�������<-�r�	1��zↄ!k�9��W�F��t �=�n�Ĺ5{��rM�K����!7 ��Nc������x:��� �@�F�U<�-q�ADu�z�>�{�൐����I�/r-�!1��`	ƀ�H�#�S�l�_������=�i�����"S�	Aj������>�''{���gY�H�jH<�����>f/	��XfI>u�)�J*�#�zh�I���:� ��1�R��1K��t�6��\�R@�(�D�DI������	m�1y2m U+���<���c�|���x��ȩ
Q�
�GQ�"��z�N-���wQ���rsV�Ya��v�8
T/��HJ�AB��\̤L./ӓ���>�mBQ�k�%4���1<�N��v�X�è||�O��P�E�N.�ԙ�p���k��2cG=���[B0�_TO��; :�/p�g1P����?�]�m�v���~Mn���Q'Y�e*�[���Dk�e����6L>�5��=P�%�u!���ešclp�ѐ�����bvUm!�E0��,��qJF�����ܹ�ZQ%i.�䥥�(�c�~��_q��%�����g(�I37sݟ���MY�e�x%���cK��V$�^E�9p�P��47@�B��'�{�]#��>8���Ô�W6���Ff'6��X$���!�	!r؉���Rܷk^�[|���H��y 7f�H���G���)����������CD7!�'��X�Nʟ��^tV�@����`�2R�g;\��M\����������X�����D
ذ9��
�ڒ��jW@<�SN˿扙ME�*�u�]	��hlc ngh�<��zL%�4���?TjS3��]'�'X�!�Պ��:?rb{�EA��O�b�<�0�#�Z���@=aJ�=�}��A��3�*w,�i<qqe�W�!O��Z�����q^� 哩c����Ѥ?�}���?J|���V�����-��{����lc_a�OF��ϙY�"aT�eڞo��c�[(E�L!1� & ٪m�jPlm�#pU��u����)��G]:B��ix�x8v��y�t�=��0ւ�]��g ��&�J��;P;4����V�O4�q�E�i"j�~���ѹͩ���?R)cفp�^v���&�W�O�̣B c�%��.��xT������E���4�Hu2�31����R���ui�E�
X3����{
�^�h8't��U��.ay�m�>�v{ZEy7��;��v����m�&� $.�U�[K�n
XCaA��>��w���v3�������`&�aUR.�����ސ!Ip�:�.�B�L��,nJ��{��$7@��&�_�#���*�}	�h���hJ��,���)F8jB���I?�<��������$? ��d �3�(�d��Tc>ԯsw�ہogwN:��Tu�r�k�@������C���ǊL�kbv��_e�Z�&���WY������gI:�V_M�h�'�ݷ�u#���Ңu�6ޡ��{o��X@ωغ�w �I�^���|׉s���b�5��7�>���5�ӽ*(y�n���` 1Y9��1_��A�`�gJX��â�qDT��a�i�1��MMv�f�?iO�:�A(/`��V#CE����aF1�?]=ƅ���nW�K��CݻQf����QҐ�J���K��9�0�3p#�q@;���vE��G���mq`���?� ��q���Ӽ�4�$.#yEo�d��Ѫt���ޖ%�CPd0
�󚀷㪧���8����j�)_�e73��,�|T�l�Wv�7�hӥ�0 �83�M�D�N,:���[Tŀ�/|��ȑ԰̈�?��1H]8���~� ��j�Q+启��3�]p׉�up0�)7��a5M���A@��P	}ͻÚ��ii��z�`�k5{19����6��=�^�jYX/�T��`R�	�>�rL&ƈA[98R���
�^�%�':,�����"���CA �xףjfl�
�8�Q!�]�� �t���{�&�ΰlĀ���L>��	{Μ�,����âR=��~Cb:�v�U���5��x�CN�q�rs^R��,��r��cp�4����Ǩ��Ф;������̒+O~ֱ�9g���(����K�	�������o����1&#���_)䱭�q�h��nY�������9w��^"%iI)*�|�m�X�'�4��ש���7��^A�'[ۛ�a�po4�j�f|�x����i:�>�-��׬M`&�WऎyeKO��M7���dKtIRSJi|�k"D��Sٻq7Ÿ�B�<� On��"�tsD�$�]m�-V�9�y�AB�~��ˣ�O
tVez�R3��#����!� ?���bv��JW�=b��v�<i��V(�>���j�2A/��[-O�,FX7�+�7x�/�9��}�8�9�u�[]}��ڍ�U8����r�o�q�5��/t�9��j�rvHg����E=9|=7f[qz���:�IA�?/J �&��m����:4��O!��%r���U�nȉ�c���{4V�(����\��޹|iPY�!���(zɴ�X�G��r�l���oP�5�ڎ�W�48d�Ge����6F��ǦF����O�J�l R�Z�$��+n|2��R��5��׶}�񻴮5峯� za�t^���KF60���N�O#��ZH�2`���Γ�x�nғUa�)�6ïŋ�6�g����n���W�r�Il*1��`���i^<�(ŧ�!g�\Se���G>Z)����<l�1ʿ��(��ی���og�p��f\������
0���[f�Ɠ��0�k��\[Ք!0s	�@����?��|�͎>����s�?���\�:Mv�p�~ s��tw�d��fφY���U]���f�Z�\��"��8�C���6�O�[��������]5�~�1��J����P�sm@��K\Xd�}�P*#���N��Ѧ�f ��gi�N�i����ZD.�. ��K�GpKa���3��o�]Iy:��MN���Z�0A��t&t�^���4�`�����ʯL�'Fnc5�yN�&�r=�غ��(3�,	8�03�_O�
����ڭ;�(����=14g.�B��>.���S�7�B�y*��Qf�����hH�:��	�<�t�:M ����nx���+CSYC��n2���|��lJ\<ة:΢-��SI�u��P"�����;h�3��c���ϻd��GJ�y�)�=�_�q��/�Ք�VS1���?�����!?{zk�<gYC+�����1OU��K0'�h�E(:�j�����6G���P50�x�T���H7�q��&_ [�L7�O��W�=�쟢P�6��a=��e�����OLxJf��,��ӂ��JN�Sq���A��51�*��=a(�X��3=��u��'���/�>���w[-�m��p��?�-&�%��r��B����W�C���S^��}��t�n�;-�(2>���5A�⭂5���訆��Y�yp�#�ՠꙞ���`4��<%��m�K�d��½g��`H*��h�!���I����BoT��2�%5�\$R�oBf)+S�����T�_�~����ۻ_MY5��-��C8��Q��-��k�n�mPg[S�e�V��Dh]���v����J�M4e-��k8Y���^�Ck�̬�ø�����~#��Y��C���9|���7�W��4d�5#��l����	�=K�Q��h>wʦ�ɜ�:1 ��%P������D
g�c4�{g�������(��.�����<�<����5�i�9M���
h�A{"=ڶC),y��c��/\����ĶX Oay7�E͟��� �A
v���b�ɨ�V򢜀S��IJ��@�xyҾ����Տ��#����<���<�Z����Y��1�v�k��YP!���20�����=]��	ؓK�͠	l/#��IX���Oz�|.�hG�}_�U���"EJ����'�W�<O�pw'B� �I�	Թ��m%R@��@�u����m��[��������8�|��u�0�x]Ws�'�(w{��:`Le�	�u��^�����r�ȳs[�y������5��g|ɋ���i8AX��@��k7�*��ǃ�d0a�&!�du�MG�[�d���k�a̤����]�؁�n8bZ��׻�T~W13n}7O��"p\�G'G���}��)��i��~�a.�_}�H�:e�� �V��m[���O��dX�x���.*tdS�
R�o�5�&%����f��%G;�Gz��Y٘�䢈��l�sMWSڿ'��G�LM��P�.BcT�m���Uo��<RGU�2�G�v����$}�Н��*�B�=������ĂK �y�|�!V����&�r�������$w�y�Q�IL��pv!1�����U��z���2҅; qrE���r^�|�6�~E��'D �T���8���=�P��[�6�*w�45$� ����}[(�8�
�*q"{`��$�|��`�ǔ�f�1��vN㆔����J�ɶ2+�y�wf��!��NcG.֊�<��z~�2�9�ڧ���.�1��	��_p�X�����b�<��a�}iC��R�
uh�K��$TTf7?�S<���L�y*�!~H������Ģ ���"M�]fz�=mY�#��<��+L�l����0��څ'�=_��8 L�7�v���Km��zV.�+�K�u#6����������a�4=Y�,I��t_Pql�=����F���#,�{�w�P�V�y~����u� �r g�� M%����gޅ��X�g�-iA,�Q�nq�e6i��Zͥ ���)���6^��?P���P���D�F���z���%��=�ww��")ގ����le�_ U�|S����";���ȼ.�v���iRKwf��9R̖�f[2��R����%�/Tr�M}v��tN�f�W	����@c,���,e�y 7�OJ�����Ve��:�{�ju-
����5�kˠ�e,�P�����D�{��2� �/дT�	��n �`��]NU��{�v,3r[�6��O�^��bZ$eRH�)�����21.���2�8Y8�^Zgӣ�'*��Dc
��v͒nKSJ/����O��_j=IU:<��{��i�������SG��{Z&�J1Y��c��`ޫ�7k�xr3b 8�	լ�R��>|�P�z�{�esb�?��S�ݑţ���*x�kdXp���w!K�46u��H��w��2�/(~�R���wZ���m`��΂��]�'�>�������L��!=��/�P����v�r�>�[�sJ���_�e7ƫz��8���H8E��i� f���>msi@���"��ӧ�i�V�T�1�ЈX $q���|q�ݐq��ވ�p�I�W�|f���A[ƙ��ց+u�&�9~��B�շ���"l��&���J�����S��iHM2� ������0v{,���as�wN��hdxo��2�[<O2S.�����+;~�x�M�b,�U�* A��W����E�&F�Kw�����ͯ$������&[^c�k����Y�3GWd���1���A��Fu,_�<��|O42�ؤw�G͎����ϒč��wW
��G]�Ӯ�N7bF!︁�od`eĀ:p�!��k2s;/�KH�j��\���L�GY�',�P��ֵ^���݇��׀K"��� p���/q.,W:�f����ZW1��*#�nW��<bΒ/7�߲x��)��Vr�R��~{�H�_�Nxw4T}��+*`k��w�%<u+y�Co��#����y��.���6Qݴ8B	n���y�00ę���Гd�QA(�=�@��D z�C�"j��ך-d�*��Y�w-QS�EiSwep��p�si���q��[�,2��b��_�x��jD��qo.�/m�f�Z��b-oYW�g���d©�7P�z�B�`U��ۑ�w
�S�{��G������_]<}9ɑ]�ww��:u�*�(�Xc�iW`ii=�H.��b�����ӯ���Y�.��p��'�:7T�$�5q����aG�{/Ǔ�.��J!Q�`��"�>��Q�%�<3���yG���nO{���c���7D+t��e|7�Q�a��E�l=VzOM%N��Gwn��w�W�Sl�<|M4=��ʣWOM��Vki�[�F�v��)3�8�UKW�!mMtn�� ����t��2��,�aƍ���y$���=��hLӅ��6�����'������A�*Na�����6G��`��������cH�~ �����\Fݷp�Ŝ`�ʒ�>q&�%f�q��,*���ƚt�"nh�Q:���uY�D��U�䂢%�;H՘�|an��5g��W�����X�{�#/�S�=�it�?�iT�2g��ȑ2_�fk(@�+%Y���7U�ڝ��)���T�O2�,Y�+�3hk�|�͡_ڋ�:qo���/���<^��������S=51Bo:~l�k��X�hU~C�����Am��u�&'�[��y׃�Q�	)q{Q���d��M[��ֱ�%ɕUz"�<G2]�wh`@��H��P(�W���0g8	���R���6݋�*Pj�{m���苟�Es]��rj0.Ì��p*��"�@�j�]�G6>R��P��k��	�G���?� �F��n��-`jŖ�pf����$�5�I��3)���t�j�"�m��lyv݉�}���~�uϗ�,%փ�:?���Y<Qtn�q��s�4kb�J����6c��	�>ɢO����� ,"�b�����@���aUX恵�4\�1_L�r�#E��ܛ�c~z`�7�4�G��e���T�g������Q��~�_���ϻ����g.��z�9xݟ~�4���V&��t\�r�gm)��ɫOiJ�M�(~�ӹM�~�[�q���#��I��R���,���g�Y(L��UVV��}���(~��~�'O���.��F{i%�>4�,M�ʹ0"���Ǘnp5�I;��9�հ���od=�
~�~��_��+QD��Td�:����Nr���1d�_�(�`�c���^�90�랄�%yb]�L����Q\�\�/�|�o>(�h���:j��(c�.�Dۼq�5`�홢��"	�O�H�p�Y��o�����<o���APF����3��M�Ib�Ro��VV;�T�e{Ut<�����~{l&��^ǜ�/46u��j�>���톙s�%U݆,a ��)N��`�����n[�q�x�x$K�RTT�p��cb��.í�!4Q����%�Nr\�0�q0#k��NcNR�#CϾh�M��	A[#�O@Y��+_�<_���Zc���o����ꯦ��i�����fbp{"��zt��C9�����Nt��rH�뙟�S`h��r;��_��	���g�\Y�4_�l�yV���@C��N߼1K�I�$qP�'�D7W�!Z��`�����wA�<�,4�#�uA��J�)}��*��k���yA5=)^�*�}<�n
�٫��M�㴕l���L���2c���&�ɇ7[��g�fX��/pú ���b3Za%Q_eA=OC�pH�f��Տhl�mW��]p|�:c�%������� ��]��Ou��b�o�ef��h���i=
,���OФ'��X�
�|���s�n��b���B��{p �H�d���Q��"��i7��r�=^H,u@�/|�&.�h�4W�{�P$
�r�3�9�k�8�P������M�:^5��S��B/S���`Dh�悡ڒJ���Fn�����u����SUx����	;)s"�Y/H��M� Ή�t�����(:�p�dym��Q%@r�F��nB� �BVh�f��8��G>���Jb�0܀nӢq"��ID�P�Ȼ0��{�v1�G���%/�j�g / ��I�d�Fr��H���B���W�R���J�֕F���)kK�>�T����͐��<>���I���6���J�фX�_9�C��&Y��_�9�2U����5��pD�[uE���#�,����. �
*b���;���I�
:s�ٕ����l4m�*CFO��ˍ2�Q�]�cw����G� j��,ñU�ӿ/9e�-�<�K���g�,�e�.�zTh3�f.꾌R�B9��B����Uu�F�+Y�����& QW~���}�?�jS4
��C�M
���"�´�V��yr�3��N��&֛���F�ٻ��z�*��pYb1�����U���b=q�������Xџ��k��}A�1R���EE\scs�ynVS|���#�[AS����<{�TV�^�7�^���`�Mo�϶N��w8A��M�#�����L��\�:l�먘t�na}��9j��|Sn�t��x�ؗ�ag8�Ȩ���tp�ާ6p?�Yh e#�p?	���=�c0?�H����_EQ2 կ���)>��<(��:EHxmc����]G�����#u�p��_vijPϛ�U"����C�>U�l=��02s_��
;�>�=,�FP[��s%c!C�n�m�e1Ø6����ą����0`W�?Aa�/�}�}��!PFJy�!u��[���3yuBO��������޲�t��3�YI����{Z�c�&�n��� YqO����:�P��N�lI��Mv­��L��� d��<����{ků��ut��ףa�s�c�=8�������6;.�\X�ε�2Ye+��a!ч��q�v���@��C�+�0%���2��$g�,�̬��@v�~�}8G��,�n��3k}�3�>D&9,�������cZ@D-?)�=���S+Q�O'�O�%�M�EZ�b`a���t*l�F�_�A�<�)9@�H
6A�rP%fg�mXʽuh�^É��ۚ��>�R�e��c���x�Q3�3��L΄���M���q�҂!�4$u7��e���T�.�Ԇ��J�� � �P4�٬�ペ���&���#������wۉ���߼����jMf͝��2]_�ʂE��Ò���ld���0D�G��A��J[v���Jئ��"�X�Y{M~�t��s�Ѭ��Wđ�?�����&_Z`W���B�z��&�l��:XPd[1W9���dm��b�ڷkbpDI�j�>�a� �.��Q���c,�"�y�v>k���H_�3���$��;���<-S�ؒ C���H����(`=�V���?q��q�TL����R1BF��,�}�G��c�u��@���_b�κ��6�w�G�uĔu��H�~���˅$Ba0OV�c�!���tzE[#���j�
v��|��I�[
q2�O7��ʉxeTL9���&���`HNl/��C�^�|#�~����#9[{S�vGG!f/]�i�dN���z~��c �٭�?� Y���7���N4��#���8�;��#��6om@C�r��1|{� ��!�m�m�B�Y-/3��+���iD�.��0Jy7F��˺�x��4gT�P#F��z����e|+@t����T�2�[�\6�uzg�b&f��D���1S�[��*ND�&��kgoT7|�����@�M�G՛n.x�Q�>��@���][/Z���$�d0᛺C�.�R�#2��ѯ_V�YL/K�㱂������!�cY��ڝE�I����ZW܀���
X���+���\j��ܘl���f�������Μ4T��j9N�yJ��L-�'TYҴ��a�r����3�]>������kM��5d�����d~�&K#�X /�ƞu��͖S�0
�f�mR�&��j�,ũ����h��<���[ڵ',�2`��F"!`a��p�����+�o5@r�.j"6�`���LY�K���T�îe���$/5�3�X�q��gA�&ۦɄ�,0�>�aT��.�kOe�����zX�tX�}�=4js�y�!�0h���.G(��)�j9�:�?�7c�5�s,�	���k�>�����HX*^�GuH;�]��C|�A�O��%P�j'�LT��!��r�!�0� ���3�ϛ;G��[� ̧�imTk�v*�������������7&G�P�-�Xr�'3δ��|Be��D߿ґ�����#gr)��E�d�֫\��v�#��H�,L��O���nu.s�qzn��=�(��3[!\��M4�G�kr�f�$����2��\3����~�?|L��*�1��H۟��,>�:.�Cq�쎖�\_��,�mES��+��̌2@J&��fJ�����&�B�?�6X�G�P~����.KJW��@����#����]H$P5��*�մ�!H|5m�`���@��l��o霥���_ ��F�\�~�]'�>>[{����Rl���ݾ���I������z��YZ��T�q�W��j� t�*�������"�/�	�P	3)�ؼ���Hl�$�4��A�߆��l;�1����[��1���c8l�.�*���5t�	L�S��Ħi�w���A��П8����T ���;���"�Ͳ���eꉻY/�~D��X����*)u��w�0�Dۊ��\��O��Y_�T��E�5 �/D�VdS������x�7Q�i���li��%���S�_M����)��|�w���˓��e(��3&�}���	��xy�0�C�g�'G_���ڸ���5�q��p8�a񠎘ض��f(�T�9ik�A�U� EfF��J��)�3�\x����GXek6'K*��n8���R/f�"��i�#�KyJ���x� x�d��/٠�zK�97�v}�� BE�. fc��.����g��^�܊SP�Jk�$9*���"+�=��:!ޓt�c�A�bd�����R�%�t(�}��E���嚏�Qo2`
;+KL�2��N<^�i�W�(�*�8.�d�����F��l���A���3*�f�S�m'qaĂ�|&��9u��0��n{<�H�#��� ��J.5?饊5�
�%�g��_=�L����lϣ��+e��z9L#X×�P4�cϓ��-�ř_-Ģ-��*T�Ά�̶׆\��g��5m��%7$��zͯ.������Ye�	��8ϯ:o{�S�`�%�[�v҅}�[��H.�;y
�a 5�m�w�+0	rɛ,��`��d)� %�me�s��Ga�c6�롧Y�J�����:(��,���x_P�0n�E^2=��X*�,�[�rҫd�k
�j<{�3&�,�+HM��@�Fy!g.mW5銅�h�J_X�)c_���'߭��7!�;np�s�~`�1P�ͱ=�6��.b�P����x��Pb9��ףB��9W���u��x,C����,��b'ag[����ASşR��_� ��h�#��)3Bs&`���ȟy���
ͥ���k����x�7��Ze�5P�"��|]ǝ�L���ש��T}P���ۛ��rŉ�r��]7cR��A�C�^��:vE�)(Z��wz�-�D�~�>-�ߴb9�����ENk�	�ȇH�֗l����ٌ�C
2ǥE����*ȊȔ�U�\&�H���I$"�I��F5���-�D�au�Xs�VSZƺg-ӡ&V���r����Z��C�poˢ�����32��������S�΄M�~D��j��zB�������(�12'��L�\O
���Q�
4n
Ă�
z�	O��1fӾ�&^����!���r�3�SC������?��ٶ�>=�*'u�ʈ���?/�LӤ[�G���s��"^.E�*�&�D�/%����� �K'��(k�&���.��$ @'+1G�03�y��<wlF��8���aSN���]����Ӟ4�12��/X��rF��O[����tC��GQ�̈́�J��@���_HW������
G���&ЁF�ٻ4�#��mm���7�����z�4TQÉ�i�.!yT��E����2�ۿU�m����b��J���~Փ�0	��,�Kr
������$�#;��qݴA7�a��#�s5��C��C f��Ep���u�WB���x�m`����E��SȾ���)��D���:�&��h`0���y�u���VA'{������DȒ�ys��g�1#�j��E�w��e��j��7�G^�W��[�)܍vPFY#�$�:�g�. w(>t��f�}"a���C��?����(�c�nѷl��!J�U�Mz]~�zB�&ܮř��ޚ�l�s�ؘ��a˴�53d8 ��Z��Nz��r��1�H,~[����<�Y����hi,�?�5&�	0B8��Bu/���� �̀�	���������4޸N۩�|sr��$��ee[��¶�5�����,�'�Ke�x�(��<�ʣ]�q�tdjK|�}ש�: ��;3c��ں�9r�1���Rցu�Ein�TV��-�snD9� �/�">��XN_������gq��e��0G.�Q���?��pq��v�G�l@J��>?j�����
���3"�yء��<q�O,�0��kYT�K!E�nO�ɖ+�\�\��ܤ�ν���D����'�8�.�R�O������.QU0��m�A����� ����xf|�*T�'��Z��u��i$���&��'<e��y���.���? �l��;�y TF'�yK^��e<�R���4�C�e i�?1�M5�N��oVA��z�\)��^Gx�Z[��ij�
�b����cµ�!x(J�������*�̽$`K��!�+;���ssV�[�æ�&Sc�n��U'3���i�wN��f��f�.���#�����I`Ʒ>�y��nu4"!��1�����L�j���ɤ�;�7 ���w�`Y�<���*vɄ�U� ���4�l���f�d��'|� ._ƏɂХ'<��!��L�Pu�1OK�X"�T���)�%�x,@���t2V���?Rr�3T��`�0^E�̤���/N��`���h��
�k�ޥ�Z��&NJ�ӌ���_���U�.�H-�:Y���Q�p�o?q'�nL=��Y$>B�s��qS'�l�`ϊ�tV����"[�գ���������D�W�w�c����˿wV:�Y3�@~�W�{�p����p�z&�.fv�E���o��?F���!�ɋGpS�z�x::�y�|B�2�`&��j�]t��"�r� �@S2�$6����Ţsű��/Ir��f��b��1�"\s�.(��O�㝐���@�ڋ��đ_ j�)E!1�I>rD��H��ݣ�K�D/�3;U��4
��j��2�HRiu��-�a�	��\���67�l��֔-��n���Ӎ�	^?� ǹ������bKMx���������3V���s�����Sĝ����W����m^�DԝQe�Q+5�AKY4D����b���#�9<�N6܎���ѠI4MdTq�0��gå�;�5)�w��u��M�D8���K@��g�(�����!#v���A`:����!Y/?,?9*�2%z��5���&�3��������G̨Bo�W��;��E�+M��`}��Z�- Fx�gO��r� ���c�����k ����i�Y���1��9��?4�YgC�_��+�{����J��Ӳҽ0��;�����Ӛ���'����-ž[��&���Y��?W,��.��-?2�OĞf�㾤����e>]&��Ck&]O��^�(e>��7$,E��)�>�F9Z8+��D��
���9̝W���[*�nU�bBz��<2�V$ U[�Ŕ��2�������z�,�ܜ�̉*�
�p���4x2��]�Jx���&�HE ���$����t���- 1�����HA��a�y�S<I�����537k���vw�ͯ�?�����o	�ˢ�^��mT�>�v�"E��!<��j��ZO��^R�a��?�K@�[�Z���W�aoSԽ�����R��̡���ˠNݐ����Y����!~�J�$����M�Y��ԙ��[&�B���ױ�B�M9%�� r?�ɊN7�R��
B=S��v�����2t�.Vg<׶;���E`%2:5ҥ�<;���0/�[A�v,ܽf�m�HrV��R�b���m*��C�����!�������rT�������1t�Ź�x��=O��a���� �n$m��馠x������*%���%d&��B��@�7mH���G]D*xY��ؾ���56�a\/�DI�x*�<��e��PXd�|�M���Y�a�3�v�ǒ�������u.�zK�~�L�hI��/M��P~�p�@��^+���Y5xٶ�h��Z5�uj��}y�;�[ �گr�Q����&^�Բ!��K�i�T������T�0��n,z���!q�`���)M6�5����-K�1�����**�I�ұ�_zm�{�3�L�1�9�*�+e:Kc.V.��M��`Z�A/���ш�q<���y^o�C�_9��߰a�J�1�Q.���P*JY���N��Ît��X�{� �������K�-�ꕤs:}����������i�m-H�Z���#�#�Yy����eĔE��f,�ͺ� zY����7��ڠ��'��ىN�����0"��G�H�hf��H���r�a����
�7��8(���`�~�sȷ�k�P+�"pi�^�\�h��@놷*"��W��Ig����t�)�`qR��#�A�z#hq�g��dS�
<��#�i�0����QQ�� (�����#��w՗���C�Fu��s4��G�ypv�d��9ap�Du9�R��s��x�;΅�{tr><�쉩9OA�w�@,�u��T�\��"������g.Y�j�3���o���Yp|s�u��@b��J����k��p�Z,Ǎt�
����W����	�E���F�����Ɛ����(9�n���0<P���HRzd{��w,��5�.f�L����s����tv��|?��D*��1��9���ц��j��yu�4`(v�t����f���'���I�G�b��.&�� ��"%L"�r���gCn��˳�R�?�v��>Z��(�fJ+�*5�j?Pps��՚�_Qc�	p��
B��G���'��J3,ɫ���B�F8�RC���-��m����ax��bJ�%��o�#:j
^�!i�%j�7RN�0B��i�]�^�yaɕX��i���/H?�'<�fb	٩�%^7�ķ���9�!+�f��h� .qN�j�[�G��Ke��C[��ф�J����j�8�n�Q����BܖXⲔ�������<Qι(�a���llH`���<s���E���CIҨ��$�{�0-�3��[6.��tB�|s�>���ra7�1��]£Q��%����ڭ�oGW����ni��3��~x wh���m�&}�wl���,�Ҿ�G��Ig[�h��,S��;��s�19�Sc�V��u���wg�8s6p���Ϥ9�\�����Ƞ����z
��p��w��vp�ݢ�Ń��t/���o4j�eX(~ر�A�ˮ}PK�i�A{{�u�a+�2��n�����ï�:~z��́�t��:̓��p������R+�<?��~*N��C�����00�gY���y���j�?�.�<u��U��,�NjDI� [�*�ob@�kF�j_�L�oR��>��!-9�4u<��˩r�����K��a����Fk���v�����hw�F���[�#���K�cdo����\n%Bi��8��Ղ?��^)��|7"�X���8�Z���N[D�M��tG&[A&��8�̿P�rϹ"�A�SRR���T�_c�ؾ=
:����j�Tz�
�]�d2Y�!�.8x*�O'o�v`��x�*,�bA��քa�ڐep��;-��0L�w�eSD?�G�܉	�o4qo��ܵ���
t���Y�b�o8�:!�3�u�3�K,�[�M�-,S9��b2��U;���s�����^�!>�Skl�$ƪ��ح=����������5DN�����$qz�!�T`�,tҞ����������S��7,�Dp2~�=�� �X�C�;�����!��ݔ�ף �_4h���x�j�ld:�D��Ҕ����*E~x�|z�%�f�2���?R�~!ߒ�QYNQ�#�K��n[²	n��V�Y�&H�$O�<������'����Kır��o�Ji�N�u���VCZ�"Ag������8D��Q�S�Ғ�}C����m�e���L�<z��&��kq|�vʎoJV(nzZ�;���}�#��1Ćʰfƅ�sBH���؛هcڍڣ@暮�F��Μ����#��K�� �Z3��L�K����E;��8��l����	%?���B�)��tu�@��q�s7/:��~�k:�>��I�<MWf��Sq6��uE7���kԉ����ڵ���.L�y�7NP��	V��Y�pl�0f*���(D��k��R�J�a�CE���B�7
(��F���$.JĢF�-�:i�Ô�(�,j��?���e�m�]I�;+d[,�K{7��Ozx:P����-黛�h��N�#|u�}������g��~umײ��{���|���]���&&�+�����\��\�3�~&H[t��P�6>�+�!�o�ZO&��+��"�+����hJ�^3��5�*9r� 4�d�(����ԇ��e&zef�H^�*��/�nK2$�� '�kp�;#�>bߣl�]����� ����.�a����DM�пN�
 DFD��&%���Nr�:ޖ�5s����(�R�P0�;��o�-���X4)w1+Na�G�]dҷ�3�-Be�~��\���L)(���cw#�ʢ�s=-��7(�2���RP`��U�}]�~��zGq3\=NlP)uI|��>oD̓D��7\�ِ7���>�ꤎ��,0��^��_q������_l��k�pAt
"�^�#Q�Q
Q+�ܦ"<����͈Y���Tq�}���)'��z<�# �
A�%���Q�**���v�����3s�����_�}	+^�JN�P���Y��o��2Z���,\���,�\�^BNZԲ5gZ��ٗ�����댾��U�9ku�I��K�Dc�������5Eá���/����(�mj�����4d��q(4l��1�v^�f�?�,��ZF�BԤ�/�ΘRoH�7���&(����Ѧf��T;�q��ah���6%�m?���I�U�f?y��^ϟ���Oȿzc�[���E1C�_#o'��� �	ѸL�	��_bַy�Bnb�K������Kx�)Fɿ���Uzn�� s���=�u�7���g9s��������v���a('d�yp��9{ag����[���w��44~�4�ЦH^<�c�LY�w��شE}K>�+�9���E�g�Nzi�±���"�K���%C�u�]���~�c�L��H0I��hۣ�l�8U�u��jq�6b����`�:�=�_HM�D&����U��.� ���X�I��<@V����{�;��/,9�k@�O�#կ�7m7&�8%�
!�w�Ѯ�J�	̝y��y% [�s�s2��:7e�D}��g���Kg��M�o�դ<7�>P��! �r_�r��,��s�roN���	tU�Lh|�ٜ~�����7������,�8���f�1�>��[�A�o7�bPT�X��C����E'����d!r�>:Ѫ�U.F����Ib7 �p�/:��xN�b� ��C����v��7ZF�ATT�w��Q[kw=��m֢�iu<���;��yf�;�n��S�%s�E�S�b�㘍�����C��J���J%������8{��غ�нM���HWF�-&W;���	Ϛ�KA@����? R�D�<=b1oKs���w=��ŗn���q�7�!��|!ω�c�|
���N�:��$�t��l����)/]2���6���)j�m�Xn��lnWw5�omc�%�V�#��^��ޟ�I�ֳ�qH=3�5dt�6,��cM�TtQ@�o>�����s�t�Wr�S�R��!.�]�K�gcy��_H��1%������/��%1sm,����TiV�S�S?��
X��@ng$�7tho�,q�+kU-\R���=���z���amS~�4>�>���ri���=3���T��\u�i�N�Y�굷m��o�	[�*O,�������Ӷ�k�/`\�J��& ����<TCa�!�~��㴅Ȍ��Pl�E��-��9��Ȧ���ńR���U2�2HV_�F蝤�G�M�I_i��,x�{���7�u��0s�����x�n��0<{�yS�ܹy���#�����}n�Τ����B�T���@O}�%i�D�{� BQ3�	�wCT�lɧ諭�1�do�����0�<O??���O�S
vS�
�)J�Aa�`Hj`a��!�M�s"��4�jF����8�]Sd_H5f
�cݞ���}M�΢fK]��*��W���/}A��X�7F��p,�\$��J���5��f��P����X��t*2H�J�!qԹ�3V��(����U���l���"�ᴌ43SV)��q����PV��ݫ^FuhK�}�����FQڏ���&/�A��C�0�����R���� �is��z 3ӈ!��Tv���Q�+�yoƢ=�^�6�1��u^E���ͨh�y�ª:Y����E_hG$��..�q�lU�K ��>+�����pB��� ��ʀ{�H�󥉅3JhY!�/Ӏ�d0�7�S�����ȅ��·�� H�Lq���� /����+���j@��'��
��_Աq�'ԅ����.�a8�?џ����3V�ʙkY`�N�À��u�l�����V!�wI"�e��c 
xw�l�v�{n}�!a��Du�[� DۊG��� pݮY�'f�f�hK�=����넋�Qr!6���*�\/�bD���/�!�3	
7��x����!���f�%�۟V��D����**z'�T6�q� /h�=���.�*ߣ)9�:�u$_��jS܍��˶)�<%ÖA�2>�RC��)�����!�����]m�m�AE�ݥ0Y*iuf��.�l��4eW& H�e���1�mo g�&��"��wb�n�N�p�Q��p�z��CY��Z��wxuQ������~+4*'R��=�x�~ej:3%��0(H�m"#0BM����/��r����Z��:~��Y����oH8~�4�6�:���#���ک"�����y�i��dE�\��,C.�t����5�AJb5W�������<���X��x(-f�Hͳ~����`L,K}1��Sa��ɹ�)������uaӿ'�`�f�4{�̯�K��Y\M�;)��L��� �C�檴��Y{�������u?>x�cp�![h���)_�Ж��0��y]�G��`1E�~ٝ�/̽��H�7")9�U�P�#�p7�^.���^4��v��Ύ����V����� ?����~�c���	��V���}�����ID�_Pq-7��cZ�k���$��_r5��<(����n���U��j�bFQ���Y�Ƿ`�@�m�G��7�"�r�̷��Ǡ��	�[�/C�<�J"V٨���4����H�@�Qi�^&=�V&���E9���t���Q��������������yU�B"q���l��c�w7�CC�	��s�[���2��"
o����˿�L�6�<�<F�o̓�ZZ<h	e!j��5A�뗮yz>:b�R��L�ӕ�t�ۂ���K΋=Q�Y����A
^���?N���`��R\��Pc�~��e�����b���@/�����i-�3��/��j�I�z���lp���y��J��N�ܾ*0ZǢj:g~��`����e$a5�p_`�
���&R��M1{���&4�2���d��H�v�������2?Q�7T\����׫�9V�]��ь�$�!�4z�i\Z'nx���L1 0-����D(����|s��m��Μ�q5�~1�r{2H����`���d�m?�fR��˿����x��5)d6�t�TU���]8�o��N�����Κ�&�:5�4A��)z�5��_Ԩ=���`�t�u.�۹�q-����Х
t?�E�(ߣn:sd����O�.�AҪ�p?��g�2k5;��[�n�������Ɩ�M�����lb����>��$ B���y�A�e2j�O�������0{��K�	�wuC|�^&�����?�iKZ�#�Y�z���/ݨWRy��ݛ|@]Gy|�%N1��k}��-�)9��`���䭷�riv}�����@�g�0M�Q<sWO.�WAH'��*lpsv�����cX]��U!ܭ@j�b
�nf�bS�wi�L䇦೯�+�͐�خ������V��x�� T:�ڸ���@3�P-)ע�K�x���uS�Mž套ӿ�p�E��,[x�R����(��O6n-xю��2�1��ß�^���N/7$+:С>a4�Z;����BOE7��`�R�2=�(�3芼�S�W�m� M4�kQP�x�i��-�I�3اW�!�6<C�K�q':eM�J��'�mwԉms�m�*8��,�����~e���VP��4Nbf�@$�Yp���,�!$�� v���a�'�[b(D�H��R5A�j�.��
~K�*bw�ZJ^�O'��j�]���0#�!���F3&�I�"nz�^��n�|Im�7��x�ʔT�m`�LW����ACڴ�����B����]�Wa{��r�^F���ʗ�C$�g�c�m�T��7�+W���kc?h�B��'V"K�MR���FA��E��O*VW�R��1�;���<��� >N�a[F7�l!�B�\�Ҕ����	�#�/�#�8R�p9���9뱉1�P��w��-gL��>Ǩ#�C�5[�T-�z��Kk�'�V�9���an0i���n�E���$W�G��G��v�v��q����>�r�.b<�b������JNc�[�d�.c�}Z�*5�khkT�&�~��E4�z^k�_,6,+Ը��T~o{l�A8z���e�x:*Փ�?+~2��ą�yA���]q#λ_��7>#H��C��C#NkRX��7�,T�:��hi=��9:���O�	�+x�Y�8���&`��>�v�^�4�X�����l`�4N/
R��xj�^=aj�_=p����9�"_W��5uwڦ�i���D��A@��Ɉ}zS[g<zG�����P��{	��Hx��&�z��F�*��y~E�7^�%M3(���{�h�F��l����r�A8b8(2�L��U��:[f�"��a�uqm���C���VM�,���k\ۍ79���b���
�qJ jB
�%��OΐX�v�����)���Ȩ2,��,�$�s���1�f���Q������1%ߣy7�����H0{������zO��GD(m�H�z6P�[wBYn�Fd���Z5�ˡ�u�&2Ǻ#;�)�<���� �tM���,�'�(Q�����n�h�lcgY�e��T# �Q�� ��&�(�_P����$͙E��E�[�jv��}�q�ന��c�O�/���6���M���L�z�a7��M:�M�s9�'zZ�X�����܈����ɽLobn�!A����O�q���P2?F�TW���)�ea[Ä�<��\�l�T��}S-��Ɂ]��NhD�˾������Sp$����U��IF�P�Ib9%.	g�ڧo�l^�������?U�4��("/t�n���.�
)��]H���$8PY�꣪��2Z'�r"ŃwM�2'e3���1D���ҧ�����S�
{�N�b`��{ګ���ؽG��/\� R�n/7��q6���S�n��N���n�jϤ��ŃN�{PH��\���ِ��]0^�'tA0^8��#����]9A���j��]YHi�t��\t3w1/�ů�	�p��p9{� �S͖O��vS�Uv�1K���n4��iS[wk�X�z�`���6x%`��8d���qm ���B��:���5_�K��������.�dd�J�qt��s =��~ρB15g�\I�a���yħ}(�lhNY�Y��[�b!HC2��fM���$V6�h��u)5Բ��W����j���{ȋ9\����TDC��E¥�Iܛ�qT烙X�"��H��.���Ql��QiǛE󇴈��X��w�AW�E�l��a�ʪ{��P���$��9]�0-/���&f@3h�;�����X5r��Ae�l돤?:l�V&���ʏ���[����>r�����D�Ѡ�b��� \�gRث^�h]����{Syb��I��i�y5����#�= r{�ɑ
K����G�\�]iY��N˼lG��F�n"��"3�B���{��wbZ��.�bIB���+v�0+���);��_�S���H	��?�\hp�x��0`���e+DS��8cc�k)����ƍ+�ͻ���ag-|�r)q�4�l�M�o��6�Hf�X�� �)��?$&�rk9-�`�FtQUd�P�cn���y���%�����l���ع�� �VI=��O@np���t�Gj�$����)�HV3`�S�Q���"����"�����;tI�y�ć�袨��i�,��V���F �e.��ԉ2�<+��X��F��o�V�8�h�)n�R��Y��^�<�"ʶ-N}� S �V:��5�x a�5OF�H��_���%�C��зW+,��ڈP�PZ�$*����(�g��N�,�J�l�"I�6j��L0̤~�%��&����L3:U���u���d�ϗv��?qF�\�����|�]$lR�|?*�ہPﯚ�n���G�m��g����Ԇ�t�9��ʶ
�o��F@��o��R����0�V�ԣ�~ql����+՛���=���n��]��F�0�Dch�?(f�ӯ7�����2�$���Rj���9��+���qt��X����èN8���fɽ!�� ������g Bl�Hk9}m��%�#��C����$f��#�x��	�׫��=���\W���+�6�";#5w�f��{mx+/��<%|[��Os�<nJO�QJ
>�+@J,��6� T�Q<K���+�2+�:�g��������-(�ꌙ
��N��|&+Zr8�C�:eP���g0�de�]���O\]�l�.ޤʞg��x�Ǵ/��;$$~;�?�(vߋ���U0m4>�9\V
�ݫt�5��vـ���o����^�G�
�L��]$9�2�ޡ�~��������+>�[LQ��J�MR���<�K��������L�<�><2Pk:�}JÝ��?y{�j�dޒ*Lx��b0�(��v��(;,�S��x�nbK���D�][�Ŀ���ɿ�z�kc�3@���g3����	��{�`�Y���"�K'3�l�q�m��+ݚjk�a�\f.՟��3Y L���5+HS�U}9��io>��Ǳ�Nvy8DH���ʇ�La9�d����hbp i;P��W�j^�=D��a��eϴ�u�`��OV]N����1����Wa"=�5W��	�@ՠYH���!w�*Oo��b�r2-�c�l��}6VP��dq]�0t�p��i�Ź�8�&���j\�2N}��'�HW�ˎ��m�e��;�Y�.�c�q#"b&���Ov����_�Of�?�k�G��ۧ���TȀ�@�#�ev�Y2V_^|����Ǚ��lE����E�,�\m������/�!��^W�"��\��{�h�N�(�k������C1 	�3꾗����!u���I9����J(.1ג�.�\�/O:Z�
4�7��l�{/n��sA�0 �	-���dq���A���h���+P'v�mw��_��������Q���$��ׯ��+7-+̴	�>?�����zk��d!ݒí74��#�U�����Rq�q��֥=�] ��c�G��H~���"�����"v�k�e������7�F1}�C����L6Z�EDJ�_8�0W}o�H��y�z1vR#I�c�ʮs����5�աy�F�w�l�P']�9���U���s��e��pÏ�7A�=	ni4HT��+W;���� |[s'�}�g�yk69�#�~�nr�Ӵ��R~�)�P�#�j��rYj��ٸ��a�CY�ǵ��Te�G��tnz9���uV��#���PW��zF��{�)�L��b�s�+%T�^�)Bz�)�;��
j[��Q�lF�+Е�N*(�]�.�Ĭ�Ck��B2�{�#ՅA�lbA|9Kz��������y��.�w�i�>�?�a�.�f �yE����2�:�Ss�c[>�Pl���8��.���G� �a3��~p�_����"��� �g�;PD{���>�����F��w4C(�,Qx:���[&z�;ܽ����v�7�u���S
���������nN�}O��6��|)��A%e�kU-Pg�	T�����M� �����������4�
��e��6{%�7�Y8%�������G��ܾƤ7��;_� �!P�-׉���r<� �\�/v��8�y��^W�l杢�[B�^+�6K��AT������,�>��q|�X�8o���Pk����0o�3��{�%������X��c�?6�J>�)���b[��c���е۹Nc�#� �CJ����L���0�.L��:0��շnx͆ł�D9wʽ�"���	�����JYX��Yػ��AHe	@Ո�)C�]�n|f����Ȑ���F�Q���I��_��Z<���}1Ӆ�s��óJBp��[C�@Gՙ_#�"z�.�xvb/��ʣQM�d��L�s�r�n��`�����4��97(�| ����.�2/�UY����cv�H�9���tf��Tt�����:D��/�s<Q��6N"lgz�Ж�+�c��P4����F�z�p��(t�9/�v#Kv�{!�a8Þ����6-���SO��5l����^����#c��n�Ų��w�>X��R�J�6�= (�2��7�i���9�E ٕ�鶈u�u�*�����NDφ�IE�&�|����V#�
c3�=�c+"�r�&����,��F)L�]��^�OtWI�����8ZL��vr#~xS�J�#u>��X1�4.v׋�O~�q�H#��z�.�r�|������~��"������j�>����4�h�~s�b��Y�^=Id$�K�&k~�ı����	I�����_BGV�>�3�T;Ɔ!;��\LW�}���QtD��d���ܭo�M)ب��)����q��砀O�����c�ݓG� .Pr6��/�<�;^&O4f>�x�pH��Iq�@ 8�������V1�L8ޥ6hC�V.7�7�W���6�~v�y�&�V����xr�������k?��a.c�ۍL~V�����5�tF�q��`���xĈf��z�{����t}��7y����q�v�q]�i1{R&�)J��*���۬��91����m�N%t`b�']vL�/,����y��oW��x��;CѴ#\%Y#	grR-s�HEڳ�;P����Tb�F�$���)�~Ò��yd��k�(>��V:�^��O��ʙ!��0"r�[�X��K��=	��Ͱ��1L"���U���i[PM���\���ٮ�^�IK�E�~��X�r����\_�A[�3��]���-��Ϩ{�G��Q&��H�\�G�{�2 !)ˢVe��X��S�d��%�c)!��{_85�s����s^0m8Z���H�����oo&l�%R~��{6�[�>�,�����}V�?c����'(y8��LG'�"J�4[�7�Ү⹒�8&���LN��ݷ�̇F�e2^���ש�'n5�R���1GzU�o ��A�m@�׸�*2<8O�dly�N�X|d��\aɰC����h{�+�N�uI��
8#�	�����=j�B��O�ߎY\�7�5l�����X�z�Ow�|7UG�&�I]`I`Ω�CC�{k�XΏ�d�P!de��">Fd� ��ք��P� K������+�2������e�A�[�>p��&��� �+W���������2o�F1�)�����d�Џ��,��mGEɿkW;e�?lCy�*�S�IH�蕷sb�9��ޙA)�qT
B
M^��~$I>�:^\��n���i
я�= �?�*2T�亮�<g�Z4�s�cҿ�㈠^P�a6ܚfy�G�@��%���(�Pb\����ܵr&�mIk�G���5�/m)��Xx��'q��l$W���Qڂ�kԋnKV�$��VӮ��r����w>V�"	�Ȧw	x}t �p�����j�����>��1���t���Rkp�}�?+��T�S��_����I�����\=3���`��L����{�[�#�^Q��@����'d-��eӬ�~%�`&w�N ��s�VHln���3LO`�quS3����6P�
9�%!{�x3����i��Ж�gD�kP0�3F�M�6Ȯ�����Oq���m���e8����ĺ��O��9��,���׿�ه����wF&!%�\1�����P�=��2�/��O�����@/��O����jm�N�������j�4OF�G|?�`k�5ϐ+��o����^T\��,'4P1d�ƞ�6f;�늎c�b7H#8���A�g�=������ƌ`WI�H�s&�����QBߛ"�?B�xCYG$��:#�N�M���;��o�������.ND���	��Xڬu<өM�'�&�\ø/(6�=��1�~	"�N*Gb�a�gK�$Pq���O	�;���Lk�K
]z���.I-}3B�>D���jZ��d���DĮID�a*��iO��PW>'�ӓ�N�$qu�h���H�M}�7��RN6����i��?
p\�%�kA�~��'�Qt��D�4C2����f0k?g��� �]�3&�#��gtCm<�TM@P\�I�D��c`���*����%=)����?���E.3t�D�Ds����\��	�{M�_ǋHׯ�:N$�ut��r
Gc\��#���L9�+��{W���*\
_�*F
X�E~Q]��OX�TS�
��	����z�9��7��qw��>��@�x~���9���Q���UKh��^Ѵ�wO��o�L �%(�����Te��T�/��N;�t5�}��V����|������lK�U/x!10!���͆D��V���L����>����&���d+Ȃѕ�#��c�°C��M~&4���>�G�ۗ]�h�t�M��Ü1y��p�z;�i# C�0v��heVD��헹��uF��d�,}�����d�	���qm��u���Sa�̑�ڴ�ȷp��l ǎ�6?Lk��Y}M-����ӻ0����߾��ޭ���oR&�ߗ2��½zu8t/��T��m��+4������Q��Z��!s�D#ศy�%6'�x�$���{7����B���h�.�Ƹݫ_��Mk�DV�Nbր��{��Kg�Ù�S���{����/�9@,���r�ڼm���oZ�{���$4���=`�\t�>35=z�F�o������'���84`�ޱ�(��3���ʻ!Ks�C�f��ܪO�L�q��n���� ��~H6Ob��h��x�qb��-N�G����"�{	[�[�>����Y�I��w�����צ�*=�)������^t��A��)�n�jVe�+_��y�8PQJ���o��+M����t:x�:2�/�+}�Z���:�X���(��ᅋB:S��)NfҴ������*%������,�ϜX� ���&0SaÍ�Վ��K&��Y5Rn$�8S��e3�t����U��2��!�g^-qv=Y������ź�-��ȿ4����Y)P9�w�"��<�"N, D�{K������0�ن��IPj��O�8bS�Mv�^)n׎c*-���0���c�n�A�;<�d�'2� ��P�"��*�Y�К2��\7����D��|�Oč�f-]��y�S ,`&�ۻv�L���	D@� ���ْ����.����;yQh�QO$![a���D����n�� @���Z"VW��e��\"�-7��OΗ���yl�'�'��8,���q�jr�����l���ڭ�
R�z(���(."�e�ū^��/��������!�����߬����Z�'Hk�U9��+k��ۍ�H�U1L��>�~�ۤ�o/��2IuK����S�B�>I.ݝ30(�	�f41.���)hΈ~+lx�2�~���U4�t��(C/r�wS��ϖ�� ���ZJP؛�/�;�G�.�h��7<�L�,R��r/d�/$~�1��{qfe.WD:�S�Yת�K��F�L��H��ni�}�AB�\�Ċ���x����)�i����fq�J�)Bst����H��^)�D"�q4���h���H�CJ�M��5� ��KFW�ڙ�c#fX���1��J)��6��	�9h�S�]�"m0&U��� Uo�9�Y�íx�����e��~�?�������m�ķ��u6,
�l{1q�Z��[^#\�6�{�D�F���tͪ���]��5���abV��mCG�[�jGʻU�MC�B�r�_��\Y�N�2�?�k���9�?���s]|�~I�� O�$׳��P�R���\�vx~���4ۖ������� �0R�E���R 7^6Zw��yT�Ts#����Q����������j3�i�3���7Z�L<����Hk�&��e����1yo_PO�}��w�/?|(��B�C"u1ە��Z刾h�Gϵw�A�[) $"�m�U,�q��xj��Y[�4�_J���8��w�n�G�L(���i��$���� ����lcb%�r���<A�|ٿ5�߆��Lծ!6��+���cy5��/�>�~��$�$���c���Rp
d#���^Np�:64b:fw#m����Z/ݞ0�&wË�G���)D�r�Y���3�F����)��*�	XK��$)T_��~���l���
���$���P�0�U6�wn�9۳1fE�)g�4|Q�a[�
���
ΰ�m9���|�nmњٵ��ݦ����\�2W��^����#~�q����T6?�ZJ�����2x�A�9H��h��2�]�X_�B�?�T�%��{��dȀ�-�f�t vvyEd�Aᓉ܈L�l'���'Qǅ<m�s��
4�;�4��%W.\�t9:����ıZ9�Ԍ%���PF�O�`���"`2\�g��o7č�8"�e:\�}3Ω�B�-�'� #f���Ll���	�@����
�Q��@|�^��.�����g��pB��_���M�!�f�&�o�MT���ߔ͓|��{�׊k�G,�	i��UD�+��0W�ǁD��[S4<�ϏA��Z�D�rk��"�kY�1��[���s�ќp���5���I��K�K��n�~�۬����Tz��a�z��G]?��E��[7,ߕe|L�e���R�,zE���b/S� �/�|�G��{=�S?ZZ:�*�Ī��v?w� ��D�a]ӈt��^�Sx�Vy�z�d�{P�MC�$����(�H%�QN7��ӯ���<����S!*�{�ބR�a��T̐��4E�pǬ9�5��p�U���G梺��� �n ��|Ãts'H�<oiu7�TR����F[��v�u�f[����V�0����XI	���9�� E��LL��Y{dN�q^�<��d6��Wi��W���'ʾ�v�y��}gn��8%o {\��t,a�}����<9jg0�Ѧ��3fs�E��t,�E� �h8S����1T�0�Q�;�1F��,���g�v�� �� C,2%�@x��O(�p��p�5�||�����qg��a�d_7���u���н<�V�F��Ơˌ���u� �~X��G��ȓK����U��:h&�v;�nd�3��{D����gh���iߡ�T=1`�=���;��E�)X�kj0[@�;�.NF� �c�Ae��\0��?"	X��.g�F䴱���;��3xS'�p+R����gm�1U�Q@�5c��R���:�,��<Ckw�J�>C�����������Qb����?�?̞e�.��n��J�N��B� ��D�k��Ϲ�����k�Lti�*���_��{��y~!˳)��`ri��R��{�u	?a��2\�i�"�Ph��J4�������v�c�W�I��k�qp�*xH�u�߮�:�:�z�l]�Y%§@m$��C��!��j�d��"�;�	$s>�Z���J�F�5˄BxrDtj���d6vI��T���O�6\*�'#E-]i3z@D�,NQ?�}--�g�Ym��Ӫ���.n
��]����c�3�INL�}D5�2�ٖ�17+�],�n�h̽�����X:��vo�w�p�GK�غ���`r��>�(=7�����S��D�DxOW��q�^�|8���,V��B����=�iS	�o�P.�`�HH)��_�&���g<`�N�V��F+
_�S;H�� ϧm|P/A�r�?��G �pK�>�P�}�v�`�Gd����Ms$L{{���m9��-��J���L��.�QtD��t�>��F��.����50N�V��1�r����@5����<����ݩ�p�b=�Y.����[,��K ��N���I�X��U����mR��z�b�O$,��\�Pk��ƢW��I���v�d�%T�z+K��.�����k��4Uu鱅��u�faEve�:�|q�He%y3O�?��y��Ѧ4@'�����2�����f���vtt��
���G-�@���N60*�1�]�D|��>��bk�Ę��w�݆��$[���c��5���+�Ⱥ�
Ԇ{�!�Փ��o��Bn�?Ч�n���_Xe���t@(�?��߆�0c�6F��΋��7k�Gr���U#q޻Ѕzi���SQ[�v��=�2���r�]�l�n��/P��}���Ĩ�;���*X{���C"B�B��4���I�=��I|?w�5׭򋺖>�\�lC�f5�Yϗ����F��R��Ƥ/E����Se
�y��ID��'��,t��\>u�/'��K��
7mCi�����5��,��g$B�u�b�������sh�qޚ�����<@��卩�4r�%h9���䵒�Þ�x�~�@�ўo�ӎM ,t�Y�ļ��B��{��N�X���W��@����M�e�X'cB��I���+�F{�u'i�*��s60u����E���ŧ�g���Q$��b���x ���ӷx�ȓ:���_5�o�!���q�J�f��[��*w����5� N�I���FS�X�'�!�!���nc�r�k-j��Mo
��4>Qn�T���R�#V���������O����&��S�9� �����xEi_�S3����X�	�<M��Qj$��<w������h��o�������+l%�����S�s�8�v�F�E����^���Y� �6Jb��	ע��o+l�5��-�>�� ��< ��p�a�oJi��Me�f�q%"Q( �������z�6���p�I��	���T�1m{'���^�q�zx]�ޢ0�����������sTv)���ߔ��#�>��� ���@$bsQ!�=����X�2VͽEF9�H�[����>�F[.
�#�ۀo1�3U��!��[tR>n���KW��q�8��
�}]�ug��
'%9:L\P~��v���4�p���5����G%~��0�H���VA�sx��b�{�/�Y���-�.l�И��0�)G��UN��֒�N�1�'9�]�rۜ���}d�Tr�2��$5�ᅡ_�X"rTD_�����(�B����Nh?����m���'��)b���%��u%W�o��bȼ�Zu�i z�4�;�(0�ͩ�7���L6��)�G1����
k�/�ՠ��jY�ڮV���EM'S_e�K�4�}L-�oԪ����hM�M�JՎ&�u�q��{O�6g�[7�7�ˡj'�M$������x��>����+�s#�-پ�l���U�*������GYP�B\_|��8�>�~�ͩz��qK+3�৑����zH�F�b0���G� <I�.� &Q�'��R
c6�4�������nXx��7�K�j�DhO��S|�B̜�K���A��a���\*$��t@�m�M����ݢ�h�.��ē�,�V~��%kEN�'�������N�]�/<�x�}$�@����Ҭd��=v� !Ӄ���ོ\q��U���la5*G���b�uh��ʻ�|����B�*H�0�+�*j�X���b�O��"a�8lE���BC���A$�A�*����x&�,ݥ�ݵ#T ���	�'�e���̙)�^�,m'�>r��rXCM�.��+�Q��8�ul����?P�r�����q��|��fL�L��}��w�E��'�Zh� �tl0n����i�{�h�N����z���:}���lA�G�D�A�k��w˸�yPX蜑�A�	w�1���v�<.h+��_��'�2d�E�S��xS�oʃ�OrͲ�|�eT���%"����;�CD�ݳ���X�0w�b+L��M��:S� �p��ìCN��V�4���s�+�Z����%�Ț�񿏟nՇ�"�;�s㰁�I�c�g�Hd�`�K��b�P"���H���W�?�)�zGdn}������\ O��q ���h�T5�1�dɰ9tL�P���� T�7QD�P��Y�0�q1V*�Ҁ��������k��(��Um��������h)�z6��a�4f"VyߩԤOObܤr&#��?B&�Yj����6S*��)��ۙ���L�j��s~����Z�b�y�I>nMW�o����VlF֐u�yLu^l��QpR ۉw�o���:5��v��f͒�VP�و��i9��Y��%Ŕ���yN��n��3%�O\���u�?d�Z{AEp|Ly�!�jç]��昃��f��^ZDܠe���b&��;n4Ǩ��<v��/��~�g����ţ1k�E��\���8�^ʴw���""�}7�B����1>�����9��8���L6T�l�� �FePV���������Z�G�]�Ss`j:�UZ9wcRk�X���V�m���^��@���,,���͓�i=0MY���� ��:�!;�Y�,���_s���+v�vp@��cNݹe.��j�l���/�h�Vo�[�)^H����h�`��*�<I9?�kes��mǫṷ0Xy�:aw+�u*�%&���-;�]��8�(��NkW�E�c�e?_!W��i ���y��Et�X������5�F���jQ���/�� ��ڈN��p�f�`{�e	���#��#�`�� U~�3���K�4�]�/��$уC�͇������<�<����qVX�aJ���!MԆ��R����Y(�,Y���׊���;��c��L���~�#jҖ��,��_&���[r��;o+�d�\���-H�bÜC�O_ ���|d���K�CgcBkC��'�@�X���IK���z%h�`����gj����VϪ�i��as�i���ϸ0K���?S�G0��Ho����ڻT����7�D���+�<S�g���c^&�U��,�#v:����G !����n�Lvg�<�3|��Kh:�iYY'� �?�r�#�ك+F+J�����>�9�KB�	�����N�{mL��FAt9�l,�[���@���F��šƚ"� �t��|*�-�Z�	ꟻ��O��5�H��U���sSZl��q�g 3��KŁ~Gt�u�KKMd��Q,�[�ˉ�U�AV+sTS�UaPX�4H��R�n@�s��,�Bxkǈ!z�X8s�;;2�[�[��j��U��kk���}��Ot�{t]��%B���P&L�Q��ʡ^�q~��_B�T[(���� S�K�X�?�OL��t�A8��j�
���`욌�t�!ԧ����Z�p,ڹ�#}㴶��#p�F�������.�edLZ{�,�[gLo�I���C�@�9���F��ҧ�vpm}z>+�c4`,��d�I�������[��9�s
4}9�r٢g8o��z������F�����D�(ᗍ�����ػ9R��:�^�4�1�!�U���|�6&��Hd�Y��+M0�����N�=V�Ȓ1�Ѡ�%ױ�^߶検Z���?J�u[ C�������yQa��?����2x�t�!��K]��Xɏd�����B�rM��N������9A�c�b�[7��6�jAW����5ǟ�W�g�/���eG���E�d��"nv���֜2��RK���C�do9ӐN��WR�Z�#~���/%�z����w�C�	�lҔ
����R�ÏT\��������.?/������� B�/{"P�B��@���7�W3Q1��|�iP&�c�ZB�g�L��8�����!'����mG&)�vF-x�RmK�ΡUX����2������t�r<f��K� �l1�_[�K(ȁ}�'P\Cv�	 �&Q�Y�ڰ��ŶC �W�wnm�����[�T�(���~[<(��
�~��!_�
�߆&�>rkW�Y���k�Ҍ����D{�vp",��ܧ�c���@�pe�q}:�8�������)�W�+�F;��zz�	g�� �>�ҏ����<@mr��8:���
��
�тdzDb�M�9;�A�ÏNϡI^��O�c��ȼʮi7��Qմ^uP@{�<�X�%^ʧ٦
��l��l�TS�����k)2WR�2ύ+��(�{X�{��pE0�;�,��1k�B�U�(Au�^�~��K�iֆ1ܼ�qc�2pP�f6U� *-���=��փ
bB���!%Z��w6����KO�y�C��AE���^�L�(�kV!���e׋�*y9�l�����î[k��T��:0������y�,�^+��5>Q�a`tⅨG-�҅ �DN�B:+ٺve���jN�ư��ʮy�6w����s��n���՛��M�a�>Fؑ���w/Z�y1҆o� #����1�X<���Ǣ��Aݞ�\fm�³��o
�Si����;�j���Oj�q�WE9�r���R����V.�"O���[4>��3���;f�B��/gM��I?�����A!������ �(]L�sҦI8�h�4P��*%U�r>�M�B���^��l�+ ���aǷNB��"6p�L��die������t)2/0��/��yUR��	����pi�:�G��ψ�"ڿ�:������3cۅ�uh�R�M.ʵ){�D�r(~�Mh��.�}��.f����֝�ɾ��V���y�S�6|Jw�m�d�P�v*�Xz�x4��8���.������$Ob �W�v$��I`/�z��yӪ�t�lh'x�g���.���	y��`�,�ݙ٧W����Z��DC+,\C�4��u���k��\`��&�r�0�Ō��2^<��g��Jc���W:��e!�g	J<�&��=�]�o�J��0�+�=߯�����1��?=�>������?!��[�@l��蔗N�5�0=B��W켦�L׏���9ЏN��+�?@��bp�`v�
\Crf�<��Tg�lX�A3!>��F&W#����ʣ@MU:"1����(I�!�[슪�ϙ'�r��D�Z�p�p�Q�=� N����� r�?��B�Ƨq�]uO��'BM��N\��(�zQ�Nn����&�TPV!��G�ٴZ�WT�	G8��yX�
�^��?C���au��g .�&���c���mii$%�U�0���'b��mJb_*m����_�~{�����7��H���3%No��-�Q��	wC~E����j�(����?е�<���F�q�B��\�d���Ho�M)9��b�;�s�\�H�sL�D�%��E��>y@|�󀦈�k�G�ɩ�p�<u)5E**��l�2��N$��\S���++��J#u���{Z�݌dҁpCD��L�OC���.{:g�AUH^���F�Y�e���ܷ�c�[�Ţ��<"���Pmo޸����j��4�(��T��k#w���yMݨ$0%|Kd�{�rN�;YN[@"�4e��	۷���.���x�D��j<oHJ:����T"���"��-�y���5���F��f�K5h��A�(��D��_g	�P�0���E`�q�u�hp��?��4�V��*U��]��ჾ����Jؔ��T��NP��Dy�kr�:?On�R����.,B�vF ���6��a�������|sR���.��&빥�J`�.1���?.����?J��27ab>Y�<��?؛e�����*޲lv��,�1r�35�|�Rtn�ޚS���l�x����x�m�{����j�Г�y�pY=�98_�B{�5�8�hG�� ���� ���+{G@Ă	���U"`%�)��{�n��t�F�;��4���|?�<��,���s�F�l�h�?�<���#�HN��oz,I����LB��	k���j4���{qY��i89{�FG�WZ��◹C>�w�
,��:Æ��bmn��C*�Pd�] 	$�#�w`���L��/�eT'\C�Wx+ }}���G� �FoR^ȶ_4�M�ڦ��8��d�(j%+e�Z����e<�
1�G����lS��Q^��B;��;��y��+~��`Kqt���*��0�zP��5��������(ʠu����̳0���z^�F�{q�L��  *�GH;�q����H?�y�f��m˅Nz�	2�IKZ�&��wj ��#ŝ�/�M��N�h؁k/&3֋\�	B���Z��BS#mk���w��
l]5���.���� A��B�'�u#Q\f)'�,/��xGu��������^�ٌ��GZ[�Fl�6)Q�1�����%���q�m L�rb��亨{��:)����W�s��9�����H��h'Hpc^�xG��%�L?PD{(���9�Ak|��"�젛L_����1g&���
�l��3��)��������������������60�s���"��X;�n�i��s���,��%CkO�#ݜV��h�.�ØRRC���v��?�����<%���[q���JU���q��?xI�2|��/���i�/gW��7��/�3���-a_ë�z�EeK���;U?e�/�)��`k$����>��ꓟ+� �����k$G���.b�+��Lg�I���+����d��GΌg��jR��+�T��w2y��%���<~�:!=��@;`�{��U'3�f�ő�ޖ�I7�K�\~�ed�X��"s&�h���	�)��Ym�/y�~�PJ�z �Z���u;����k�$@�j[1@�2��u�t��oODt�0�$Z���˽�C��J�z�~����˝����3��q����ekӶ|a���|�s�]�����S�g�Q��l���)c������Y�9<S���e*E!*S�\�]��:,���+���}jI���X���)tn?=�4�)�(+��h%)�s8�u�vǷ�f���0�I�'�&�d�<��y|����A�D҈��_�N5�ʂ
f��WL/���=\���,1D���R�~��N�ZSB�z���.�sl�J�z�,vP'�� ST��R�L�<.p���l��u֌~��j�a�n
(ƙWRk+̲��|d����Ɉ�u	����\���i_�I��rã����-��$����@�+�!_bB�r��MA���/(�ո��~��g��ML�Z���ᙘL����r��(�Ţ���i`1,Rۜ(�^Nς}���Eg�����;^^z�ڭ��8�����}~m.Z��Y��T�O�ȼ�5��eK��T�:W�;Z�6R;�bvKk�d{�fд�+;l�=�v����5hA�z��0Ea����\����R�[�w)��&D�4!4#Ǣ\�4SO��P����b�(zs���Ej�3Ѣq��;���E&QC4���l���h*��ao3:����]f ��z`ku1���u5KJ# Y*.����>� �egC�'�pb�:�A��������C�M1jI�k��w�R�����29�U���!�vK���H�����2���OP���H��2_l��>)�V&�h�?��2��]}9��*�7�*��
ar�f^�2G����6��A�wM.bo�V<h;�h|���)�@��ph������]-+��~!@���<��W{�s�@�����:	���������CXb:̃�!3�̈́��~�M�(���WÏ�g�#����!Z��V{��nx蜇��)��PM@~l>�r	�����JX�]��_h�co���<긼?n��v�F�
�{�S޺@����E����E4j| J}
Ȥ��mS���Tf�m��G�����M������S����AEt��ȌۢUWB�A9�ڨi�.<��'��+�!�B�-�;�����5�*�X������#��!�N��m�X<D��o���	��ٍĠ�:�غ�>M5!��*o6��m���>�����Yes�����h�vs�'Ue�~{��e{6#e;wa�vQ���ou�����c�����B���^	���]�`�b#����.��S�3� O�T���D7T�8�c�}�����h�,�E����8�Z$�ߦ"��,'09�p���y��kc�S�����;$ϒ�G[������{l&k�8\P3�6�*"V�'nlh�r&��L��A~%J���e��uVl'�H�v�Qԅ��R/ո�3�%61��'��(��=���lC��#�c_��#D����#��ٕ��_<���u$���姦��W܈�ǅ�B1�� q&�W�`��`�{��19�r�z@;��<e�/�[���cMR=,ѳ��y�ߑ󓵳Oa@S�Jy(kK��=^{��P�s^qy�޲u=F�~ř{�nw�Zbc�n� ��W�a�����nc�վz�~tH�<CU��ή}S�6�.�x:0��L���6��5"o������U��k�H��ʻA�.!��0Qp>��X��O��E�]����z
���YE�KV@�ڞ��%FϺ�6D�[�&y^����.!H�6����X�d�p\�C��`��Lt|f(������i�T���nc�&�P)���������~��� N8�uY��_J� y(�H���$#p�V�����"ӌ�+���g�åG�.`�#��!�|���B�!W;�������|6���qI(�8C8bND����w!zI�3V�F�0T78�L�%��'X���MzXJ�����u_s�eK⟰��[�_j\�y��Rk��mH�2�!�,8^zp6�����옠$*|����wJ��ϣ$[}s�Q'�Kiߌ�U���~�z
}㖔�C�P�����8N#���N}��4�܈@�*�6�Իu�M��	B�� ;qد��9�F>}n����3���ӣ���?��Q��Q�?�, � �K}X���w�I�I9I�'��%L�$-<S��OP�`�-�ym��;2q[�F�F�)��+�O|S�v�<�B���i�g�4! s�󯖭r�s*䈿�N94f �w�u���a�rg	�#�;����@P��s��0�eJ]cֹP�&����ŶV��zZ�Q�<eQ��L����0�Vl������\`��1��)��������%8��j��#����H��#b6�s	��T��Z��pǢXNn�&7\g�4�O^q)�'�?��&���#t��"�<A�A��5���ͬ&�AY+9Y����]h��wFv^�D�%2�3Mڍ
�g��ܬ:�8�u�HV�!,�VS��&h��B���(��b �+'�w���<�։�;����x�d����7�F2b*14voMd��*:?il�Qf�Gг��Ky(�PX=�T�L�M��y"�_~��x۬Hh��	G]���8�5�ߦ>�K�����H҉���.�j�+GÏ>�ɘ&�S%� �c�>�ݯu2��	�+�k<���P� �Jн��Z	�J������
����:,/A��?���!��f�Ƴ=�cx���2�[�iYg�Cˌݠ�o�4��>�b��������5=5[ڔ4<l�V�[���Nro9���.���ֈ��+�D�
���"[�(B1���! S�8�(��H��B# �:�������02���/�X;��qit�a1z&F�؟py��cCڷ�Μ�]��Cz�&e�,�7i�W�ܴ�q���JK	��(�w���lɕ��'�#�u�15���X݆j#�`��Q�z�YF��&U�GҴOL��������!��t,�T'���\=[��ь�wї�s��m�\���`����36�(�E��]@oA�oc'i�服�_$_y+g4�	��:i��kx���F��0^��F/�f�@��*�j�"03p����=
O�9�4���|�nJ����U��AW~��&6Hgs%�}!�"u���"t��1�--�-�S@��_F\ST.u.��l�i���8�2i�������"��J9�n�I���7
n�6�=nc"S�>��bg��&�F����Py�X6#���`G�03�"�	�&��Q�Qg268~���ʛ�!��<���M
�hA0��?F��D(�-��'D�(���'v�y<2ټ*���n%IRO'��*X:����!9ܩ�D<�?�a,�fՂ �M�0���i�S�w�����d�A޻���q�H��t�B���Y��d��Ή�h�%g��6�ܹ+ǰ�YQ�B+�͖W` Wp*��<"���_�������Ů+�s1��x���Zت��e�pZQ��H>o�z	L(��o���*lpE���"[��|t���B5��#�O�^��fғ�!�alp��Z@E�,��G�=E��e���-$�K�W�%$`�R'��W�Whҙ>c�k/�Ԩ�U�"����Q�$�i���w]',��XJ��+F$����a��!#��-U���O�*{=w�g��<\��mͱbiZ����9_�H#�n�]�e1=�M�BBt�-I#������,,>�om 0�o֠����e����X8h�Yy��'�O��Uֱj7z�m��a�qm"��>����y��D�lC	�Z��#����z[�1�`̐�?��)������I���вV�s�Jp� �<?)������Gs��]u1��p�}*�3,(��I�Q�� ��/|���Vm-�"��Ƿ{���KC��Ge�	��k=��+ ǅ��=�ԍ(�imЪ8���.YiW�X}e��,]o��V��LlU�$�-�k�����9�R{�����9��D;�k���q-��DSp`�՗�5��*�e����i�j1wn����w�?&r�Fj�{?3��E%�p���w����4�3&�{���k��	�����=u��
�7&䖇jH�-� y(J�~�ҷ��jM��7��Y�屙;�&�M�V����	��-�Է���mdU��������!]g
4�ؓ��7�8N��t���E�Ϊ:C->�9���>7:�M�#O%ThqZ1��&�!9�ϒ����<��x��\8�R��&�o5�ƚ�ɩ�
*GL�  �+�5���}2�Ĝ�8lU��q��М���/(q�ꆥ��c��ū�M���>sٰj,q����^��fN1}� �5�Y�����ߵ�[���Gp��v���h�]��a()��4�Vj4}�b�F��! �j�FeS �[+L̐�9"22��̒��$��]sֲ,�
�Ƶ�Ƌ�Wt����2B��X�Q�ޝ�{��6OGD����E�ާ�����W?�KE��np{�g/U������Ԣ���]b�͟IgIi��(�uP�ͥ^D�r���f��#.ҧ�|�<z
�ueM�s������|�=e&e��A�13�3���&�~�FK�MB$�1�EBM.q'|������r�B���F������(T����'�	o쇩S��&�0�ؠ�hOZ�lZ ,��J$4`%�e<9y���䱎N��B�ai���;Q�޸��k�ܺ_^�J��߄���K�쯯@�$�Q��5�4 H`�	fM�A���:/�KƉ���Joh,���1�����
cB\�9�>�OE�ZRX��Ls�����	���dsV'`�״�t��ާ�]�ИdB�z������b� ���49H�A���)��rie��m�}c/"ʺҵ�+����)bx�@]e�,��Pp�x�h�J?�^j� J[o�y���@����J�^���j��Fo���:0d�G��$�l��"�����
�Iebe�OC��#��y�?�珳�8a����"�	8l��L>2Q�D�h���Cu�Eat&���x��c���x���9����*%���1�`ⶇ/�V|F������5��@Z�/tl
�&�p��/;8_[��P=��Α!�c��Ơ��|>��v6�s�����L��n8�IZ�v���.��n�J�j��0z���ҵ��л���ZUG}Ӑ������#�ϖ�Q���F��i�@��O�8:�E�3xE�Z�:�B��I�6�ޟ[o�˵i�Yx�iEb�(j���-)	f*���P|��͜f	SL���P��D
h�N�$�����g�� =go����>���\��2:1dN�*����<��a��A�h-Y�n�h�u
+A����3O:��Nl�0[r��o����8�8<�2�L�B��Z�q��Q�`���R����!7�EՎS(A:#a��!Ϛr5���ǁ����.������&
F�f�&o��b5�󦞭^"��8h@I�?
��&��Q�6l_#l��3�!���2�a�S���%�kn��p��5�[1qh���$�!�Gn_��K�K�n�Z�wä@��]� ��./�,�1�6���;�=z;����X[w����.#O�8Y9�W/n�/��nI��E�W���h'4'��̠�^�*�q����3�M��jF���P��8�N��R��`L�`E��(��fl�7��`�l��wH���9qg�jv����M f��z'BQÔ�\���gG4�ϖg�l8�I4�I,�BA�G{��L4�SO�DT��O���Y�9� ��@R�sH10\5.౸���w��"R�K����+���l�U��I��Ac]tanDWe!��ޫ�=�l�{�p���"��m|5�������5���%��u/��\�'��?S ���ܽ1&/g���x������ֻo���Xg1 �j�4qw����xɐ�r`ȡ�T:M �=��*"��	8k�ހ�kmR�?�eub�(���-�F��3�Ay��R�X��7⌦�K}�<�^͞��3EI,��B��wg�v	$�u��O�8J�!;�A�L��'1T[�����g�pg�����#W��s��f��p�򉱤G|�@���0��n�2�7k�:R�G��-���>6�o�n��2�T�	@���C%� Q�F�Ƶp�`������)4h[.`������*�@�g�1�b�Вյ^���o��2�'7��ܮ��<�@�;v}!�#�R�>qǅ��-R%�4�݌:`ٴ��}����d(�Q_w.~V>u����!�J(���aQ�I��$^�7T�+�C��?��JX�;��Y;A����m���	}��U�n,����=���B�`@c��k�;�<ö�wd�с�c�����Z+&y"r$u�!_�lae�I�QN~ċݍ0��`$h���G��J�n�$�
΢�[��l/�~��:�����E�u�`4<r�!l�Jۈ�c���,���˒ܰ52��|V�Y�df�󼌱�H�;B7Xa'B!�(�B�ұ�"����4}�\�AB�.R�iI�G�洍
��(��-�����`A�7i�.���~�4�3�2���h��Q���G� �����rJ-V�B8�mC#߅.���נY<-S���X���)O���<2�/ז��B��V�����A7F���Ҥ�]q��Y�G�¯��=\�^�k�x�>��X=Fd���W�{�HM�E�!n��#�-��?����	�-���䤽�?`�#�8��vzH7n�O1c;�����`XJ뀸��XFP*+�7΍��>���&wP�P?��<�i��kn�� _,�$o�L�$#�a�b��`!�����]]<0_�-+�G0�	C�76-m{iV�z�F��s�q� S@��N$*Z�v�e�����D�X�����#TF��,v���҅=փE�jޏ���"^��׺� �cj��|��e��`�J��rU��{Α_\f¢�G-F��W$�M�✐ N��!s��[+��/�.�p<�d��|�Pc�Z�p�K��T�u<#��y��m��B����2��T�Ԏ]�2	0{��M��
�ou�M��s��M�aa��v�>�k꽸2�e���Q->��\tC�*r���FLi���:;��P%Ap-6�i��Do�aӜ�ҭ�-��V+�Fy�
�[CX���k��o1Ї����4n-#��&��Ԣ�9¾s�8Հ����7���eYVP��	�L��arr�����&����Pv�"N�h��6D�$�㬊	L�[��r��W�d�$_�L�&�P��+�A}x��k<��m��}q%h�
��2="��u������@Għ��/�?S͙�5Ye׷9%LƂ�@3�N3AHo������j5Ѯ��usnڥhs*�)y��K�4�ڐn,�]#t|\J3��H �&�-�j��u::��ϩSɹ�1��'Xؠos</�ta`���Ƶ���C��6|t��|���W˂.p)3^R�^r8���G�д,P��"s��Ka��ҢҴ~��$��]�	�n�PH�����B靛�ǵ���F�`�/(*���gi��1��pT��ZO����t�J���x�=�ߚS��A<9�ot��h��(�l��P����tȒ�5KO-Y%�!3.�*�����x]��~��a���1��đ�f� ��>D��@���V� -Uq!�<PҤ�As�r*����Μ<��$���rݔ��o���/jA�^ꀉ���ñ����y�xoX��h\�G�C���8��_^N�����F��>\�v���,�ē�V��]֛�E��:%nE��iĤ��-�`J�0넟ǈ]�㜒.���eŇ����k��.^���:}���6�0O>/ʁ��5a�b�i@��b��@;r$�e/Z�继q�j��_��$�IE�C~-2����"�N��`�+��t���bƛ�H)���p]��e�J�y���6�t)�P��E��_���+��E�'�lT��oR)р�lץm,/?U+��1�Iym1:�Q��� ��uhkx�����
�1��!���jt��.�,s��Qkh��V�@Ҩ̤p�9
R�X/�Z�Kt1)/�Vjih~V��&`^U$�&��Q�躃��H�oG�ۙ�� ��QJ���"��2:"7 �}����%I���䤋�����w�Z���!
z,�����^:�fP?��vs|MG5��oVQ��?_q���=�m���dؼP�7� �j���|U�G����T[��5�,�y�[�؟�V۵�>�q�:({y%�bA[r�?M�l��uKf�����c�_ӡ)
R!;v~�>�O-*�x�o�ߩᏬ?3FN�Y�ŗp�Sq:a,�Q�Y�������@�/ϓh��:41ǌzI��ع��.� ��>�At2���9C���F����	�$�U/ڔ�L!�8E߭�
į@ַ]V�KJ^Sl�RO�0��H��Q)�������m4As'֍s2���_�C��x.���2O,��?,e���[Sן��x�1���H՟��f(�P%�?xv��d��:���*����ſg) C�P^$��poha�>z�"R���=��ʗ��c+�SV�N�=�({��"V�2��fc�ynV̅���,�/��] ^D<:��JTq�<l�i�r�n�h�u���b��2C�9�~䯀�%��24�`�28��ͧ���Hl��k�0�y"���=��	�������`F�ymk�A��^u�*fu ���8:���@���{ HV�8�u���6jL���'+���v�����ZU�;׀�\��܍f]�Wh�A���I̷��w�����g �4��c�w�!�vo,f4jZ��XW�#��0�`��ciM��`�����Ļ\Q��T���#�G_�J��~��챚wu��,C�[��D���B0�Dv.��p��rU����޴�0#.�)H�H&E�=��xZ�j�Gj��u��}ɲ�v]�Dj��x`N9�����ɣD��#܊yk�$1p��D��[�\�V��/j� �Fj
}!�s���l��ցٚD~m`ۂ@x����=�++jRs@�WCZ Rf^� ��Nݍ{�3��QΈ�D�9���ʝ��JzPճZ�'�+�!��`��]o�}Vٓ��L����L?�v5�����m��ڍ`w���gO�C�ˉ�L��g�6jW�a��o*ɾ@L�{F�ha�D�>$9	%
��T��d޼�	��ʉ�+��Ջ���.C�ܽa?X>=1E�#����p3=xlB]�W��Aڋ�Z�����A�ᚖ������J6�4��97?W9dJ����h���� ���a�t,�����F;�ˆ8�<�5�\l��u���x�u�i���&�	`IS���=��q��퉏]�I+|�SH�� ��B����_4{�Kz�%�t�'�V�	�@����p�n�Ih��g,�����1�������qoQ��';I�e$��?Ј�O�g��MCg-!o�HPM�V�e.���'��;���~�3���,����-�}$��"��z�h�i�:�曟��V�:�^��0.�9G��\#�9L���@�5��0S7,$2�d�
r�B\?އ���8 �T��-��.��x,Kov���+�"ـV2��9�mٛ�M���F�6��+�7�����e��C�(��,|�>ݸ�Fhɲ�/�wϒW���2ϡ��%O��'d��P�����ڙ�sT'��DT��m8ϿϚ�'��AS�1�)�$�=��� ���ǲm(΁j`Ot��{�}\�@i� ��o��
&$0�C`6��S@�����o�	u�C��K}��AC�4���&k�C�=���ńx�����0���A����,��Z���7��͇W�)�Gq٣�;,	9�����}���/U�O�ڿ_:��!FVyB�w,�֯�e�	_�Zz�;�xz��������iqo�'��p����M�w\�O=�Y'傥&�����m�[׳�VR�|�}���?&�v	d,^R 3�<fy��=vY��~��?���Ob/�cL�L��082sk�ϙ����Y�s����:��h^8et��3�H8�"<��N��ɤ����6	O��C�v��,��~T 4R��5�F��lɗ�&|�ޓ�`����dp;`�6,��p���'I��eK�s���X%���ǋ��>����4�)���L��{�kH�~t-.M�NL�� #���t��z-p���M�@ ����'�*$�AQ���tJ�Ű'yw�
�z��"�)���#�>N�� �8����a!�㉒�Ω�����f��685m�!8Μv�w��w�Do"��Jl51u���ڃ��f��O�2_(�r��x���HcЬ���D$�ȴ����z�M�:�:����KQ����IMe�i���h����s,M%����8
���4~;hf��84�e}n&�����F��N ��)G�vf|��dFd�qz�������A%��e	�0���\�%#���ԗkY�/�n<�B��	�a��O�xX�I�#fFН�2ٺ���W���8Bl/7L�\�0��hrt�ȿo���'}00UO�T�~:dR�26�q��92�4s�	���B�E0N�.T+nP��>�������
Ix��Pr�/���
X�G�-�NH3ಀ�}�z���P��pQ9������U?|��"��%%��
��]��s�QM7��bg��S����t�>���z�����V/vx���Շ��+[<�y�3
/����x�kk�>?�T�G��k�[M�.���El�aP8*�PP�O2'�2�C��Ņ�'sg�}�m�SJ�l�.�g���>?�������%t�'_�:ج7��`�૫s�&\���ǁb��Y��w�TX�De<��	���}%� �/���$�.��E�QS����P���Y�"������>�Ie5���0�2h���,�A�O��gv�(�H�]��G��,�Q3���8�w�!=�Ko�t���F�fgU���n�����ѐ{�� ޽�:1sh�*e]�Ƨ#���dRppSc��]��"k�i
 }�Q���g-Bj)yP�u�2�ѷ�* =7ۨX5�Y�<�GaN��dH�3Id"R3��rq�;! '~��!�Tf�:����"��]�ڂLF!O:9ԫ<�xƊ)�C����em�E�M���gC���_L��4�bނxC���F�I9��}xz�3&����ɏ]"qh�FZl��j�q��%4�b�G�d�e�b�K��;mju��W�L��6^�����WȪ>���[a�Q�3��j!�r�Yp�_�1Ӷ.��ux`J��S���]d��*&T��"�&��>mBf��1�;�R	�Ak����
m,�r%,���i"28~|�㚰��@T�߃���f?\lT����P��q\���MM9��&�@��5�caZ�K=ީ滖@�x�	�O��"�-C�ѡk�2�FnL�~Z�%���ǲ�M��K*�ȵێ��bx8���*}���?�l$����j޺&6�V��)k�Ly�I ߒQ3%_4��]�S�2�u�k�?&��"��Pn�ך��`j�80��1"¿ꏧ���L]f]�Ml	�j����*f|x]ʞ��^��ۊ்%�&���=���{Ƙ��1Q�f���ˆ��}�kzW�ȯ۴�t�@uGz�Z�L��Xq�]l���A�����{ �3	Z֝�%����2��
��skBk7�~o�*�X���!��6�I�A��G&yl1��u&̈́V���;N�?i$KNB��j�¿Z����aA��;VY�Q���jQ�ցA�I攤q���?����i�~b��hP�?�ᤍ��e���ާ�3���+aj�WPC�B?	I}��o��+��G"j6t�Յ�O��'E�~Eb��	�k��S����I�y�i.����g�TO��,"��S��eT,M�t�Z����Xb��c"�@ݺ���]�Ru)�������f.X>�V��i���6�mO�{F�b�f�Ӓf[�d��p v���X!�J�����+�Z�̪A�y��j\���w�I[з>\�Ck>"3�qt�6͛���f���	�7f.S
/�����%'h�p�3�l�$��`^d��=F(�9�'�W�d�����{��V��n\�n��`n�4]>^P�n<?9��߯��m�q���0]����pO9K\�(��,g�7[%�r\������߇���t�����ϱ(�oa�bgU����:�b�%��48�>����)r��ͦ�COq�߹��1>�h���u�k���jY�������w�i�ؑa�郡!�X9e�<���h<�Hg1�����t3	�A����i-C>���	�$IFapN	"��&vd
s����t��6&�͖�`�?��2G�4"�v��Wra�
�(�ۜ#_�3�矬p�^:���
��fz�����%�#�镘f�QG��yO�[�Ѭ=v��X�S��qmܕ�폞�E��$Ŕ�'�Ts��89�Q�
�I�7_sO��lþ��'��������Ta���ʣ��
�I<����N'ƍD1D�W=�Y�佯���ۉ'm"Oj0㚩�B������Ҁ�Q���F-nZ�e����Z��Tq:c�b�g4��)��gQ�V��1V��)䉪�M���s)FODj,�'�@��N`�E���m>����}���D�r�iĦ�5,b]�l`^�X�VOT��be��?璙	�l%���+]:5�rT*�O�m���$��m�9z�[׿���>��)2�R-�:�1��GS|��"�ن�Q��j���s��q�	^	�����/h�Lh:*�I`�q� @öd� ���9�@,4���ʏ��H�����0�n��!d��Y�X�ly��աx�u#f� ��M.�FaM��v�?�C�`Ꝑ����%�%��
�ԋ:��EM�g�>��A�}i���'><o�+tO��ݵ��Y�ɒ�����4�	�gO�Hgċ��A�w�ǖ���l��$x&�|�R��EB�UJ
}��ɱȤ� �<Vod�F=nlBf1�A�����/����?���X�CI�=[�r*�ޠ���`C�����yg%tP賘#�Ⱦ����n�X�{e�;q��|�Jn�K�#�,I<��T�0�{���\?���T��Z�8�����Ic�b�SK��w�
N��j��?*���4R�����o$Y	������,����B��������v�"*�Q?��������)uvk�E�����D�Z�-W+o 燿��=����j%-^���Y����^Qڍ�M�5nZG��W7�~�"�JD%�����[P"]ZQ�^ONXuŃlT~�4�*F8�?X�:;�Qr����G"|�9��,䛅á�i!�+�u)jD�f��.��l-%a�i��YT�p�u-.��Fa`4ۭ��~��~NT4�M��h�y?�Qc�0$��T9t,�;�������E�D�Q����ͷ�����y�?R��ϥN�_���c$��r�p�l�f��7p���Z�_e�mV�A�(>�M򎐿�F�q�'���ľʱ�[Xk�*�[�;��!�ͻw�U���X��w�[�'���*R׌���l�s�1���/�@2߭�7ϑ0���#2:U�'7��;	����5���%�O9����Ȁ���l�ƴDl�f�Z��뿻�"J3B>��	��A����~'
�0`�?�m�N��@�f�r��w���� #/Q�Ҝ���,�հ>�OD���h�E5߬`!i��8��]ͼ\`����=�f�>Z&_@��BB�p���/!��r�y����S>
o�����2S^d0Zۤ����DKl5��GX��i�on�hu ��
fq��2è:)K��x��eֻ)"a8�w�8:���&Z����a�^�~3 ���ɫ7d!��a3QO�f�"FG}AŅoK#��C��Q�.F�Y-'�P��i�c���0����rL��������i�LA ��=���t;@W����K�!,P�S������X����5��dIZ�_���T[��:��k�?hN�����B{���HٚPo���;x��9�{�Y�;�4�;���~�E{�9�S�k�~�v�`@���+c����ә�:"w�g;�D����\�W�픣k��Oݑ�㮝�(���谦���s������5��mQQT����ق��>u@�Tz#�X��yb�d�����|v��|A��snMyn�¨ˬ��]8w"d ��
�"��9��~�g�N;�Kq{����?��TE����S�K���;h���۬6�f!���'c�&͑������R��jqg{�8��7�o��v����d/>�d���_%�M'�4k�?7�!KDNP2�I����*�y��4���8��EO�>j�.�r��i��+�5���c��@8�Q�ѕy���]���I���>� ������}TY`�j�Z�������F�&��6+�9��.�$�S�e�i���|�� !#2��ua&�6S.���rO�Z�p��Jk���nL�����K�R�n 5=�e�re=A�w��Ŀ��W��^�K���%ƿ�uX��Ƅ�)F�t�p� z���x\VAD�~�%R��f�p7��Dž���TC��|pؖ��[����K��i�o�&�*��i�G	��u�
�A��77�Y;�פ�cg�9�7��)�)j��z���B�W!ek����$'�q�H�@7�m�ʤ����#�!�^�7Y��@�S���Z�Qv0�]N���f���G�Z��⨫ u�ڀ�ji\�b���W�VΘ�ܢ�_af�9p�^v��K��ӊ���)r�R�^![,�h��%P��qff+�>JW��կ���S��IHH���w�(E�_2�Օe��o�4�]��B'��ѝ�ڤc��"R4�)9��<-@�&i�A4��~y(�Ӣg""Ul%�A�����Qt>kY�{+��{��ByS��A6�|wO&��>z��'v��lDs�>��O !�sG�ǧ�����Jx�]?�; �L��� N��5���$�ƺ;N��6ݨe��;���H^���?k�zݰ�В����&8I_�����s�\�-�.>��A�⺟EF��{r���y���9e9���F�&��F�'7�w��Ar1dlGi��_��;Q�n������{��|q`_<9�~QK�Ph{]���I?>�2>kt�����U�&	�7���4?X��#6o�HLlKV�[��M��.vH#D�u�)�X��Ev��D�!�хa)'��K�R�����J�Pg�zm�
݃��8�紨uE�����x�ݢ�ʺDr]u����[�jM�x�ڌ)�)�μ�ٖ��F`5�O}�.n&�8c8�T^�:֎c�ZG����.�P�ESh��G5 �a�֜�l��`����LeU6y�8~R��+v���0����h���VP�ƌ�׉�v8=�N^�d~_�VܫFg?����h��y�q�j�n�S���^1I��異���<��+�I/�گ���.j�N�y ��M�"���f�}i�kj�m`ћ��S�H�d�K�c?3��X^��t���
ew���U�w�.��q'����>�����a��?�^�����ի�1���zCS
���J�agq�`EO��ő\rnK�:3�?�
=Ԭ<�e��\߅�;�+F���)f&�]Q�#^f��Ү�J	ߠ
!̄e�wwE�DN
_ؑ��[�mqO5��Dՠ�႔i��1�L����s��܏Ս4�S���H���~03�%���|'�Ӣk41��4�D��٥ԥ?�#���hTy;-'�7��p�N����:U��"��kO≹o��sG��s������(/{��*���b����"�PBx��5l��S"1��2���4Q�H����P��&�n�P�k�w��P�}*e��c��gW~v��FA��W�K�2\"w��J��8���F�Wǎ�0���j��� +ټ<(t��4�M�d �kF�,Sˮ
����o���"��<&�D�`/
�CHP��Y&�*��|Ʊ��UE��a� !��љ+$8:�y������^`�`8�ݴ:���FW����M ,��%�V�.�����Yp�a:A!�6"��̰'��:��a��9bV�EnA5����+��)��w�Y^���z����
��^I�\��]��7���ۿ��x[�ӡt;e���_F
�:���U�e����%��_~���wԂN���z&��C�_/<��S;7�Oą��~/�v�<Gf��˃O����]�X���f�f��t���>z�L9-�g����Ơ.=����ݶ�B��Rk�+��}5R�~�����Ow��&1z�0�=�S��_	��$���C�sA�����K1�
�!�Ì��J��4�k.u
#��j`y�r~�0'���}���L�
�"���/�ԚS����pS̏k��p���,dt@ϩ|t�N�i"�����^C(��ܜ/%n�i�3osӓ= 0=Z��a�~�#QR`�C����&[;�No$�����wӘZ5�5�0N,[����d�I0C�?�k5n _)�pu�X�_�T��xc$�C�;�8u�0�w �4T��J�Y/E*Q�w�Z���0����iy��S�x�
�WtH��O�+R�īu#	`��3�K�(�`����
����* ��s+\�u#�[�1�^p<�g���('���D�tL�p��(P��1�� Tv��3�ɇ���\m��3x$�
#������8��p�@����kn3J ��M�W>"�|��H3�$� ��X��ve��O��:ǝ��R��,�z�غE`�(��������b"�9���%���4C��4�V|�|�P��#lO�UDAȧ6*��<��$3vI�A1��N�\ìM�2�2��������m��)v��>/�O�1�����]8�"�\�]��|�xsW
&D2|.�S���?_`^z�0j��S�0\,�p��N�L�3j[e��*GW�А!�����*�E����"�����[�9Nv`�R?��x��<%����,u��aUlC�ݴ�^��Ft�G��ZPS�_�H�|���>�q��섓P
K���xu�Oz��s[_��.�n/� q�����чo�Y�&.�=����+oL��q-9�����(qK�V⢋����\5nP/�k�@]�u���j�)�]����N �����:�Yg�N9ob��v���o�:�2���M�B`4�&!E�ň�x�Υ���NI���>V����
^��@�'J.��XQ%W�~�lj$��a�+���w�
�o��p҂5e�U�G"% �`���U��9�Bʢ�N���Yݧh����>3%N��5;�1竛�Γ@!YN��5��$��"5��+�UN?���0̚rs�SA��d�bi@�:s+Ȧ�(�f����elT�;��u����.�����I��'ҿh2l�w�����蝱,�2�Lw9��Af6y�gj��s�.l��(�p"X��/��l�h�EQ�V3�T\a��K�!^��}�H�������^�h*zj�H���,%T��[�����%F@M�A�)�0z����e��"�N|b3&�0s��uw�3
_����W���O�N��l��:��"Tƅ�X�h�R��Ϋ)�4�I�[bO����\���7��6{�/&%�&���.3A�(�eT-��ފ�%.��њ\mua�Y9`4?�-l�Ǧ4E�r͉���1S$]��$/�l�,b���_�_S��wFEN�vq�\���<�{�ZC�W�f\L�1)�7�}��r��%��)�퇒�l9�p�ܒ"M;�(t=�3;<˔��~Û�*�
)8'T�Q��-�kFM�	(��
�rbf�׏�5�tI�˯y���K��0���{�rHWL����q+OӺb��Q
�k1_�Ck��B����8��m�I�5\�3�i���I��ぽ�J)�X*�g�Vw�f�
�Gc�c�MQ�����c��QY����[{�Rt�f�M�[E����y����Կ�*Dz5�E���ك��cO�?�b׊G�~��3��{\�^�_�h� R9�jV�LV;y)`��kS�9���+�;�{}�.��9y��s�V%�n|ӵ��&��Wb���yuP>��4#@Qw�+=kA���,^-e\�]�b�xP,~�qJӿ�C1nq����Ӻ5��v�K�<@�?��$xo@l{�O>�	Kzޒ2�5Ľqg�mʀ۬��n��}أ��`Q��ďTցhn��:z��*ٴӐ�t�b�J�{�^�PY�􄳪�J:��+̄�| �ʖ�pvە;��`�f�,�a�S�MӉ{m'P���ɽ�g����+���cW�?U<��3!Y�����&��J�;iKN+�����R�ב�躨�wA��d.�GN��7��E��Q!`��@��ěCZ��ІG"�`z$S��M��0��bj��g�~�}{�t��Ų_ݶr��ܰz/
Cb�K�H X�uH�?�k>O�zk�G�C��ϳH���c \�j�Q��ގ��61Yf$��=�V�U��]�@�_l����>b�K����ƕt\�^ǅ�?�]X�_^I�R��>�v� ζ['�pԺ��>c���g��}���Z�]ou��E[�3�&�����֫�,	;��V-i���T������ݹ�O�O�p�f*|[������H)�ε VCq�Ta�b�7c�~�Y}4�l��>��[�W�[�S�;R��`�18����N��"����P��'�����E�A�6\�.?u���v�a��Ƭ�fozp��ʩ��΍�ް%���t {�\c8A��"�T��U��%8�Ϊ�@��S�F�X^�CQ�6"j7�_���k��Q��P���5�2,���'�rwٚ��{m����Z��4��m=?��UTߧ�7ro;���ʿ�����(U���o���2�2 DҏF�����P��ʬ���j'�����v���湑�>p��݀�<�3��6% �7j��$��#�?0��wr��.�H/�L�;����{��g�/�R9 6}��:��n��t�J_4̗^�a�X�!��`���Ez��%�k ��;��i�=6�S	���m`H�<��P�����6�	��L�`�p*H���w`�`����%�_\SGf_�uM�@�]��@g��l������B��@��v���@�U�p�8�Ɏ3��s\�&'h�i�(^���v��O���͓մ$�C�	J��s�z@%S.X�ir:�j�#8�����7���bGF������)i�茾����I{�ԳP�t��k}�@�&������zy�|�<zr#��p�h���q@��pf0��ܝ�� 1�ZUzn7�)B�����H�;5w����	���W�A�`y�����
������X������ZW�١�u��G��UM,ݡFs[��yڂ�J`�#���ҕdk��rG�re��AQv<�i��-WV&uXP#3]XS�d�O����J2&���)	-��[�.�)��-�*��Q��fQ�����e�9��K�ʹ����օl�g�Iun�i!�+���@2�=��g�-�˃�f5��P�ϔI)ɚƿ��SC3m�� Q\3��,IY��`��|�k)������; �j���ݩ�룼FƇ�,�� ��,�Ӂ^��y~%��-?m8ņal`k,�~
��v:F V�tGʎx��m��� Ԧ�c�n��#�bBoʺ�u��.n^=W�j���ٔ�b��~)`��e��]D6��H/I���A���r6� ��|�"F����3O�cG�&?wz�j�}�K�Y�*ScR�;�`���w{]+���� 6�Э\B��@/��)��^��Kz��it^��N,[R��wy�6��䏛A�A�~�e���l����L���s�cTS�r�B����k�G}a;��Т��O�"�
w���Z��Y��k�G�5���l��\ i�E{�-�m�>�X���I�w�L6ڱ��S�%����ǋ$]#|�.M"� "g��0� ���FAO)����V�J���Sgx�p�Ћ��ƼU��3T9�<�Y�􁌩e	_�sx�<.Px��~�xn˻���z"Z/�S���+��*�.����Ü�������$'�$zG����۷Rm�b��y�������U+��S�X�7�b��]�s��&nֽ�FEl[#s���bVJ�LFt#T*�r[�/>��0�Sq�fh>%hڶ3>����:[��
�k'�$�W���yqx�Wc�&�t>Vwn�`R9�xn�x�V�ΊE�Ra>����7�\�U���,���j�Aj�=N٘���c�=�:�r��r#�żW[?�f�Ty���
�HB�>F?����Ϙ��E�9���k��ˆO
;�#6�)b��3̼��<��{��8"���3q��%�f8�F	�Q��r�ST���]!�U��L_x�u:�����#�ś�#t�mvoA��U9�W.��PW\~����@�d�=��ў<��!SP��
d�������!b��`T6�8�����m8��ffI�X}��s�p��]/)�vd<�D3,�W���l�D��m���u4��7�[�9A�%í+��؀���y%\*�ƃ;�q��v7:v�)�n��6�i��3�KF�h��l>3������_��uX;N���oe>�W�x�zc��4[��<)�_���x>+���g$�������EW��ns��n�׃ �0+�h
������	|��hRϷ1���&1���m�����j��iThIи���	�@jq@>�������]ha� C��j��0V@z���+���/B�h���TG:75�\m��/���Fh2=���+]!Ut�{�`w�4��}����É|�b��]��=���(��g����<GK�aF��6��4�"x4y�9U�u�׀q�k5�q	��	yR�fl�TKǈ��u� ��7Kj3����������jb
���F�ܣ������"H��9���I���.�rL|
��V�{�X����";���f���g򛭺�(8A^e�7��=,-}4=��:�UIBR�]UvpCdv�l��w��i7�ʞ�����uEN��sH����!x7��k؂�xd��@%E�mz��c���h]�,� I����΁�̼>r�)����*�Џ:z�OOJP�3��K��е�o�^�{;�ߢ���0�Q� ��r�"�(l?�H,�Uu���X���S�/�J�b�=54K�Y��E�W w���[�W�]7�ϬÐ'�Q-������na��I�4�i�/pKJe4�:1f�1a��<�=�\��5�#6U_sج��?.E�_����9,�vZH���y0'C���Bh��c�l��Hv��JzP.",$Һ�q���O�8"�ԿP��W�GxH�v-߸�Tc���gJo�M�,b��X����:�����L�\�x�W!ߑ����P��Q��p�+xvL���,�|G�A0� ����l��K�R��˖����;z`���]Ge��lM&��.�k��j��첦=�����f&�(��A�̏9CcK�(>n��Mb����0֕�K��_�}�Nm�E0��w�Lܖ�[�Oa�%ŦeoSAoZ,����ulS>ʐڞĠoM�D��%��\:��6#�VR��`��c��Ս�T�[ҠUf��{&o~т����D��������%������vi�j��\5��^k��Z�{I��!w����l����ODc'^��%��3p��X�݅63+|�!\��?��+ʥ�(D��A�ĝT/  ?��`f(���̒�߉{�R�΅��kd˔�>5�͢�v{��h~&�Y.��e�8!����(7���@jw�
)hb��\0)q�Q��no��k�#���Jo�������m�;M��9�{���Z�D?�d#���iK��h
*,B�)��׉KXS �7��~i����f6L��翝0]i6M�A�M��漓�D�VK�/�hC�`�tk^����ifi���Vٰ��0{4��V��&K�A�� �	�I�t�;p�lI9鈷(-���oP�1\X^o��o߉��&������{��� ⥰��S�I(ԠKۉ�Z���T�?�m�a7��y'�*����e��-<
��<G�h���SȾ���5RMo�p{#Z���rpG�%5w�(���T����Py���Kl� �c\{��з�/�_Pa�\
���h8���v��m<â51�b����c^}̂qkZ�Q8~FJ��?C����(}n���<J/(�E���a�!���IҌedքS����3�?�`�>T!J�}|��%�F�s���X�
�.� � م���N��Ç(:�F��Lu�4���j9K@X���R=�9(�b�$�F�+�kS�����_!���ۿ'�	�:vw�*_J4�g�po��q�!�Q��d��)�3h�����_p \�N�=X\�v��˙��+l^(�D�tR��� WY,�+f�G�	[1���Ja�%�mEA/�u`���=_��I���tD�������j�ZS%E?,?�d @b�aem��������M��-Q�/<6��N4��б�i��ʓ�C��o)52+*��9��t�BE*�t�Ԭr�֏�9�+і�I�w�(����gY�H�^x��-�,K��1˖��m�D� ���3AHf�/HL���	��J�d#�pk�
nZ������%7 �'6�}r��W߿�M>A��k�'=\%�3W����9��[Q��o�0�Ӻ���M���iwiW^\[���6�J�*���u����*>��f͍_9c{�9�� �-, 7_r>J��:�H
.���_��ة~JH�_��u|���2�E~�˨�i��T�u�Y��J���A1E>����Zr`ԛ���l����0�G�F�Z�	]:���+�	mU��Y�΀"�"��/	a]� p
3�,�hU�ّ�0��3^����.���u�Ͱw8�W�,���L�y��L��PD�!l�8�<����T� *m��9T?F�w�#���pyjk��\�cF۟�
�C����B�,<���>��E�X���;9T��vNMd���L��×��ں�L���?�̉���B<�����[��j.Y*q��n{L+I�y��	�x��J����5o��&~�<T��<l�	?�~��ɂzs��P�ů�3@�M�X��d�Z���O��Ih2%UMm�N;f��#���j����\W���H^r��<����޲(�ɼ�{7�T�i
�=�f!��{���:�S?["\���?�/�*T�horX ��7�m:!Yo�Bl�-��QI��Õ�exE���tP&b�C�Y�p/�+�'�k�m]QH#��Iv�Yȗ3g}�"�=�r�e�5�I�P�0"X�C����3��$z�*2Q+4��� |V=�gM�b�<��z�25�' ��:�JErK�@���>Y�����!�OS�{�|or���ҁە"��CJ�Ó_�&��tPp#��gnVNa���G^���σ�����з�}.���Ӝ��$�%��ğƢ�V�X3ߞ�am@�a���k�9c�Z/�r�"TX�]��I�X>�_��X�y���08q�-��y$����01e�U� �6�;�Q.���������Ϛ|B������6ps��4��1�F/�2�YD��RZ��i�'�����t�`]2�h���lQ�̖���%��O|�kӑ��Lѱ\�Y���|N�T��z��$�]����K&��)|��E#��QPL�w�]������?K�˺P�w��������<w v'L]a�W��7E:Um�u�9Q�ԙ�<��͵�n�r�O����[�:������\���(���EC�͊/<qg4Ke0t}�d�?)�>�5�5�����r/R@�PjӜ��]�Rg��N���R�K�O@�/0N��S2����d����>$��;n䞁�l�`�C��D,����)fS̄�FYI��v���tbVM�[89���g��������{�5s����]��]�U���YlJqO���g�G�q]���I�c��&����3Am~dW���S[`J*/'��S�4�T��cAԃ}B�8t�	�Y+yo;��L���^au!λ�u|	�+>(W*�"���T�����l�a{�ג�d�l�n����4o�����E����i*N�T��Y9����MG�) w���.=�kz�|��GW§��=��w6l(m���#��>��F�}����R>��4��s�걩k�3���O��g�<I��\�˕wG�6tME|$a-)CɁcg^���s��:���V�yʾ����_gpfh��$�-����@3[����tb��1l��]vw(���s "0����fi�5�p���������)�?���շd�%�X�DXA�+F���Gb��3<�������\�O<8j>��B�(�ԝ��X��6mU�~'����ƿ�Y�����ER�O�� AK����F��
 a�� :�zQ'��5�Ȳ+W"] d���V�j>�/P����-y<�Q�Ŕ�BF{E�v�W��c��'6'�۝��=�(Pԝ����?�4�/��H%ծ
�av��w���?	�Vg� �H���D����U�>q��aө��40Mx�o�#$2aHD��m�g�{�v�c$"����Н<2�_2�` ��l����!lsB㜒�Ŏ�g�`	�@{��9��B�ľ�ֽ�C��Cs���G�cå%֋��b�x泩������Y^W+�"n�<m�[f��#Y�[�.OY�A�s٬X���ѱ	���z�W��x*�:����6ԎŊ���|�Q�}P�٧��9w�ʵJP��(��q����F׏R�R��rM����m$ھ��q����x#x.Tt#?'�z��] �t���*�U���h���ñԠܤǇ���9/�:D��%�ɯ��,5U@ZT��8��������rg��W�p&T[�r�t!4�Cr���@)^�~�,J�V_�6�#�h}�,:A���u��Ly��X��"�$+ S���v�,חN�F�ǳ��c��Ф��S����,Ò���֛K�L���KdM��Se���*ˎAjwhkA�Dd��IL��<���(��N��L����}�rm����f�:Hؗ�IL�E\�&(�jey�m�eD��ը�vj�����w�h����Q�6|-���
�8�5s�kL�K��"/�8�9��I�mr&O�p7���������eH�=�+V�(x��zg���ɸ��=� :�"^�u��&M^(/w��q}��b�;���>ƅ��T p�±�8��C�%_-w��E)�H��n���	Ӡ��/�7�v���ݧ��֣m����hU��l��?k,s�X�h�n��[�����F���\gNx���k�iA��WFc[�$J=7�,�S�GY;��	K,�B��W������h�_K���ٖL�BQ�8�Ԋ-ƶ��
3��?+�>Gv{�W�������q�aMQ��H�YlA��:oC-��k/O�w�|YJ.j6S�q�8
�����2~�������g��%�<���?xU��V_@��+�a0��J��Bg�}�LT�q���k������p��D>�5X����kZ�N�#3t�=��<�U�\��ND�̪d��rF�����}%Zj���AO��g�8�k�h�<$���×LJ���x�T4e5mi(A-�Q��+p��:��Bm|�험c��Z��m��3pu���H�í!mZ��8ɡ]^ie\��|�P �?����!�J�o�Yʐ ����-Y��f+� x�v�wv3(�E�$�ڀGC�G�Ϟ�4�#p��k�h(1gT��-m�!�m�B�h �L	!h����U���ފ�H#S�z.���j��X)w�Z�����!x?���Oudy�ě+ƙ
Z(H~eΊ�J ��$U��)����7Z�<�'7q�jD+X�{�  �$0I�z+����T�/d#��]�QC�>����C��������M��5�Q�� �����x���Edj��L:�@��`�Sv�1���3V�ETL�Ȳ�%��͌刚�c!�Tt��f9EL��������;q�{�.����@��Z\�ƻ#��rv��9�l�F�6��߻t�[�-�3tI[�k*;��S�ʳCi��v*�rH`}�5�j?S-;Ȭ�,���U�Z}��y�	�����:g�HGkY
=�ΝD�M|Z^�Y"a�,Y�)֔*�;sm�Șb��Z�r���Cr.�pGA�2�&�\;�}@0"r�6�<:����O�'���'9�s��q"�e�W����lj��.����`�������c'�<ө�<|o�x�| ٮ�	(Rӊ��ڹՅyE��I�>��t�ꐘP�*�^t*2h���%0�C�u$U	G��8��uM��e�j�c��� �	�.*ޞUH�8.��H���6Z(O;���:/f�yx+/�������^#(��6+���ˈ�GR������*�׍����0�I��I��F
.aS��&O�6/�
�cYb|����G�yH�2\�~J��Ӆ���CB���v��dg+���M�6����8)q&3d��a�H�uT�q�G�sLxT�p��ũ��p] �jy���AJ��R��*��܌Z����-�7�����	;
��0[ i���=�͓��s�L�:��Vh�r]�i�$=p9���Lj-�N�q�O������ ��(2�ݳi��}�ɓ���k�/P�Q�\��78LE�*�]v�0<��^���`���ik�uƶt�$FE ��d�.�B)X�p��:1p��wi���3�˚���A�ї}��HO��tS��h��>S��N��hV
�����tJ�6����nР���$~�7��<��:Y8�k:pE�A�P}44)�&��ϟ��jR��*T�q=�`y��&iAڑX�ۣ�/���d�8�'�T0.2�����Bdx��TeO��o(S�, �{L�P�!j;Qd���
��ZD�S��~�.�	Ǫ  <�j�ih���{B�̽Rm��>E|]�c+͘������yl�X��wD��r�U|!����OH�Cq��h��xd�9H>'@�ۭ�3_�#)p�i�p�Ot���S}K=<|`�]-��d�WZ����|�J���˓��S�|G`��Yq��9|,�EE�W��������ܞ�=�G�_������@u\hv)�pǆ�w2��񪆀��� Q�,膤�����t�d����$�B��R!~�rcB�yy���~�B�a��SJ3qS�җ�%{{:�3��8 �_4lJ6'#�� d�*��t�q/i�[�jwڍ܋ �'b�'��Q&�Ι͐*���ZAB���o����C����943����<k�م6Y^u�!�Қ���WF�?�s��:S.8��������O�F��'� �g���~u�Ϣ���%����W�iIȦ��]��Ӓ�P���W"1r%"%��e_�&r�K7O7��Ii�Z`z���?]�0�I���nc�#*wZT����p��ka�߭;Ii(m�t���.��k>��&o���v�0��?$A�QX��1�T	���N�,M
�?�� �n��ݷ���e�q���H�z��2����;?�z�	P˔��-��I�n�G0
Y��|�ڋ��h�7aLV(6��IoD�V������e��|^۬)��E )�@O�h*�H�Yb���d\���b�$��1#�J�:�����h���'B"@���3�.w�p�Y��m��X����0
Tᙬۓ�,)2�J �%�3�����=�s��'d�9�K>�]���c6�H�yt��85{Y!4�m�!��pZ�Ѭ�6��G}���Y��B��~X���l'ޭ���=�tqk�w&Vw�J�F�䞲#�*5�D�� W|��o�حI�x����U�X���"�?�uP/!��_őϜ������gܣL�bIK16��e�����A~୩��dd`w�)4Z#I�H=I��)
1z'a�E��!
�m����dvzd�D�a���rȲ�a(�U"��p�fYu�	������]��q�9X�u����Cspa5�¾�6yl�W��J��~�@�s�h�� Go4B�[�W������������Ξ�+�\��H&�uf
��/ cS�7�ˏ~M-����W���)����$zy��08��+wCq�p�{��F�3؈ކ8lea����:V('7�E�S@���aa;H��I6�Fa<`U�h�j2)��4��t)�+�!cԊJ@R��L����H� �쫌����(�r�=�$*g����<'ٍE�JAF�s9�=C4@��d �,���U^�So���vb��C˂S���yǍʒM˜T�q>��kO2[I:����A����_�$aT^�0�@p�o#W�e)R��PkScٗ�k5�=҆�6߯��f���D�wv ֠�<��){^��l#�8�L�R�上���S��n�,@��@�(-ᕥ.<c
�[luu.�֪�l��xC���'�/���Ѥ�6vVZ�60^��,:FI�rF��2�uk�0R��Uq�B�j%��dT��r��hR�wɼh�[��U5l�Z�?}@����Q <˴�+�WSS�w����A&h_?�[�ɰq� ����Hf7$���ťoX��"��j�?E����l.OFӌ�D�	�1��]A$d@�c/=.�[��50�`Bk��NM������S����,�A���F�[*��ʙ���4��C�%��Ƴ��z��pM[��m�2�?]
7��<�~ֿ��!�)PNЫ���Z��7qW��[�6��s$��6��_P��gߓ�f���z�3�Q}�	-ґK�T�Ya@�
�\PE����?U��`��+{��K"�42ֆT_}�h����h���z�d�\
�/�y�̒�K@	��\F_Y$�x�(B}�!��eN���=z����q�%�)q$���^q�TU���:�"5��k�@jnu�H"gB��1�>
UOe� %B�zԬQ��"���r��'�+.Z�%��FA�h�ک�<*-ֈ]���P��&x�X�D����ۀ�h��D��.�aFL��ݪg1N��QG|�a�$��mq� �h; b��ԧ磪+��]G׾^���S�ħ�"�F��;i�B�'x8��d�F|�I{A�'�.~��&�'�8<6�3����M��7���n9�6�	��Y�G��`��U��f��V���e�� l؟�z�S���F�Tac�'#ֹ7�A%�Y:�EAK�D�10��]�� \�'7��x��ad�aDd�Y�'���S:�V�9�C�GA�t�*�4��m!.ij�Z+V	F�'�DK[�����\P�olk���Q�̗8��x�����|L��^�ВZ��!���^��Yh?��A�,+�i�n��~ ��6;?ˉ��z#V@����� �d*��i��c��$��-(Kj0׼[�1�<8�O�q<�}�~�����x�f\�	X��ܭ{�3�+d�����#����c>W"r�q�ҐPM�n랴g�{���\��d������.{+��-P/>��J��|!�����H$r��U�T��E����jY�����X�8(�Ue����T*/�[�>�\��/����⸂sD��Z>JC�K0�H�}�	���a�Yi�b��lZM���Ӣ+�B�������['[c����W�J��H���j�������N���zn T�R�{<�@�����v�Z<���biMX�d��n[)P�Z{�:��:�+\	;V���7��"������A��⧫z�	d�9�ׂoJ[Y����#A�U���6.�r�����t׭����e��IXƝ`J�;#%xD2��(��бc�:̀<����$mJ�B���$�+A?�2<^O�"���<0�$}9Ò^'^	~�݆ ��J��Jm�N}\�]�}������3̜M�J�ME$R�������&3[K<9��Hy��B}�Z�'�ç�RBQ��('V��R�u�Q��nۮ�<v�%%*��CN��zu9hN<�ت����/Z##lh���'��&[e֊���ر�q�7öU��y؜��Y��H�
k�A1�0��@�:|d�������D߸��KO�M��MMs΄º/���;�j��ݓTq���
�E:��:�)��JtJ]C#�Gt����,�-X3��@�<q�vDǧLY���ۍ�M��} ̈���<;�����pVV�T����{�މ���ƍXXC�Wk�BG����2�MSW��йd��OR�+�p
�q�N"u�T�����9^Z͊!�/3!O��˵ܿ�D}�
y�d��$]Q[�� ��u��TPvv��=R�RG�&
<)�Kf]9��'R4y���u! ��R�LsǗ93q���FE��L�2����S|����^��^�&�T�]��Z ��@Sl��s#��7�W��u<O���jG�~�rY{���H J��=�,Q�����u"$l����,$���ڏ���^:���i�iN5� ٽ��Z�/�Ŕ�r�ِ��eAs<~��=�$>��l���=���i��	���X��O2 �3��]{�Y�!��_�̭zSW�=���־p����h��g�_� �K�)�`V^5��]%.v�� ted�X�v5�"����){��P�mY�(��;�P���0�&�	���qDڒ�=�� �I��+X�qc���ɞ���|n|.o[i0ސ�6�8����Ōȍo�]�a,a�T}�9��5��G�h�?�͌y����A_���.�9-�C���#�����B�/�Q��M2����L� ��yo�
�BJ�����zi�2�0��<C^ ��̍nS���ߧ�g?�7��6fL��I'p���b���"�����Er�Q1{��������KW���Rm\@ȿ � �Itӓ<��:����$��@I�w/z���)$���bMZ�����yP ��f`������I��@tw>7|YޥԞf���_��ND��B%b`X�J9��-^���KM��}_�Ѳr���st7L4@�Q��%�/w�!�����ԧ���(4��ܧ�#����Fm�E��QHНm!�a�	I�{��zݫZ�f�Q�q\���g��9ABa����/��]b�d��,�ا�t���g�pZ�cQ[Bj�M���r�&�.p��0�j��v��C����	��o�t�RN@���D懑j2�EY�R0�H6�q��π��}��FS����m��� ٌ�Fzy�]�ah��\_�D�FG���޶]�(���yDK�&ɦֶR�D�\a���lu����J���#�Ix[ޣ��nn%� ��R.˹������5�b_Ɣ~}�gX#q�X~W��:e�Ñڧ��8���Z���. �"�������[�� ]¡�{G̮��[Xb��H���x,e��?��n�} ���AƛT#�j*���k?��]�6d�]\�*M�J6�3lf�j��͍!�+$o�b�X+����Mc�)�;�F���۔y��Y���p��ܿu@˜n��ؙJ�=��Q|1�+���d��L�6p3��D13<S��Gb�w$P��xy����+W9)�ׂH-:{��M��l��2���qm�īaA�(P/X��_�-������6-�pT��v3`��1D � �3��$�;N��|m�2s�9�����ϭ��i?�J2�g\+�͵��2�(�_Lv�U�x����yb�<p?O �o��8)�Q`��Ʈ$���$�7���Z�Q۾7_h{/D6���� ,���_H������~<�8n�>�b�&��9�\3R,�������!<���T�I����j��鋍-)g0*x)�5aܔ������9մ �zz�H�M��<��v�;ٶ�)�x5-�eI�k�P(�}*���KZ��O�xum�ɩ�V�Е2	��&�}���#["�*F��)�}�$�'���z����&Mx��
�
q��S[[��5� ji��NPw>�z�Y���?ӽY�l�o +�ؒ�}Q2.�J�nv,� �>@�t�SL���ĵ�#n	����y���_��
ꓜ��
7I��xV�u	4����ξ�}~	���?}n0"��af�67|���4zs&��aR�"�ofO�'/��:���EMM�yA�z��$J�@�mCm���L�Mτ��e��s3�s2Q5��X��,��ti�d�ɵ�\-e�T #i	���#�4�D	�jz����r�\�<+ �O�P�+=������\�4z���J-��]`�'&�8�+r>E��gᚁ��nimŶ�����VKi�Rwq��E�|��a�߷�wv�e��SK�׌�Ws�g@~���x��˗[��D�O-��F��:�h���,�{tk�1�Xgl,ܴ��k�پ�o�̸��h��V#�	�A_О���˚�2�nf�N��*����t2B��-՗�>_xX���A%@���Y�q����Ҕ�{fZ��Fsj��'ӳ��Sl��� �X�cnᤛ����bfZ�q���$��=�"���!�+�fnl+�gJ&�`�I�����w[JK�����Y��C ����]�܉A��3�R����ud�Pq��J�@i�Rj[4H��U�:wk�G5��س(���E����t{���z���\��5b��SoP=ZK�U_ko�E�l]�4�~(}�V_�3�2Ԏ^`�}b�%v����,}ޖ�J��h�A�$����<��=
�_1	��d�#3<#�y��d8(��7?<�����l=Q+�Y`R=�ɛ0"G4F���J�
�P�^2Qz��g����C��O"�ڻ_򶥡W��.�G���@X�Ua�qA�/�fs� 1	}7��H"�rk�B)��;H~�P�/�|h����0�������)���t.�8�.��Ǽ����Յ4W`(��Y@�T�YH~ii#���/�j�a�#�{�}��$vZ�;]��=��%V(�}�<��P��d��G��Ap�M�3+��I$��%��?�pGƃ���@�%�rF4����X�pK'�--��<��:p4Y�+����ؿ/`+��+�m�����W������|ۿY)�G���̠Q�Sq�{&7�+�lj#����po��}���>�k���&��v��5��jhާ��v,[I�ܦ�L���z��%&OXJ�^Cc��گ�g��]V�S#C���\V^I��[���y ]�uC�8 g�*�� �HX$1��Hn�G�G����_��t/��v\�7�����x'i����I,�٦CI�+,�Y夃�`�]��Ŝ��^�k���4��^Ώ,d���*[��9�g)"�E�j�v�B �R�i�Z
ԍU�إ������iP��OvB��/�חF_j��.�������ݙ��oK��3�Z���`��^U!�B��#��f���հy�/����z�fK&�k�m�\'.:��JG�Ϫ/��B����ͼ�e #���K�@D!~����r�%w�gQ=д��I+=%�mrK�~�tW��IU��l�.Of�u�h�J:�Y����%��X�d���ϖ����1j��2I��{\_W?<�ly�/�3�lC=5��xW��؂����T���kz���J>0�ٷ]J9Y�k�$0�{��E�Nd�|�<�hႺ4��%����bo1[뽲��lM���pAa׆?D�u���%����UK^?/�Sށ����kLs��%�l	p�����)x-���'�=��W��	�%VgS\�H��/�pZ/�oQ8꟢S'*֗����D�Z.�F��-����$�7Z�?��uB)�Aڄ���M�jm1Pjr��J�+7,
&�#+C�;y���]xj�g�u@v���x�E�Kzc㴞Ta��~)�+\����Mef��U&��Jv��4�v̈i|kn�vDG��ʟpgI��U���SL��T@e�lуE��2��/�K�d�!�fӛ�j�w&;e,vɋ�u9mg�F� O)���	{�pCTiex�6'&��J(��(�����X�=ϳ�d�x�e���8�ϒEp�C�1����˕j`��/ ő�J0�ա�.G~.�{;���H�X���ӿ�.h6n���6~�0�<Sр�ԶB�Oa�Kՙ�A��p����8ݼ��QP���	j�yS��K�����l�څ��u/�!K"�{x^�]@�:ң�T�-�S�m�-���p5r��ׂ;�(/�&������)��m��Tz����a9�ՙ�5�<��������EE��/Y�����L�O]�ǽ����ǥ,��SED��]KH�A/��P�GYRG'����a3��K���VK�����]Uc�yF�K�NUj(0g!>c'���E�A�F�;�Gye.�(�<�I�q>��!)fq�&����!�,"�gb�4k+�t�N�wz-��"��yǴ4ץ-��Sp\y}�qܜ�4-��* Y�O�E�u\�>��"oa;qp}*��%�Ĵ�mx� �$�2��?��"JSg���K=
�W�ؙ��I�z��D΁>o/�Q��}�Ě�#+K�oa'ЫΧ��_:G��ba�Z;Eݞu�:�����vs�[�?��������S��>���B$�h�H�r����Ɏ��0K��sa2õ�/����l,���|��F0(a�2RجN"c��s0$RWm�p�����O䤤�~�^_<�$t�,��f�0��X�]�6ͼX�ʻ���/��/����1��:4>���D4Q�wy,g�<2B�3���S�`wAt�L?+�W�x%��X_�[�){��N�T��v*��/4��W+d��'P�Y\��i109�H��9]*��˿�+,��Q"���Re�*��#��{WT0�N��ܑ��Z~g���H�-�w�D��e9�O���~7�Hs`Z�zك�w��&��ǡ���ӧ,=���������w�n������O=������ �S<х|�q��C�Yi��UH����h�5�YRȰ�"�%�!}���C����`�2������/������14�ޖq4�
�@�2�x��1���%i���R�����f�Oeg-�`��C���o�lɼ;�a�U�&�qyI3��a^�`�b%��8R��1/S{P�/�D�
�zz;�DO/4�z�A��yD.=�
��3·�v��I�%&z}=����T�휂��0�ޥ�`y�����$-y@�2bL���ź��d��ЂN��=�-�C���{��f{��CFn���iB����䧛,��e���p�IM���-0��wy*M����H�͆��ezp���r��PLY��{n>{�rN4��9�)
7G'F�s�Z���<��=��"��)�o&1C^M�ph,͢�{^v����h¢	dA�omVQE��.X.m\I��}rְ6i�SГ���Ӫ~-6�ĝ�_��d���Pz�Wz?G�D�!�6Wjk)�I����;d8�S!x��X�&�g q̲�B��У֮��!-��>\Z��q�B�! ��VE����՝�^n�Լn������
��Wwψ�y�*����@�DE������u���RM�^h*��%9f7Ss��I�pânN,ڦݻ
˞���Y�DP��o�u.EJ%�<�rR5�O��wJߣ%#�'�۝9Q�$ۙ�4ƹ{S��HgQw���T�1*�֚�=S�=�¨�2b:�˺Bǜ8��Bs��wD�:��]b@&�#�q�ň*y
R��n%%��X_��7P�Դ]�q2օc{��#.ϤqB��ru_�b�4���O���X���!�U �se�.��3�"=������'t8��c?w��f�q�.<���eNe�{R�WU��p':!dl���I p��$���pa^��G]t�]�����w��j7�� �9�=	Qv���N�t%"�!�y%#�5�������{�ր���{�9'�����,�M��A]��į��6'OA�ئ2B�.7�r����q����Uhv^�f��S���Ec��ǻԶp���x)��4Gö��~���7UqY�$>�7�i��L(:��ax�6��M��
b���?7�ԐSB��ڒlͩ'�Cq��F��Z��>�Dh.U��pr�[��犠�.W�)X���^���\�롉"�jJ'Q�#T}\-
~B��JH� ��2��+��K1��-�K��d���(�&ky�tb'�&w�!�~֏g�jI8,��V��O ��zf������x:z<s�Z��Co�{�Z,�³��kŞ��6�˅Ϝ?�C<��Z���i���%P�%�L�ۇ�p�� r5FI��[�v}Q����c����^�!?���%����_`�G.t���>�2��F�Y�F�P �.��<?\�W"�3ۭ �r�3�i�ڜ z},���sԗ�1Cc7 �o�����X�13?gW9|����/�3L���"�);ӊ��b��}��&L=���6��<��,1��k�G���N4N|ق��5!�W1� -1A3�B�d~j��� �X[8���o�H7�;(	AS��u��n�j���1nж��x����?�l��R�^���{�)�<'1�K�
��'Bw?�����3�"���&��e�4�ef��# ]9Q��� �-�k�i=d@5�7�#DO
x�]��Z�x�.f�`Zhr(˪�dGz��1�a]��С�qRӯ��`�s]w�H %������߉ I�ȏmɊ��	ee���`۟��ջ�w�L�qG(ᷜ�?�:�j,"��O�,�ùT�kA�#��o��@�]EE�7��x=qg�Q��+j���~��;p[�p�$��R����
?�-��_t>+ U���TeXgE��9�P�L��T�(9d����M��Ya�`��59�W�O(ݭ&�V]���l �J�4�E!~�PN�^�e	���'���(À1�� �X����{m �4����ѵSP��� �y6�9��s��v��:���BW�9��7ID�����An�o+i��6�uLƁ�|�VC�v޳Os`��������ꥩ|W{����a9�i7����:l;a�.��4��ޥHC6��26];�{�U�|�fZ����1�/��
�h�<��Vk�=@o�e#�g����h�����g.H�Y���L�Lb��~�\'đ��>���C�����(���5����>�j)�gq\W�:I������ɒ�6��[���,�U��Yz�V�S�4�V�ch����s����\@{�Yk�2�(������7�����J$��3����T�Ȝ�;���1-j	3�l�	7	����e�ز��}8����S��˰q�w��	���}A)��c7(a#��� ��@�Ū0�$�3^�6��vV���� �2�'-���du�$��O��S\u���a�=X^޿�_ꌖ�X�3D��2cB��QO�-��,���Ry����fJ����TE
�����
Q<`:�,����ﰀ�T�?sҜl*!&��!]'t+ܶ�!p��ߠN���1���D���`^J�T��J��.��̵��B��Bߘ��[�9"ðx��.:\�YH�mu��vZy:�=2̭X|Y6���HNsa��-��Ņ�dL�KLk��$̾Wѿ4Ô��D�u�Jo�^����� X��o���ߡ��a)�P���M�����;��D�섿������C7�E��~$Nۧ�Xy�M�?��˗,���Jdm�$CJs.�f�1Q`��������-�2�%����z�.^�JB���5�i5��^1�,]�F�M��WR����;ٖ3�fI4�/�@�� 0���p|�h(F����q}�z���l�6��3d�=�`L���I+'��Ul�q�'�P�u���w��n�����#��o����6�+կ�Й�`����c��|*�T�y9t�Â	��4�n/���*�/"����V=ϗ�L�����iI��&��ԕDC-r��D5(�ͬX�2��������Q�{"I�_y�����6Ôsذ��w2p���3�k҆fp�$�]���S��B\���(��]MM�t��r�F'�z4�҃��Z+Ks�j�3�U��l9��X����;<]Q�F_�͍�T�YKeheJu�eg�gDkCp��+�SX��S�%�3�	m�tRH2�9
�3�q�Jb)���jeS����:N�"�Xi{�n�@��Yp��Z�K�,3~�7 #�S� 8��LY�w�0��"��ݦ������	��ց�˵r?ׇ�P�=tL5Sj�ěysIi�
9ו�%i�bs�!5�bm����QE%�4�?��Hs�'���8�F(�PzTj4b2ʒ����f��:��%2�5[��Fo��C��L�����^�]#BG?[�� �s�C��	G��I̶��H��5�8ETG�N!(aJpd�ߓvf�B�5J������&��-}P�I��"|�m�����\5b���3��&�Y�&>x8��b%����9��ϝ��Kn�^*M����w�?"h6>�;d�FrU��9s�&��g�9jڜ7�Z���k��Tš����)1Z"�H�Ms��b�d����0'j�rc���wÏk�އ�>G5\�	N���D�9���� :���l����mIm���h̒��qb�`YF����"Ih`wCP������ I�T&F������W�T�:�0�Z��v�$�gO�KςH��!,�2fm:�j��X��>"1X�M�߶$tG!ԗ��=ckc�8���o�N����b�+��:"�iX�/� ��o�?����߹{�iP!�ǥ��0�Y6RF��~��ː܏|�]u85��\�9����C:�iv�fX�L��H����8�K�9�p��o࿂Md0�K��.��^lm0-�Lᖥ*e�U��Z�*���k�5��-g�.�/]��H���M�@���K�Ğ�w:P����.I������
6��^�	��r���ruB)�kZ����W�P�6BqkR���D���X�A��Po���t��W���霜����-�b5�g����q�j+��eM�ͺ�6�8�t�)�/.]���d���X9���_�.m	��_8��"��z}e��
�2F��yy�����~vb@��JշZ��a��r���y6����xN�������'_��{�;���b�;�\�L�IV0���	G�_�B���p�nJ̗�3O�Jc~l�l�TD_�bB��t����VYۃ��\g!�K m�L%U�-]V�.r�3[?o�`V|���������j�^�Z�C[cP��*��ܙ�@�����?}�'�A�OX.�ͪxH{l��>Ѣ%��doA����}�I������,yXñ4��
�Bx��K�.K+Y�6��7����I�;M�X7^���5$}�o(��#����{�ɉ��K��F���"%:�1�1Y�)�
p@h݁���Δ��L�ybJ��_�g��@�ej�5��{Ku�ǆ��]�w
��:���2kPpѷc��S�LK�M�90K��:��7to*})��������3MuFj�gQW���7����'̖'`��.�ܨe��X�*��-3��ɭ�[�j��X~8����ں�N��p��3�W ����>�2�0�V�}y�/�tV�FQӈ(��޸�����u���J`�xtd9+����oo:�����R����v��G�〴� NY���~E�w�b�8��{~�C qz�J�,�6m��v_��Lp��o&�����cdQj�xW4�!&�tV�k6:2mY\��^+l�g��\�왅$�-�/0��P��DL�z��\H�5���~	�B�O���9�4L	����֚����_\ĮF·�s6G�\)���(���V|��bk�*�����u&m�.��y^�Nq]�\}��`�1>2?��~�*�ҍ"�i�������[�UW��W� ���S��Q�\���b�YQ�zG��~�̒;�x�vT��o��\���发�I���}�������rU�ךE�}�XJ	�{L����"����c�(�^�7M���j �����-�=�-��ML��.��c�!��O��ݳǥش��Z��ҫ�N(xo�)�r�n�G8��{���j��ljo��J.��;]rv�S<��N��P��]�ؘ:�EQH����݅h-����H���i���}y������@���H6����Sx��W�-�u�7���{ ����I�s?