--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity AV_Config_avalon_av_config_slave_arbitrator is 
        port (
              -- inputs:
                 signal AV_Config_avalon_av_config_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal AV_Config_avalon_av_config_slave_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal AV_Config_avalon_av_config_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal AV_Config_avalon_av_config_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal AV_Config_avalon_av_config_slave_read : OUT STD_LOGIC;
                 signal AV_Config_avalon_av_config_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal AV_Config_avalon_av_config_slave_reset : OUT STD_LOGIC;
                 signal AV_Config_avalon_av_config_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal AV_Config_avalon_av_config_slave_write : OUT STD_LOGIC;
                 signal AV_Config_avalon_av_config_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_granted_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                 signal d1_AV_Config_avalon_av_config_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : OUT STD_LOGIC
              );
end entity AV_Config_avalon_av_config_slave_arbitrator;


architecture europa of AV_Config_avalon_av_config_slave_arbitrator is
                signal AV_Config_avalon_av_config_slave_allgrants :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_any_continuerequest :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_arb_counter_enable :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_begins_xfer :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_end_xfer :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_firsttransfer :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_grant_vector :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_in_a_read_cycle :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_in_a_write_cycle :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_master_qreq_vector :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_non_bursting_master_requests :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_reg_firsttransfer :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_slavearbiterlockenable :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_unreg_firsttransfer :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_waits_for_read :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_waits_for_write :  STD_LOGIC;
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_AV_Config_avalon_av_config_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_AV_Config_avalon_av_config_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_AV_Config_avalon_av_config_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT AV_Config_avalon_av_config_slave_end_xfer;
    end if;

  end process;

  AV_Config_avalon_av_config_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave);
  --assign AV_Config_avalon_av_config_slave_readdata_from_sa = AV_Config_avalon_av_config_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  AV_Config_avalon_av_config_slave_readdata_from_sa <= AV_Config_avalon_av_config_slave_readdata;
  internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000011000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign AV_Config_avalon_av_config_slave_waitrequest_from_sa = AV_Config_avalon_av_config_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_AV_Config_avalon_av_config_slave_waitrequest_from_sa <= AV_Config_avalon_av_config_slave_waitrequest;
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave <= CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register_in;
  --AV_Config_avalon_av_config_slave_arb_share_counter set values, which is an e_mux
  AV_Config_avalon_av_config_slave_arb_share_set_values <= std_logic_vector'("001");
  --AV_Config_avalon_av_config_slave_non_bursting_master_requests mux, which is an e_mux
  AV_Config_avalon_av_config_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave;
  --AV_Config_avalon_av_config_slave_any_bursting_master_saved_grant mux, which is an e_mux
  AV_Config_avalon_av_config_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --AV_Config_avalon_av_config_slave_arb_share_counter_next_value assignment, which is an e_assign
  AV_Config_avalon_av_config_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(AV_Config_avalon_av_config_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (AV_Config_avalon_av_config_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(AV_Config_avalon_av_config_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (AV_Config_avalon_av_config_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --AV_Config_avalon_av_config_slave_allgrants all slave grants, which is an e_mux
  AV_Config_avalon_av_config_slave_allgrants <= AV_Config_avalon_av_config_slave_grant_vector;
  --AV_Config_avalon_av_config_slave_end_xfer assignment, which is an e_assign
  AV_Config_avalon_av_config_slave_end_xfer <= NOT ((AV_Config_avalon_av_config_slave_waits_for_read OR AV_Config_avalon_av_config_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave <= AV_Config_avalon_av_config_slave_end_xfer AND (((NOT AV_Config_avalon_av_config_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --AV_Config_avalon_av_config_slave_arb_share_counter arbitration counter enable, which is an e_assign
  AV_Config_avalon_av_config_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave AND AV_Config_avalon_av_config_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave AND NOT AV_Config_avalon_av_config_slave_non_bursting_master_requests));
  --AV_Config_avalon_av_config_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      AV_Config_avalon_av_config_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(AV_Config_avalon_av_config_slave_arb_counter_enable) = '1' then 
        AV_Config_avalon_av_config_slave_arb_share_counter <= AV_Config_avalon_av_config_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --AV_Config_avalon_av_config_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      AV_Config_avalon_av_config_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((AV_Config_avalon_av_config_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave)) OR ((end_xfer_arb_share_counter_term_AV_Config_avalon_av_config_slave AND NOT AV_Config_avalon_av_config_slave_non_bursting_master_requests)))) = '1' then 
        AV_Config_avalon_av_config_slave_slavearbiterlockenable <= or_reduce(AV_Config_avalon_av_config_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master AV_Config/avalon_av_config_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= AV_Config_avalon_av_config_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --AV_Config_avalon_av_config_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  AV_Config_avalon_av_config_slave_slavearbiterlockenable2 <= or_reduce(AV_Config_avalon_av_config_slave_arb_share_counter_next_value);
  --CPU/data_master AV_Config/avalon_av_config_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= AV_Config_avalon_av_config_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --AV_Config_avalon_av_config_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  AV_Config_avalon_av_config_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register_in <= ((internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave AND CPU_data_master_read) AND NOT AV_Config_avalon_av_config_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register <= p1_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave, which is an e_mux
  CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave <= CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave_shift_register;
  --AV_Config_avalon_av_config_slave_writedata mux, which is an e_mux
  AV_Config_avalon_av_config_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave;
  --CPU/data_master saved-grant AV_Config/avalon_av_config_slave, which is an e_assign
  CPU_data_master_saved_grant_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave;
  --allow new arb cycle for AV_Config/avalon_av_config_slave, which is an e_assign
  AV_Config_avalon_av_config_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  AV_Config_avalon_av_config_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  AV_Config_avalon_av_config_slave_master_qreq_vector <= std_logic'('1');
  --~AV_Config_avalon_av_config_slave_reset assignment, which is an e_assign
  AV_Config_avalon_av_config_slave_reset <= NOT reset_n;
  --AV_Config_avalon_av_config_slave_firsttransfer first transaction, which is an e_assign
  AV_Config_avalon_av_config_slave_firsttransfer <= A_WE_StdLogic((std_logic'(AV_Config_avalon_av_config_slave_begins_xfer) = '1'), AV_Config_avalon_av_config_slave_unreg_firsttransfer, AV_Config_avalon_av_config_slave_reg_firsttransfer);
  --AV_Config_avalon_av_config_slave_unreg_firsttransfer first transaction, which is an e_assign
  AV_Config_avalon_av_config_slave_unreg_firsttransfer <= NOT ((AV_Config_avalon_av_config_slave_slavearbiterlockenable AND AV_Config_avalon_av_config_slave_any_continuerequest));
  --AV_Config_avalon_av_config_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      AV_Config_avalon_av_config_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(AV_Config_avalon_av_config_slave_begins_xfer) = '1' then 
        AV_Config_avalon_av_config_slave_reg_firsttransfer <= AV_Config_avalon_av_config_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --AV_Config_avalon_av_config_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  AV_Config_avalon_av_config_slave_beginbursttransfer_internal <= AV_Config_avalon_av_config_slave_begins_xfer;
  --AV_Config_avalon_av_config_slave_read assignment, which is an e_mux
  AV_Config_avalon_av_config_slave_read <= internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave AND CPU_data_master_read;
  --AV_Config_avalon_av_config_slave_write assignment, which is an e_mux
  AV_Config_avalon_av_config_slave_write <= internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave AND CPU_data_master_write;
  shifted_address_to_AV_Config_avalon_av_config_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --AV_Config_avalon_av_config_slave_address mux, which is an e_mux
  AV_Config_avalon_av_config_slave_address <= A_EXT (A_SRL(shifted_address_to_AV_Config_avalon_av_config_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_AV_Config_avalon_av_config_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_AV_Config_avalon_av_config_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_AV_Config_avalon_av_config_slave_end_xfer <= AV_Config_avalon_av_config_slave_end_xfer;
    end if;

  end process;

  --AV_Config_avalon_av_config_slave_waits_for_read in a cycle, which is an e_mux
  AV_Config_avalon_av_config_slave_waits_for_read <= AV_Config_avalon_av_config_slave_in_a_read_cycle AND internal_AV_Config_avalon_av_config_slave_waitrequest_from_sa;
  --AV_Config_avalon_av_config_slave_in_a_read_cycle assignment, which is an e_assign
  AV_Config_avalon_av_config_slave_in_a_read_cycle <= internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= AV_Config_avalon_av_config_slave_in_a_read_cycle;
  --AV_Config_avalon_av_config_slave_waits_for_write in a cycle, which is an e_mux
  AV_Config_avalon_av_config_slave_waits_for_write <= AV_Config_avalon_av_config_slave_in_a_write_cycle AND internal_AV_Config_avalon_av_config_slave_waitrequest_from_sa;
  --AV_Config_avalon_av_config_slave_in_a_write_cycle assignment, which is an e_assign
  AV_Config_avalon_av_config_slave_in_a_write_cycle <= internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= AV_Config_avalon_av_config_slave_in_a_write_cycle;
  wait_for_AV_Config_avalon_av_config_slave_counter <= std_logic'('0');
  --AV_Config_avalon_av_config_slave_byteenable byte enable port mux, which is an e_mux
  AV_Config_avalon_av_config_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  AV_Config_avalon_av_config_slave_waitrequest_from_sa <= internal_AV_Config_avalon_av_config_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  CPU_data_master_granted_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_granted_AV_Config_avalon_av_config_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_AV_Config_avalon_av_config_slave <= internal_CPU_data_master_requests_AV_Config_avalon_av_config_slave;
--synthesis translate_off
    --AV_Config/avalon_av_config_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Alpha_Blending_avalon_background_sink_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_background_sink_ready : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Pixel_Scaler_avalon_scaler_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Alpha_Blending_avalon_background_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal Alpha_Blending_avalon_background_sink_endofpacket : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_background_sink_ready_from_sa : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_background_sink_startofpacket : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_background_sink_valid : OUT STD_LOGIC
              );
end entity Alpha_Blending_avalon_background_sink_arbitrator;


architecture europa of Alpha_Blending_avalon_background_sink_arbitrator is

begin

  --mux Alpha_Blending_avalon_background_sink_data, which is an e_mux
  Alpha_Blending_avalon_background_sink_data <= VGA_Pixel_Scaler_avalon_scaler_source_data;
  --mux Alpha_Blending_avalon_background_sink_endofpacket, which is an e_mux
  Alpha_Blending_avalon_background_sink_endofpacket <= VGA_Pixel_Scaler_avalon_scaler_source_endofpacket;
  --assign Alpha_Blending_avalon_background_sink_ready_from_sa = Alpha_Blending_avalon_background_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  Alpha_Blending_avalon_background_sink_ready_from_sa <= Alpha_Blending_avalon_background_sink_ready;
  --mux Alpha_Blending_avalon_background_sink_startofpacket, which is an e_mux
  Alpha_Blending_avalon_background_sink_startofpacket <= VGA_Pixel_Scaler_avalon_scaler_source_startofpacket;
  --mux Alpha_Blending_avalon_background_sink_valid, which is an e_mux
  Alpha_Blending_avalon_background_sink_valid <= VGA_Pixel_Scaler_avalon_scaler_source_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Alpha_Blending_avalon_foreground_sink_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_foreground_sink_ready : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Alpha_Blending_avalon_foreground_sink_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal Alpha_Blending_avalon_foreground_sink_endofpacket : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_foreground_sink_ready_from_sa : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_foreground_sink_reset : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_foreground_sink_startofpacket : OUT STD_LOGIC;
                 signal Alpha_Blending_avalon_foreground_sink_valid : OUT STD_LOGIC
              );
end entity Alpha_Blending_avalon_foreground_sink_arbitrator;


architecture europa of Alpha_Blending_avalon_foreground_sink_arbitrator is

begin

  --mux Alpha_Blending_avalon_foreground_sink_data, which is an e_mux
  Alpha_Blending_avalon_foreground_sink_data <= VGA_Char_Buffer_avalon_char_source_data;
  --mux Alpha_Blending_avalon_foreground_sink_endofpacket, which is an e_mux
  Alpha_Blending_avalon_foreground_sink_endofpacket <= VGA_Char_Buffer_avalon_char_source_endofpacket;
  --assign Alpha_Blending_avalon_foreground_sink_ready_from_sa = Alpha_Blending_avalon_foreground_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  Alpha_Blending_avalon_foreground_sink_ready_from_sa <= Alpha_Blending_avalon_foreground_sink_ready;
  --mux Alpha_Blending_avalon_foreground_sink_startofpacket, which is an e_mux
  Alpha_Blending_avalon_foreground_sink_startofpacket <= VGA_Char_Buffer_avalon_char_source_startofpacket;
  --mux Alpha_Blending_avalon_foreground_sink_valid, which is an e_mux
  Alpha_Blending_avalon_foreground_sink_valid <= VGA_Char_Buffer_avalon_char_source_valid;
  --~Alpha_Blending_avalon_foreground_sink_reset assignment, which is an e_assign
  Alpha_Blending_avalon_foreground_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Alpha_Blending_avalon_blended_source_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal Alpha_Blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                 signal Alpha_Blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                 signal Alpha_Blending_avalon_blended_source_valid : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Alpha_Blending_avalon_blended_source_ready : OUT STD_LOGIC
              );
end entity Alpha_Blending_avalon_blended_source_arbitrator;


architecture europa of Alpha_Blending_avalon_blended_source_arbitrator is

begin

  --mux Alpha_Blending_avalon_blended_source_ready, which is an e_mux
  Alpha_Blending_avalon_blended_source_ready <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Audio_avalon_audio_slave_arbitrator is 
        port (
              -- inputs:
                 signal Audio_avalon_audio_slave_irq : IN STD_LOGIC;
                 signal Audio_avalon_audio_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Audio_avalon_audio_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Audio_avalon_audio_slave_chipselect : OUT STD_LOGIC;
                 signal Audio_avalon_audio_slave_irq_from_sa : OUT STD_LOGIC;
                 signal Audio_avalon_audio_slave_read : OUT STD_LOGIC;
                 signal Audio_avalon_audio_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Audio_avalon_audio_slave_reset : OUT STD_LOGIC;
                 signal Audio_avalon_audio_slave_write : OUT STD_LOGIC;
                 signal Audio_avalon_audio_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_granted_Audio_avalon_audio_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Audio_avalon_audio_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Audio_avalon_audio_slave : OUT STD_LOGIC;
                 signal d1_Audio_avalon_audio_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave : OUT STD_LOGIC
              );
end entity Audio_avalon_audio_slave_arbitrator;


architecture europa of Audio_avalon_audio_slave_arbitrator is
                signal Audio_avalon_audio_slave_allgrants :  STD_LOGIC;
                signal Audio_avalon_audio_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Audio_avalon_audio_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Audio_avalon_audio_slave_any_continuerequest :  STD_LOGIC;
                signal Audio_avalon_audio_slave_arb_counter_enable :  STD_LOGIC;
                signal Audio_avalon_audio_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Audio_avalon_audio_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Audio_avalon_audio_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Audio_avalon_audio_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Audio_avalon_audio_slave_begins_xfer :  STD_LOGIC;
                signal Audio_avalon_audio_slave_end_xfer :  STD_LOGIC;
                signal Audio_avalon_audio_slave_firsttransfer :  STD_LOGIC;
                signal Audio_avalon_audio_slave_grant_vector :  STD_LOGIC;
                signal Audio_avalon_audio_slave_in_a_read_cycle :  STD_LOGIC;
                signal Audio_avalon_audio_slave_in_a_write_cycle :  STD_LOGIC;
                signal Audio_avalon_audio_slave_master_qreq_vector :  STD_LOGIC;
                signal Audio_avalon_audio_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Audio_avalon_audio_slave_reg_firsttransfer :  STD_LOGIC;
                signal Audio_avalon_audio_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Audio_avalon_audio_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Audio_avalon_audio_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Audio_avalon_audio_slave_waits_for_read :  STD_LOGIC;
                signal Audio_avalon_audio_slave_waits_for_write :  STD_LOGIC;
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Audio_avalon_audio_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Audio_avalon_audio_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Audio_avalon_audio_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Audio_avalon_audio_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Audio_avalon_audio_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Audio_avalon_audio_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Audio_avalon_audio_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Audio_avalon_audio_slave_end_xfer;
    end if;

  end process;

  Audio_avalon_audio_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Audio_avalon_audio_slave);
  --assign Audio_avalon_audio_slave_readdata_from_sa = Audio_avalon_audio_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Audio_avalon_audio_slave_readdata_from_sa <= Audio_avalon_audio_slave_readdata;
  internal_CPU_data_master_requests_Audio_avalon_audio_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000011000001000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave <= CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register_in;
  --Audio_avalon_audio_slave_arb_share_counter set values, which is an e_mux
  Audio_avalon_audio_slave_arb_share_set_values <= std_logic_vector'("001");
  --Audio_avalon_audio_slave_non_bursting_master_requests mux, which is an e_mux
  Audio_avalon_audio_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Audio_avalon_audio_slave;
  --Audio_avalon_audio_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Audio_avalon_audio_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Audio_avalon_audio_slave_arb_share_counter_next_value assignment, which is an e_assign
  Audio_avalon_audio_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Audio_avalon_audio_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Audio_avalon_audio_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Audio_avalon_audio_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Audio_avalon_audio_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Audio_avalon_audio_slave_allgrants all slave grants, which is an e_mux
  Audio_avalon_audio_slave_allgrants <= Audio_avalon_audio_slave_grant_vector;
  --Audio_avalon_audio_slave_end_xfer assignment, which is an e_assign
  Audio_avalon_audio_slave_end_xfer <= NOT ((Audio_avalon_audio_slave_waits_for_read OR Audio_avalon_audio_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Audio_avalon_audio_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Audio_avalon_audio_slave <= Audio_avalon_audio_slave_end_xfer AND (((NOT Audio_avalon_audio_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Audio_avalon_audio_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Audio_avalon_audio_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Audio_avalon_audio_slave AND Audio_avalon_audio_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Audio_avalon_audio_slave AND NOT Audio_avalon_audio_slave_non_bursting_master_requests));
  --Audio_avalon_audio_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Audio_avalon_audio_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Audio_avalon_audio_slave_arb_counter_enable) = '1' then 
        Audio_avalon_audio_slave_arb_share_counter <= Audio_avalon_audio_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Audio_avalon_audio_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Audio_avalon_audio_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Audio_avalon_audio_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Audio_avalon_audio_slave)) OR ((end_xfer_arb_share_counter_term_Audio_avalon_audio_slave AND NOT Audio_avalon_audio_slave_non_bursting_master_requests)))) = '1' then 
        Audio_avalon_audio_slave_slavearbiterlockenable <= or_reduce(Audio_avalon_audio_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Audio/avalon_audio_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Audio_avalon_audio_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Audio_avalon_audio_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Audio_avalon_audio_slave_slavearbiterlockenable2 <= or_reduce(Audio_avalon_audio_slave_arb_share_counter_next_value);
  --CPU/data_master Audio/avalon_audio_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Audio_avalon_audio_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Audio_avalon_audio_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Audio_avalon_audio_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Audio_avalon_audio_slave <= internal_CPU_data_master_requests_Audio_avalon_audio_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register_in <= ((internal_CPU_data_master_granted_Audio_avalon_audio_slave AND CPU_data_master_read) AND NOT Audio_avalon_audio_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register <= p1_CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Audio_avalon_audio_slave, which is an e_mux
  CPU_data_master_read_data_valid_Audio_avalon_audio_slave <= CPU_data_master_read_data_valid_Audio_avalon_audio_slave_shift_register;
  --Audio_avalon_audio_slave_writedata mux, which is an e_mux
  Audio_avalon_audio_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Audio_avalon_audio_slave <= internal_CPU_data_master_qualified_request_Audio_avalon_audio_slave;
  --CPU/data_master saved-grant Audio/avalon_audio_slave, which is an e_assign
  CPU_data_master_saved_grant_Audio_avalon_audio_slave <= internal_CPU_data_master_requests_Audio_avalon_audio_slave;
  --allow new arb cycle for Audio/avalon_audio_slave, which is an e_assign
  Audio_avalon_audio_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Audio_avalon_audio_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Audio_avalon_audio_slave_master_qreq_vector <= std_logic'('1');
  --~Audio_avalon_audio_slave_reset assignment, which is an e_assign
  Audio_avalon_audio_slave_reset <= NOT reset_n;
  Audio_avalon_audio_slave_chipselect <= internal_CPU_data_master_granted_Audio_avalon_audio_slave;
  --Audio_avalon_audio_slave_firsttransfer first transaction, which is an e_assign
  Audio_avalon_audio_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Audio_avalon_audio_slave_begins_xfer) = '1'), Audio_avalon_audio_slave_unreg_firsttransfer, Audio_avalon_audio_slave_reg_firsttransfer);
  --Audio_avalon_audio_slave_unreg_firsttransfer first transaction, which is an e_assign
  Audio_avalon_audio_slave_unreg_firsttransfer <= NOT ((Audio_avalon_audio_slave_slavearbiterlockenable AND Audio_avalon_audio_slave_any_continuerequest));
  --Audio_avalon_audio_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Audio_avalon_audio_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Audio_avalon_audio_slave_begins_xfer) = '1' then 
        Audio_avalon_audio_slave_reg_firsttransfer <= Audio_avalon_audio_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Audio_avalon_audio_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Audio_avalon_audio_slave_beginbursttransfer_internal <= Audio_avalon_audio_slave_begins_xfer;
  --Audio_avalon_audio_slave_read assignment, which is an e_mux
  Audio_avalon_audio_slave_read <= internal_CPU_data_master_granted_Audio_avalon_audio_slave AND CPU_data_master_read;
  --Audio_avalon_audio_slave_write assignment, which is an e_mux
  Audio_avalon_audio_slave_write <= internal_CPU_data_master_granted_Audio_avalon_audio_slave AND CPU_data_master_write;
  shifted_address_to_Audio_avalon_audio_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Audio_avalon_audio_slave_address mux, which is an e_mux
  Audio_avalon_audio_slave_address <= A_EXT (A_SRL(shifted_address_to_Audio_avalon_audio_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Audio_avalon_audio_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Audio_avalon_audio_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Audio_avalon_audio_slave_end_xfer <= Audio_avalon_audio_slave_end_xfer;
    end if;

  end process;

  --Audio_avalon_audio_slave_waits_for_read in a cycle, which is an e_mux
  Audio_avalon_audio_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Audio_avalon_audio_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Audio_avalon_audio_slave_in_a_read_cycle assignment, which is an e_assign
  Audio_avalon_audio_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Audio_avalon_audio_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Audio_avalon_audio_slave_in_a_read_cycle;
  --Audio_avalon_audio_slave_waits_for_write in a cycle, which is an e_mux
  Audio_avalon_audio_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Audio_avalon_audio_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Audio_avalon_audio_slave_in_a_write_cycle assignment, which is an e_assign
  Audio_avalon_audio_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Audio_avalon_audio_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Audio_avalon_audio_slave_in_a_write_cycle;
  wait_for_Audio_avalon_audio_slave_counter <= std_logic'('0');
  --assign Audio_avalon_audio_slave_irq_from_sa = Audio_avalon_audio_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Audio_avalon_audio_slave_irq_from_sa <= Audio_avalon_audio_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Audio_avalon_audio_slave <= internal_CPU_data_master_granted_Audio_avalon_audio_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Audio_avalon_audio_slave <= internal_CPU_data_master_qualified_request_Audio_avalon_audio_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Audio_avalon_audio_slave <= internal_CPU_data_master_requests_Audio_avalon_audio_slave;
--synthesis translate_off
    --Audio/avalon_audio_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity CPU_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_debugaccess : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal CPU_instruction_master_latency_counter : IN STD_LOGIC;
                 signal CPU_instruction_master_read : IN STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                 signal CPU_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_data_master_requests_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_instruction_master_granted_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_instruction_master_qualified_request_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_instruction_master_requests_CPU_jtag_debug_module : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal CPU_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_write : OUT STD_LOGIC;
                 signal CPU_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_CPU_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity CPU_jtag_debug_module_arbitrator;


architecture europa of CPU_jtag_debug_module_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_instruction_master_arbiterlock :  STD_LOGIC;
                signal CPU_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_instruction_master_continuerequest :  STD_LOGIC;
                signal CPU_instruction_master_saved_grant_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_jtag_debug_module_allgrants :  STD_LOGIC;
                signal CPU_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal CPU_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal CPU_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal CPU_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal CPU_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal CPU_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal CPU_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal CPU_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal CPU_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal CPU_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal CPU_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal CPU_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal CPU_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal CPU_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal CPU_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal CPU_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal CPU_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_CPU_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_CPU_jtag_debug_module :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_CPU_jtag_debug_module :  STD_LOGIC;
                signal internal_CPU_data_master_requests_CPU_jtag_debug_module :  STD_LOGIC;
                signal internal_CPU_instruction_master_granted_CPU_jtag_debug_module :  STD_LOGIC;
                signal internal_CPU_instruction_master_qualified_request_CPU_jtag_debug_module :  STD_LOGIC;
                signal internal_CPU_instruction_master_requests_CPU_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_CPU_data_master_granted_slave_CPU_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_CPU_instruction_master_granted_slave_CPU_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_CPU_jtag_debug_module_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal shifted_address_to_CPU_jtag_debug_module_from_CPU_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_CPU_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT CPU_jtag_debug_module_end_xfer;
    end if;

  end process;

  CPU_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_CPU_data_master_qualified_request_CPU_jtag_debug_module OR internal_CPU_instruction_master_qualified_request_CPU_jtag_debug_module));
  --assign CPU_jtag_debug_module_readdata_from_sa = CPU_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  CPU_jtag_debug_module_readdata_from_sa <= CPU_jtag_debug_module_readdata;
  internal_CPU_data_master_requests_CPU_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("01010000000000000000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --CPU_jtag_debug_module_arb_share_counter set values, which is an e_mux
  CPU_jtag_debug_module_arb_share_set_values <= std_logic_vector'("001");
  --CPU_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  CPU_jtag_debug_module_non_bursting_master_requests <= ((internal_CPU_data_master_requests_CPU_jtag_debug_module OR internal_CPU_instruction_master_requests_CPU_jtag_debug_module) OR internal_CPU_data_master_requests_CPU_jtag_debug_module) OR internal_CPU_instruction_master_requests_CPU_jtag_debug_module;
  --CPU_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  CPU_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --CPU_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  CPU_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(CPU_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (CPU_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(CPU_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (CPU_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --CPU_jtag_debug_module_allgrants all slave grants, which is an e_mux
  CPU_jtag_debug_module_allgrants <= (((or_reduce(CPU_jtag_debug_module_grant_vector)) OR (or_reduce(CPU_jtag_debug_module_grant_vector))) OR (or_reduce(CPU_jtag_debug_module_grant_vector))) OR (or_reduce(CPU_jtag_debug_module_grant_vector));
  --CPU_jtag_debug_module_end_xfer assignment, which is an e_assign
  CPU_jtag_debug_module_end_xfer <= NOT ((CPU_jtag_debug_module_waits_for_read OR CPU_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_CPU_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_CPU_jtag_debug_module <= CPU_jtag_debug_module_end_xfer AND (((NOT CPU_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --CPU_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  CPU_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_CPU_jtag_debug_module AND CPU_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_CPU_jtag_debug_module AND NOT CPU_jtag_debug_module_non_bursting_master_requests));
  --CPU_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_jtag_debug_module_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(CPU_jtag_debug_module_arb_counter_enable) = '1' then 
        CPU_jtag_debug_module_arb_share_counter <= CPU_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --CPU_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(CPU_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_CPU_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_CPU_jtag_debug_module AND NOT CPU_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        CPU_jtag_debug_module_slavearbiterlockenable <= or_reduce(CPU_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master CPU/jtag_debug_module arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= CPU_jtag_debug_module_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --CPU_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  CPU_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(CPU_jtag_debug_module_arb_share_counter_next_value);
  --CPU/data_master CPU/jtag_debug_module arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= CPU_jtag_debug_module_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --CPU/instruction_master CPU/jtag_debug_module arbiterlock, which is an e_assign
  CPU_instruction_master_arbiterlock <= CPU_jtag_debug_module_slavearbiterlockenable AND CPU_instruction_master_continuerequest;
  --CPU/instruction_master CPU/jtag_debug_module arbiterlock2, which is an e_assign
  CPU_instruction_master_arbiterlock2 <= CPU_jtag_debug_module_slavearbiterlockenable2 AND CPU_instruction_master_continuerequest;
  --CPU/instruction_master granted CPU/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_CPU_instruction_master_granted_slave_CPU_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_CPU_instruction_master_granted_slave_CPU_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(CPU_instruction_master_saved_grant_CPU_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((CPU_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_CPU_instruction_master_requests_CPU_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_CPU_instruction_master_granted_slave_CPU_jtag_debug_module))))));
    end if;

  end process;

  --CPU_instruction_master_continuerequest continued request, which is an e_mux
  CPU_instruction_master_continuerequest <= last_cycle_CPU_instruction_master_granted_slave_CPU_jtag_debug_module AND internal_CPU_instruction_master_requests_CPU_jtag_debug_module;
  --CPU_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  CPU_jtag_debug_module_any_continuerequest <= CPU_instruction_master_continuerequest OR CPU_data_master_continuerequest;
  internal_CPU_data_master_qualified_request_CPU_jtag_debug_module <= internal_CPU_data_master_requests_CPU_jtag_debug_module AND NOT (((((NOT CPU_data_master_waitrequest) AND CPU_data_master_write)) OR CPU_instruction_master_arbiterlock));
  --CPU_jtag_debug_module_writedata mux, which is an e_mux
  CPU_jtag_debug_module_writedata <= CPU_data_master_writedata;
  internal_CPU_instruction_master_requests_CPU_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(CPU_instruction_master_address_to_slave(27 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1010000000000000000000000000")))) AND (CPU_instruction_master_read))) AND CPU_instruction_master_read;
  --CPU/data_master granted CPU/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_CPU_data_master_granted_slave_CPU_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_CPU_data_master_granted_slave_CPU_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(CPU_data_master_saved_grant_CPU_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((CPU_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_CPU_data_master_requests_CPU_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_CPU_data_master_granted_slave_CPU_jtag_debug_module))))));
    end if;

  end process;

  --CPU_data_master_continuerequest continued request, which is an e_mux
  CPU_data_master_continuerequest <= last_cycle_CPU_data_master_granted_slave_CPU_jtag_debug_module AND internal_CPU_data_master_requests_CPU_jtag_debug_module;
  internal_CPU_instruction_master_qualified_request_CPU_jtag_debug_module <= internal_CPU_instruction_master_requests_CPU_jtag_debug_module AND NOT ((((CPU_instruction_master_read AND ((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))) OR (CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register))))) OR CPU_data_master_arbiterlock));
  --local readdatavalid CPU_instruction_master_read_data_valid_CPU_jtag_debug_module, which is an e_mux
  CPU_instruction_master_read_data_valid_CPU_jtag_debug_module <= (internal_CPU_instruction_master_granted_CPU_jtag_debug_module AND CPU_instruction_master_read) AND NOT CPU_jtag_debug_module_waits_for_read;
  --allow new arb cycle for CPU/jtag_debug_module, which is an e_assign
  CPU_jtag_debug_module_allow_new_arb_cycle <= NOT CPU_data_master_arbiterlock AND NOT CPU_instruction_master_arbiterlock;
  --CPU/instruction_master assignment into master qualified-requests vector for CPU/jtag_debug_module, which is an e_assign
  CPU_jtag_debug_module_master_qreq_vector(0) <= internal_CPU_instruction_master_qualified_request_CPU_jtag_debug_module;
  --CPU/instruction_master grant CPU/jtag_debug_module, which is an e_assign
  internal_CPU_instruction_master_granted_CPU_jtag_debug_module <= CPU_jtag_debug_module_grant_vector(0);
  --CPU/instruction_master saved-grant CPU/jtag_debug_module, which is an e_assign
  CPU_instruction_master_saved_grant_CPU_jtag_debug_module <= CPU_jtag_debug_module_arb_winner(0) AND internal_CPU_instruction_master_requests_CPU_jtag_debug_module;
  --CPU/data_master assignment into master qualified-requests vector for CPU/jtag_debug_module, which is an e_assign
  CPU_jtag_debug_module_master_qreq_vector(1) <= internal_CPU_data_master_qualified_request_CPU_jtag_debug_module;
  --CPU/data_master grant CPU/jtag_debug_module, which is an e_assign
  internal_CPU_data_master_granted_CPU_jtag_debug_module <= CPU_jtag_debug_module_grant_vector(1);
  --CPU/data_master saved-grant CPU/jtag_debug_module, which is an e_assign
  CPU_data_master_saved_grant_CPU_jtag_debug_module <= CPU_jtag_debug_module_arb_winner(1) AND internal_CPU_data_master_requests_CPU_jtag_debug_module;
  --CPU/jtag_debug_module chosen-master double-vector, which is an e_assign
  CPU_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((CPU_jtag_debug_module_master_qreq_vector & CPU_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT CPU_jtag_debug_module_master_qreq_vector & NOT CPU_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (CPU_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  CPU_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((CPU_jtag_debug_module_allow_new_arb_cycle AND or_reduce(CPU_jtag_debug_module_grant_vector)))) = '1'), CPU_jtag_debug_module_grant_vector, CPU_jtag_debug_module_saved_chosen_master_vector);
  --saved CPU_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(CPU_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        CPU_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(CPU_jtag_debug_module_grant_vector)) = '1'), CPU_jtag_debug_module_grant_vector, CPU_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  CPU_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((CPU_jtag_debug_module_chosen_master_double_vector(1) OR CPU_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((CPU_jtag_debug_module_chosen_master_double_vector(0) OR CPU_jtag_debug_module_chosen_master_double_vector(2)))));
  --CPU/jtag_debug_module chosen master rotated left, which is an e_assign
  CPU_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(CPU_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(CPU_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --CPU/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(CPU_jtag_debug_module_grant_vector)) = '1' then 
        CPU_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(CPU_jtag_debug_module_end_xfer) = '1'), CPU_jtag_debug_module_chosen_master_rot_left, CPU_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  CPU_jtag_debug_module_begintransfer <= CPU_jtag_debug_module_begins_xfer;
  --assign CPU_jtag_debug_module_resetrequest_from_sa = CPU_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  CPU_jtag_debug_module_resetrequest_from_sa <= CPU_jtag_debug_module_resetrequest;
  CPU_jtag_debug_module_chipselect <= internal_CPU_data_master_granted_CPU_jtag_debug_module OR internal_CPU_instruction_master_granted_CPU_jtag_debug_module;
  --CPU_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  CPU_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(CPU_jtag_debug_module_begins_xfer) = '1'), CPU_jtag_debug_module_unreg_firsttransfer, CPU_jtag_debug_module_reg_firsttransfer);
  --CPU_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  CPU_jtag_debug_module_unreg_firsttransfer <= NOT ((CPU_jtag_debug_module_slavearbiterlockenable AND CPU_jtag_debug_module_any_continuerequest));
  --CPU_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(CPU_jtag_debug_module_begins_xfer) = '1' then 
        CPU_jtag_debug_module_reg_firsttransfer <= CPU_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --CPU_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  CPU_jtag_debug_module_beginbursttransfer_internal <= CPU_jtag_debug_module_begins_xfer;
  --CPU_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  CPU_jtag_debug_module_arbitration_holdoff_internal <= CPU_jtag_debug_module_begins_xfer AND CPU_jtag_debug_module_firsttransfer;
  --CPU_jtag_debug_module_write assignment, which is an e_mux
  CPU_jtag_debug_module_write <= internal_CPU_data_master_granted_CPU_jtag_debug_module AND CPU_data_master_write;
  shifted_address_to_CPU_jtag_debug_module_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --CPU_jtag_debug_module_address mux, which is an e_mux
  CPU_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_CPU_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_CPU_jtag_debug_module_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010"))), (std_logic_vector'("0") & ((A_SRL(shifted_address_to_CPU_jtag_debug_module_from_CPU_instruction_master,std_logic_vector'("00000000000000000000000000000010")))))), 9);
  shifted_address_to_CPU_jtag_debug_module_from_CPU_instruction_master <= CPU_instruction_master_address_to_slave;
  --d1_CPU_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_CPU_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_CPU_jtag_debug_module_end_xfer <= CPU_jtag_debug_module_end_xfer;
    end if;

  end process;

  --CPU_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  CPU_jtag_debug_module_waits_for_read <= CPU_jtag_debug_module_in_a_read_cycle AND CPU_jtag_debug_module_begins_xfer;
  --CPU_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  CPU_jtag_debug_module_in_a_read_cycle <= ((internal_CPU_data_master_granted_CPU_jtag_debug_module AND CPU_data_master_read)) OR ((internal_CPU_instruction_master_granted_CPU_jtag_debug_module AND CPU_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= CPU_jtag_debug_module_in_a_read_cycle;
  --CPU_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  CPU_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --CPU_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  CPU_jtag_debug_module_in_a_write_cycle <= internal_CPU_data_master_granted_CPU_jtag_debug_module AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= CPU_jtag_debug_module_in_a_write_cycle;
  wait_for_CPU_jtag_debug_module_counter <= std_logic'('0');
  --CPU_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  CPU_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_CPU_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  CPU_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_CPU_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  CPU_data_master_granted_CPU_jtag_debug_module <= internal_CPU_data_master_granted_CPU_jtag_debug_module;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_CPU_jtag_debug_module <= internal_CPU_data_master_qualified_request_CPU_jtag_debug_module;
  --vhdl renameroo for output signals
  CPU_data_master_requests_CPU_jtag_debug_module <= internal_CPU_data_master_requests_CPU_jtag_debug_module;
  --vhdl renameroo for output signals
  CPU_instruction_master_granted_CPU_jtag_debug_module <= internal_CPU_instruction_master_granted_CPU_jtag_debug_module;
  --vhdl renameroo for output signals
  CPU_instruction_master_qualified_request_CPU_jtag_debug_module <= internal_CPU_instruction_master_qualified_request_CPU_jtag_debug_module;
  --vhdl renameroo for output signals
  CPU_instruction_master_requests_CPU_jtag_debug_module <= internal_CPU_instruction_master_requests_CPU_jtag_debug_module;
--synthesis translate_off
    --CPU/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_granted_CPU_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_CPU_instruction_master_granted_CPU_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(CPU_data_master_saved_grant_CPU_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_saved_grant_CPU_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity CPU_custom_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal CPU_custom_instruction_master_multi_start : IN STD_LOGIC;
                 signal CPU_fpoint_s1_done_from_sa : IN STD_LOGIC;
                 signal CPU_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_custom_instruction_master_multi_done : OUT STD_LOGIC;
                 signal CPU_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_custom_instruction_master_reset_n : OUT STD_LOGIC;
                 signal CPU_custom_instruction_master_start_CPU_fpoint_s1 : OUT STD_LOGIC;
                 signal CPU_fpoint_s1_select : OUT STD_LOGIC
              );
end entity CPU_custom_instruction_master_arbitrator;


architecture europa of CPU_custom_instruction_master_arbitrator is
                signal internal_CPU_fpoint_s1_select :  STD_LOGIC;

begin

  internal_CPU_fpoint_s1_select <= std_logic'('1');
  CPU_custom_instruction_master_start_CPU_fpoint_s1 <= internal_CPU_fpoint_s1_select AND CPU_custom_instruction_master_multi_start;
  --CPU_custom_instruction_master_multi_result mux, which is an e_mux
  CPU_custom_instruction_master_multi_result <= A_REP(internal_CPU_fpoint_s1_select, 32) AND CPU_fpoint_s1_result_from_sa;
  --multi_done mux, which is an e_mux
  CPU_custom_instruction_master_multi_done <= internal_CPU_fpoint_s1_select AND CPU_fpoint_s1_done_from_sa;
  --CPU_custom_instruction_master_reset_n local reset_n, which is an e_assign
  CPU_custom_instruction_master_reset_n <= reset_n;
  --vhdl renameroo for output signals
  CPU_fpoint_s1_select <= internal_CPU_fpoint_s1_select;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity CPU_data_master_arbitrator is 
        port (
              -- inputs:
                 signal AV_Config_avalon_av_config_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal AV_Config_avalon_av_config_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal Audio_avalon_audio_slave_irq_from_sa : IN STD_LOGIC;
                 signal Audio_avalon_audio_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_address : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                 signal CPU_data_master_byteenable_SDRAM_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_byteenable_SRAM_avalon_sram_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal CPU_data_master_byteenable_nios_system_clock_0_in : IN STD_LOGIC;
                 signal CPU_data_master_granted_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Audio_avalon_audio_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Interval_Timer_s1 : IN STD_LOGIC;
                 signal CPU_data_master_granted_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_data_master_granted_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_granted_nios_system_clock_0_in : IN STD_LOGIC;
                 signal CPU_data_master_granted_sysid_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Audio_avalon_audio_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Interval_Timer_s1 : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_nios_system_clock_0_in : IN STD_LOGIC;
                 signal CPU_data_master_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Interval_Timer_s1 : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_nios_system_clock_0_in : IN STD_LOGIC;
                 signal CPU_data_master_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Audio_avalon_audio_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Interval_Timer_s1 : IN STD_LOGIC;
                 signal CPU_data_master_requests_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_data_master_requests_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_requests_nios_system_clock_0_in : IN STD_LOGIC;
                 signal CPU_data_master_requests_sysid_control_slave : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Expansion_JP2_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Green_LEDs_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Interval_Timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal Interval_Timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal JTAG_UART_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal JTAG_UART_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_irq_from_sa : IN STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal PS2_Port_avalon_ps2_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Red_LEDs_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal SDRAM_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SDRAM_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal SRAM_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal Serial_Port_avalon_rs232_slave_irq_from_sa : IN STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Slider_Switches_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_AV_Config_avalon_av_config_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Audio_avalon_audio_slave_end_xfer : IN STD_LOGIC;
                 signal d1_CPU_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Green_LEDs_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Interval_Timer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_JTAG_UART_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_PS2_Port_avalon_ps2_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Pushbuttons_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Red_LEDs_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_SDRAM_s1_end_xfer : IN STD_LOGIC;
                 signal d1_SRAM_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Serial_Port_avalon_rs232_slave_end_xfer : IN STD_LOGIC;
                 signal d1_Slider_Switches_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                 signal d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer : IN STD_LOGIC;
                 signal d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_nios_system_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal nios_system_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios_system_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal CPU_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal CPU_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal CPU_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                 signal CPU_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_data_master_waitrequest : OUT STD_LOGIC
              );
end entity CPU_data_master_arbitrator;


architecture europa of CPU_data_master_arbitrator is
                signal CPU_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_run :  STD_LOGIC;
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_CPU_data_master_address_to_slave :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal internal_CPU_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_CPU_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal internal_CPU_data_master_waitrequest :  STD_LOGIC;
                signal last_dbs_term_and_run :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_dbs_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_registered_CPU_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;
                signal r_4 :  STD_LOGIC;
                signal registered_CPU_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave OR registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave) OR NOT CPU_data_master_requests_AV_Config_avalon_av_config_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT AV_Config_avalon_av_config_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Audio_avalon_audio_slave OR registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave) OR NOT CPU_data_master_requests_Audio_avalon_audio_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Audio_avalon_audio_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Audio_avalon_audio_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_qualified_request_CPU_jtag_debug_module OR NOT CPU_data_master_requests_CPU_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_granted_CPU_jtag_debug_module OR NOT CPU_data_master_qualified_request_CPU_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_CPU_jtag_debug_module OR NOT CPU_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_CPU_jtag_debug_module OR NOT CPU_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave OR ((((CPU_data_master_write AND NOT(CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave)) AND internal_CPU_data_master_dbs_address(1)) AND internal_CPU_data_master_dbs_address(0)))) OR NOT CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave OR NOT CPU_data_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave OR NOT CPU_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  CPU_data_master_run <= (((r_0 AND r_1) AND r_2) AND r_3) AND r_4;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_qualified_request_Interval_Timer_s1 OR NOT CPU_data_master_requests_Interval_Timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Interval_Timer_s1 OR NOT CPU_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read)))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Interval_Timer_s1 OR NOT CPU_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave OR NOT CPU_data_master_requests_JTAG_UART_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT JTAG_UART_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT JTAG_UART_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave OR registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave) OR NOT CPU_data_master_requests_PS2_Port_avalon_ps2_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT PS2_Port_avalon_ps2_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((CPU_data_master_qualified_request_SDRAM_s1 OR ((CPU_data_master_read_data_valid_SDRAM_s1 AND internal_CPU_data_master_dbs_address(1)))) OR (((CPU_data_master_write AND NOT(or_reduce(CPU_data_master_byteenable_SDRAM_s1))) AND internal_CPU_data_master_dbs_address(1)))) OR NOT CPU_data_master_requests_SDRAM_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_granted_SDRAM_s1 OR NOT CPU_data_master_qualified_request_SDRAM_s1)))))));
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_SDRAM_s1 OR NOT CPU_data_master_read) OR (((CPU_data_master_read_data_valid_SDRAM_s1 AND (internal_CPU_data_master_dbs_address(1))) AND CPU_data_master_read))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_SDRAM_s1 OR NOT CPU_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT SDRAM_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_CPU_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((CPU_data_master_qualified_request_SRAM_avalon_sram_slave OR ((CPU_data_master_read_data_valid_SRAM_avalon_sram_slave AND internal_CPU_data_master_dbs_address(1)))) OR (((CPU_data_master_write AND NOT(or_reduce(CPU_data_master_byteenable_SRAM_avalon_sram_slave))) AND internal_CPU_data_master_dbs_address(1)))) OR NOT CPU_data_master_requests_SRAM_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_granted_SRAM_avalon_sram_slave OR NOT CPU_data_master_qualified_request_SRAM_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_SRAM_avalon_sram_slave OR NOT CPU_data_master_read) OR (((CPU_data_master_read_data_valid_SRAM_avalon_sram_slave AND (internal_CPU_data_master_dbs_address(1))) AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_SRAM_avalon_sram_slave OR NOT CPU_data_master_write)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_CPU_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave OR registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave) OR NOT CPU_data_master_requests_Serial_Port_avalon_rs232_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave OR registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave) OR NOT CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave OR (((registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave AND internal_CPU_data_master_dbs_address(1)) AND internal_CPU_data_master_dbs_address(0)))) OR ((((CPU_data_master_write AND NOT(CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave)) AND internal_CPU_data_master_dbs_address(1)) AND internal_CPU_data_master_dbs_address(0)))) OR NOT CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave OR NOT CPU_data_master_read) OR (((registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave AND ((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0)))) AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave OR NOT CPU_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --r_4 master_run cascaded wait assignment, which is an e_assign
  r_4 <= Vector_To_Std_Logic((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave OR registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave) OR NOT CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave)) AND (((NOT CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave OR registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave) OR NOT CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave OR NOT CPU_data_master_read) OR ((registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave OR NOT ((CPU_data_master_read OR CPU_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_read OR CPU_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((CPU_data_master_qualified_request_nios_system_clock_0_in OR ((((CPU_data_master_write AND NOT(CPU_data_master_byteenable_nios_system_clock_0_in)) AND internal_CPU_data_master_dbs_address(1)) AND internal_CPU_data_master_dbs_address(0)))) OR NOT CPU_data_master_requests_nios_system_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_nios_system_clock_0_in OR NOT CPU_data_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios_system_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_nios_system_clock_0_in OR NOT CPU_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios_system_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_CPU_data_master_dbs_address(1) AND internal_CPU_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_sysid_control_slave OR NOT CPU_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_data_master_qualified_request_sysid_control_slave OR NOT CPU_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_CPU_data_master_address_to_slave <= Std_Logic_Vector'(CPU_data_master_address(28 DOWNTO 27) & A_ToStdLogicVector(std_logic'('0')) & CPU_data_master_address(25 DOWNTO 24) & A_ToStdLogicVector(std_logic'('0')) & CPU_data_master_address(22 DOWNTO 0));
  --CPU/data_master readdata mux, which is an e_mux
  CPU_data_master_readdata <= (((((((((((((((((((((((A_REP(NOT CPU_data_master_requests_AV_Config_avalon_av_config_slave, 32) OR AV_Config_avalon_av_config_slave_readdata_from_sa)) AND ((A_REP(NOT CPU_data_master_requests_Audio_avalon_audio_slave, 32) OR Audio_avalon_audio_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_CPU_jtag_debug_module, 32) OR CPU_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave, 32) OR registered_CPU_data_master_readdata))) AND ((A_REP(NOT CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave, 32) OR Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave, 32) OR Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave, 32) OR Green_LEDs_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave, 32) OR HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave, 32) OR HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Interval_Timer_s1, 32) OR (std_logic_vector'("0000000000000000") & (Interval_Timer_s1_readdata_from_sa))))) AND ((A_REP(NOT CPU_data_master_requests_JTAG_UART_avalon_jtag_slave, 32) OR registered_CPU_data_master_readdata))) AND ((A_REP(NOT CPU_data_master_requests_PS2_Port_avalon_ps2_slave, 32) OR PS2_Port_avalon_ps2_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave, 32) OR Pushbuttons_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave, 32) OR Red_LEDs_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_SDRAM_s1, 32) OR registered_CPU_data_master_readdata))) AND ((A_REP(NOT CPU_data_master_requests_SRAM_avalon_sram_slave, 32) OR registered_CPU_data_master_readdata))) AND ((A_REP(NOT CPU_data_master_requests_Serial_Port_avalon_rs232_slave, 32) OR Serial_Port_avalon_rs232_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave, 32) OR Slider_Switches_avalon_parallel_port_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave, 32) OR Std_Logic_Vector'(VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa(7 DOWNTO 0) & dbs_8_reg_segment_2 & dbs_8_reg_segment_1 & dbs_8_reg_segment_0)))) AND ((A_REP(NOT CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave, 32) OR VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave, 32) OR VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_nios_system_clock_0_in, 32) OR registered_CPU_data_master_readdata))) AND ((A_REP(NOT CPU_data_master_requests_sysid_control_slave, 32) OR sysid_control_slave_readdata_from_sa));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_CPU_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_CPU_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((CPU_data_master_read OR CPU_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_data_master_run AND internal_CPU_data_master_waitrequest))))))));
    end if;

  end process;

  --irq assign, which is an e_assign
  CPU_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(Expansion_JP2_avalon_parallel_port_slave_irq_from_sa) & A_ToStdLogicVector(Expansion_JP1_avalon_parallel_port_slave_irq_from_sa) & A_ToStdLogicVector(Serial_Port_avalon_rs232_slave_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(JTAG_UART_avalon_jtag_slave_irq_from_sa) & A_ToStdLogicVector(PS2_Port_avalon_ps2_slave_irq_from_sa) & A_ToStdLogicVector(Audio_avalon_audio_slave_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(Pushbuttons_avalon_parallel_port_slave_irq_from_sa) & A_ToStdLogicVector(Interval_Timer_s1_irq_from_sa));
  --no_byte_enables_and_last_term, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_CPU_data_master_no_byte_enables_and_last_term <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_CPU_data_master_no_byte_enables_and_last_term <= last_dbs_term_and_run;
    end if;

  end process;

  --compute the last dbs term, which is an e_mux
  last_dbs_term_and_run <= A_WE_StdLogic((std_logic'((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)) = '1'), (((to_std_logic(((internal_CPU_data_master_dbs_address = std_logic_vector'("11")))) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave))), A_WE_StdLogic((std_logic'((CPU_data_master_requests_SDRAM_s1)) = '1'), (((to_std_logic(((internal_CPU_data_master_dbs_address = std_logic_vector'("10")))) AND CPU_data_master_write) AND NOT(or_reduce(CPU_data_master_byteenable_SDRAM_s1)))), A_WE_StdLogic((std_logic'((CPU_data_master_requests_SRAM_avalon_sram_slave)) = '1'), (((to_std_logic(((internal_CPU_data_master_dbs_address = std_logic_vector'("10")))) AND CPU_data_master_write) AND NOT(or_reduce(CPU_data_master_byteenable_SRAM_avalon_sram_slave)))), A_WE_StdLogic((std_logic'((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), (((to_std_logic(((internal_CPU_data_master_dbs_address = std_logic_vector'("11")))) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave))), (((to_std_logic(((internal_CPU_data_master_dbs_address = std_logic_vector'("11")))) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_nios_system_clock_0_in)))))));
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_CPU_data_master_no_byte_enables_and_last_term) AND CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_CPU_data_master_no_byte_enables_and_last_term) AND CPU_data_master_requests_SDRAM_s1) AND CPU_data_master_write) AND NOT(or_reduce(CPU_data_master_byteenable_SDRAM_s1)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read_data_valid_SDRAM_s1)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_SDRAM_s1 AND CPU_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT SDRAM_s1_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_CPU_data_master_no_byte_enables_and_last_term) AND CPU_data_master_requests_SRAM_avalon_sram_slave) AND CPU_data_master_write) AND NOT(or_reduce(CPU_data_master_byteenable_SRAM_avalon_sram_slave)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read_data_valid_SRAM_avalon_sram_slave)))) OR ((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_SRAM_avalon_sram_slave AND CPU_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_CPU_data_master_no_byte_enables_and_last_term) AND CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_CPU_data_master_no_byte_enables_and_last_term) AND CPU_data_master_requests_nios_system_clock_0_in) AND CPU_data_master_write) AND NOT(CPU_data_master_byteenable_nios_system_clock_0_in))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios_system_clock_0_in_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios_system_clock_0_in_waitrequest_from_sa)))))));
  --input to dbs-8 stored 0, which is an e_mux
  p1_dbs_8_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)) = '1'), Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa, A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa, nios_system_clock_0_in_readdata_from_sa));
  --dbs register for dbs-8 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_0 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_CPU_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
      end if;
    end if;

  end process;

  --input to dbs-8 stored 1, which is an e_mux
  p1_dbs_8_reg_segment_1 <= A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)) = '1'), Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa, A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa, nios_system_clock_0_in_readdata_from_sa));
  --dbs register for dbs-8 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_1 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_CPU_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
      end if;
    end if;

  end process;

  --input to dbs-8 stored 2, which is an e_mux
  p1_dbs_8_reg_segment_2 <= A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)) = '1'), Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa, A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa, nios_system_clock_0_in_readdata_from_sa));
  --dbs register for dbs-8 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_2 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_CPU_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
      end if;
    end if;

  end process;

  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_CPU_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_CPU_data_master_readdata <= p1_registered_CPU_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_CPU_data_master_readdata <= (((((A_REP(NOT CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave, 32) OR Std_Logic_Vector'(Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa(7 DOWNTO 0) & dbs_8_reg_segment_2 & dbs_8_reg_segment_1 & dbs_8_reg_segment_0))) AND ((A_REP(NOT CPU_data_master_requests_JTAG_UART_avalon_jtag_slave, 32) OR JTAG_UART_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT CPU_data_master_requests_SDRAM_s1, 32) OR Std_Logic_Vector'(SDRAM_s1_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)))) AND ((A_REP(NOT CPU_data_master_requests_SRAM_avalon_sram_slave, 32) OR Std_Logic_Vector'(SRAM_avalon_sram_slave_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)))) AND ((A_REP(NOT CPU_data_master_requests_nios_system_clock_0_in, 32) OR Std_Logic_Vector'(nios_system_clock_0_in_readdata_from_sa(7 DOWNTO 0) & dbs_8_reg_segment_2 & dbs_8_reg_segment_1 & dbs_8_reg_segment_0)));
  --mux write dbs 2, which is an e_mux
  CPU_data_master_dbs_write_8 <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_writedata(23 DOWNTO 16), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000011"))), CPU_data_master_writedata(31 DOWNTO 24), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_writedata(23 DOWNTO 16), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000011"))), CPU_data_master_writedata(31 DOWNTO 24), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_writedata(23 DOWNTO 16), CPU_data_master_writedata(31 DOWNTO 24))))))))))));
  --dbs count increment, which is an e_mux
  CPU_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_SRAM_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_nios_system_clock_0_in)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000")))))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_CPU_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_CPU_data_master_dbs_address)) + (std_logic_vector'("0") & (CPU_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= ((((pre_dbs_count_enable AND (NOT ((CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave AND NOT internal_CPU_data_master_waitrequest)))) AND (NOT ((CPU_data_master_requests_SDRAM_s1 AND NOT internal_CPU_data_master_waitrequest)))) AND (NOT ((CPU_data_master_requests_SRAM_avalon_sram_slave AND NOT internal_CPU_data_master_waitrequest)))) AND (NOT (((CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave AND NOT internal_CPU_data_master_waitrequest) AND CPU_data_master_write)))) AND (NOT ((CPU_data_master_requests_nios_system_clock_0_in AND NOT internal_CPU_data_master_waitrequest)));
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_CPU_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_CPU_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((CPU_data_master_requests_SDRAM_s1)) = '1'), SDRAM_s1_readdata_from_sa, SRAM_avalon_sram_slave_readdata_from_sa);
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_CPU_data_master_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  CPU_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_dbs_address(1))) = '1'), CPU_data_master_writedata(31 DOWNTO 16), A_WE_StdLogicVector((std_logic'((NOT (internal_CPU_data_master_dbs_address(1)))) = '1'), CPU_data_master_writedata(15 DOWNTO 0), A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_dbs_address(1))) = '1'), CPU_data_master_writedata(31 DOWNTO 16), CPU_data_master_writedata(15 DOWNTO 0))));
  --vhdl renameroo for output signals
  CPU_data_master_address_to_slave <= internal_CPU_data_master_address_to_slave;
  --vhdl renameroo for output signals
  CPU_data_master_dbs_address <= internal_CPU_data_master_dbs_address;
  --vhdl renameroo for output signals
  CPU_data_master_no_byte_enables_and_last_term <= internal_CPU_data_master_no_byte_enables_and_last_term;
  --vhdl renameroo for output signals
  CPU_data_master_waitrequest <= internal_CPU_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity CPU_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal CPU_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal CPU_instruction_master_granted_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_instruction_master_granted_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_instruction_master_qualified_request_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_instruction_master_qualified_request_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_instruction_master_read : IN STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                 signal CPU_instruction_master_requests_CPU_jtag_debug_module : IN STD_LOGIC;
                 signal CPU_instruction_master_requests_SDRAM_s1 : IN STD_LOGIC;
                 signal CPU_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal SDRAM_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SDRAM_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal d1_CPU_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_SDRAM_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal CPU_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_instruction_master_latency_counter : OUT STD_LOGIC;
                 signal CPU_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal CPU_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity CPU_instruction_master_arbitrator;


architecture europa of CPU_instruction_master_arbitrator is
                signal CPU_instruction_master_address_last_time :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal CPU_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_instruction_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_instruction_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal CPU_instruction_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal CPU_instruction_master_read_last_time :  STD_LOGIC;
                signal CPU_instruction_master_run :  STD_LOGIC;
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_CPU_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_CPU_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_CPU_instruction_master_latency_counter :  STD_LOGIC;
                signal internal_CPU_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_CPU_instruction_master_latency_counter :  STD_LOGIC;
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_CPU_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_instruction_master_qualified_request_CPU_jtag_debug_module OR NOT CPU_instruction_master_requests_CPU_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_instruction_master_granted_CPU_jtag_debug_module OR NOT CPU_instruction_master_qualified_request_CPU_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_instruction_master_qualified_request_CPU_jtag_debug_module OR NOT CPU_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_CPU_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  CPU_instruction_master_run <= (r_0 AND r_2) AND r_3;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_instruction_master_qualified_request_SDRAM_s1 OR NOT CPU_instruction_master_requests_SDRAM_s1)))))));
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((CPU_instruction_master_granted_SDRAM_s1 OR NOT CPU_instruction_master_qualified_request_SDRAM_s1))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT CPU_instruction_master_qualified_request_SDRAM_s1 OR NOT CPU_instruction_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT SDRAM_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_CPU_instruction_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_CPU_instruction_master_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(CPU_instruction_master_address(27)) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(CPU_instruction_master_address(25)) & std_logic_vector'("00") & CPU_instruction_master_address(22 DOWNTO 0));
  --CPU_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_instruction_master_read_but_no_slave_selected <= (CPU_instruction_master_read AND CPU_instruction_master_run) AND NOT CPU_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  CPU_instruction_master_is_granted_some_slave <= CPU_instruction_master_granted_CPU_jtag_debug_module OR CPU_instruction_master_granted_SDRAM_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_CPU_instruction_master_readdatavalid <= CPU_instruction_master_read_data_valid_SDRAM_s1 AND dbs_rdv_counter_overflow;
  --latent slave read data valid which is not flushed, which is an e_mux
  CPU_instruction_master_readdatavalid <= (((CPU_instruction_master_read_but_no_slave_selected OR pre_flush_CPU_instruction_master_readdatavalid) OR CPU_instruction_master_read_data_valid_CPU_jtag_debug_module) OR CPU_instruction_master_read_but_no_slave_selected) OR pre_flush_CPU_instruction_master_readdatavalid;
  --CPU/instruction_master readdata mux, which is an e_mux
  CPU_instruction_master_readdata <= ((A_REP(NOT ((CPU_instruction_master_qualified_request_CPU_jtag_debug_module AND CPU_instruction_master_read)) , 32) OR CPU_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT CPU_instruction_master_read_data_valid_SDRAM_s1, 32) OR Std_Logic_Vector'(SDRAM_s1_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_CPU_instruction_master_waitrequest <= NOT CPU_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_CPU_instruction_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_CPU_instruction_master_latency_counter <= p1_CPU_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_CPU_instruction_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((CPU_instruction_master_run AND CPU_instruction_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_CPU_instruction_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_CPU_instruction_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= SDRAM_s1_readdata_from_sa;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_instruction_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  CPU_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((CPU_instruction_master_requests_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_CPU_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_CPU_instruction_master_dbs_address)) + (std_logic_vector'("0") & (CPU_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_CPU_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_CPU_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  CPU_instruction_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (CPU_instruction_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (CPU_instruction_master_dbs_rdv_counter_inc))), 2);
  --CPU_instruction_master_rdv_inc_mux, which is an e_mux
  CPU_instruction_master_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= CPU_instruction_master_read_data_valid_SDRAM_s1;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_instruction_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        CPU_instruction_master_dbs_rdv_counter <= CPU_instruction_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= CPU_instruction_master_dbs_rdv_counter(1) AND NOT CPU_instruction_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((CPU_instruction_master_granted_SDRAM_s1 AND CPU_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT SDRAM_s1_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  CPU_instruction_master_address_to_slave <= internal_CPU_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  CPU_instruction_master_dbs_address <= internal_CPU_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  CPU_instruction_master_latency_counter <= internal_CPU_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  CPU_instruction_master_waitrequest <= internal_CPU_instruction_master_waitrequest;
--synthesis translate_off
    --CPU_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        CPU_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000000");
      elsif clk'event and clk = '1' then
        CPU_instruction_master_address_last_time <= CPU_instruction_master_address;
      end if;

    end process;

    --CPU/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_CPU_instruction_master_waitrequest AND (CPU_instruction_master_read);
      end if;

    end process;

    --CPU_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((CPU_instruction_master_address /= CPU_instruction_master_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("CPU_instruction_master_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --CPU_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        CPU_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        CPU_instruction_master_read_last_time <= CPU_instruction_master_read;
      end if;

    end process;

    --CPU_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(CPU_instruction_master_read) /= std_logic'(CPU_instruction_master_read_last_time)))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("CPU_instruction_master_read did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity CPU_fpoint_s1_arbitrator is 
        port (
              -- inputs:
                 signal CPU_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                 signal CPU_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal CPU_custom_instruction_master_start_CPU_fpoint_s1 : IN STD_LOGIC;
                 signal CPU_fpoint_s1_done : IN STD_LOGIC;
                 signal CPU_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_fpoint_s1_select : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_fpoint_s1_clk_en : OUT STD_LOGIC;
                 signal CPU_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                 signal CPU_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_fpoint_s1_reset : OUT STD_LOGIC;
                 signal CPU_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal CPU_fpoint_s1_start : OUT STD_LOGIC
              );
end entity CPU_fpoint_s1_arbitrator;


architecture europa of CPU_fpoint_s1_arbitrator is

begin

  CPU_fpoint_s1_clk_en <= CPU_custom_instruction_master_multi_clk_en;
  CPU_fpoint_s1_dataa <= CPU_custom_instruction_master_multi_dataa;
  CPU_fpoint_s1_datab <= CPU_custom_instruction_master_multi_datab;
  CPU_fpoint_s1_n <= CPU_custom_instruction_master_multi_n (1 DOWNTO 0);
  CPU_fpoint_s1_start <= CPU_custom_instruction_master_start_CPU_fpoint_s1;
  --assign CPU_fpoint_s1_result_from_sa = CPU_fpoint_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  CPU_fpoint_s1_result_from_sa <= CPU_fpoint_s1_result;
  --assign CPU_fpoint_s1_done_from_sa = CPU_fpoint_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  CPU_fpoint_s1_done_from_sa <= CPU_fpoint_s1_done;
  --CPU_fpoint/s1 local reset_n, which is an e_assign
  CPU_fpoint_s1_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Char_LCD_16x2_avalon_lcd_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal Char_LCD_16x2_avalon_lcd_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                 signal CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_address : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_chipselect : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_read : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal Char_LCD_16x2_avalon_lcd_slave_reset : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_write : OUT STD_LOGIC;
                 signal Char_LCD_16x2_avalon_lcd_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer : OUT STD_LOGIC
              );
end entity Char_LCD_16x2_avalon_lcd_slave_arbitrator;


architecture europa of Char_LCD_16x2_avalon_lcd_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_0 :  STD_LOGIC;
                signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_1 :  STD_LOGIC;
                signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_3 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_allgrants :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_any_continuerequest :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_arb_counter_enable :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_begins_xfer :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_end_xfer :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_firsttransfer :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_grant_vector :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_in_a_read_cycle :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_in_a_write_cycle :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_master_qreq_vector :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_pretend_byte_enable :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_reg_firsttransfer :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_waits_for_read :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal internal_Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa :  STD_LOGIC;
                signal wait_for_Char_LCD_16x2_avalon_lcd_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Char_LCD_16x2_avalon_lcd_slave_end_xfer;
    end if;

  end process;

  Char_LCD_16x2_avalon_lcd_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave);
  --assign Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa = Char_LCD_16x2_avalon_lcd_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa <= Char_LCD_16x2_avalon_lcd_slave_readdata;
  internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 1) & A_ToStdLogicVector(std_logic'('0'))) = std_logic_vector'("10000000000000011000001010000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa = Char_LCD_16x2_avalon_lcd_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa <= Char_LCD_16x2_avalon_lcd_slave_waitrequest;
  --Char_LCD_16x2_avalon_lcd_slave_arb_share_counter set values, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000001")), 3);
  --Char_LCD_16x2_avalon_lcd_slave_non_bursting_master_requests mux, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave;
  --Char_LCD_16x2_avalon_lcd_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value assignment, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Char_LCD_16x2_avalon_lcd_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Char_LCD_16x2_avalon_lcd_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Char_LCD_16x2_avalon_lcd_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Char_LCD_16x2_avalon_lcd_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Char_LCD_16x2_avalon_lcd_slave_allgrants all slave grants, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_allgrants <= Char_LCD_16x2_avalon_lcd_slave_grant_vector;
  --Char_LCD_16x2_avalon_lcd_slave_end_xfer assignment, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_end_xfer <= NOT ((Char_LCD_16x2_avalon_lcd_slave_waits_for_read OR Char_LCD_16x2_avalon_lcd_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave <= Char_LCD_16x2_avalon_lcd_slave_end_xfer AND (((NOT Char_LCD_16x2_avalon_lcd_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Char_LCD_16x2_avalon_lcd_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave AND Char_LCD_16x2_avalon_lcd_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave AND NOT Char_LCD_16x2_avalon_lcd_slave_non_bursting_master_requests));
  --Char_LCD_16x2_avalon_lcd_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Char_LCD_16x2_avalon_lcd_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Char_LCD_16x2_avalon_lcd_slave_arb_counter_enable) = '1' then 
        Char_LCD_16x2_avalon_lcd_slave_arb_share_counter <= Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Char_LCD_16x2_avalon_lcd_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave)) OR ((end_xfer_arb_share_counter_term_Char_LCD_16x2_avalon_lcd_slave AND NOT Char_LCD_16x2_avalon_lcd_slave_non_bursting_master_requests)))) = '1' then 
        Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable <= or_reduce(Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Char_LCD_16x2/avalon_lcd_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable2 <= or_reduce(Char_LCD_16x2_avalon_lcd_slave_arb_share_counter_next_value);
  --CPU/data_master Char_LCD_16x2/avalon_lcd_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Char_LCD_16x2_avalon_lcd_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave AND NOT ((((CPU_data_master_read AND (NOT CPU_data_master_waitrequest))) OR (((((NOT CPU_data_master_waitrequest OR CPU_data_master_no_byte_enables_and_last_term) OR NOT(internal_CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave))) AND CPU_data_master_write))));
  --Char_LCD_16x2_avalon_lcd_slave_writedata mux, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_writedata <= CPU_data_master_dbs_write_8;
  --master is always granted when requested
  internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave;
  --CPU/data_master saved-grant Char_LCD_16x2/avalon_lcd_slave, which is an e_assign
  CPU_data_master_saved_grant_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave;
  --allow new arb cycle for Char_LCD_16x2/avalon_lcd_slave, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Char_LCD_16x2_avalon_lcd_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Char_LCD_16x2_avalon_lcd_slave_master_qreq_vector <= std_logic'('1');
  --~Char_LCD_16x2_avalon_lcd_slave_reset assignment, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_reset <= NOT reset_n;
  Char_LCD_16x2_avalon_lcd_slave_chipselect <= internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave;
  --Char_LCD_16x2_avalon_lcd_slave_firsttransfer first transaction, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Char_LCD_16x2_avalon_lcd_slave_begins_xfer) = '1'), Char_LCD_16x2_avalon_lcd_slave_unreg_firsttransfer, Char_LCD_16x2_avalon_lcd_slave_reg_firsttransfer);
  --Char_LCD_16x2_avalon_lcd_slave_unreg_firsttransfer first transaction, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_unreg_firsttransfer <= NOT ((Char_LCD_16x2_avalon_lcd_slave_slavearbiterlockenable AND Char_LCD_16x2_avalon_lcd_slave_any_continuerequest));
  --Char_LCD_16x2_avalon_lcd_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Char_LCD_16x2_avalon_lcd_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Char_LCD_16x2_avalon_lcd_slave_begins_xfer) = '1' then 
        Char_LCD_16x2_avalon_lcd_slave_reg_firsttransfer <= Char_LCD_16x2_avalon_lcd_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Char_LCD_16x2_avalon_lcd_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_beginbursttransfer_internal <= Char_LCD_16x2_avalon_lcd_slave_begins_xfer;
  --Char_LCD_16x2_avalon_lcd_slave_read assignment, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_read <= internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_read;
  --Char_LCD_16x2_avalon_lcd_slave_write assignment, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_write <= ((internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_write)) AND Char_LCD_16x2_avalon_lcd_slave_pretend_byte_enable;
  --Char_LCD_16x2_avalon_lcd_slave_address mux, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_address <= Vector_To_Std_Logic(Std_Logic_Vector'(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & CPU_data_master_dbs_address(1 DOWNTO 0)));
  --d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer <= Char_LCD_16x2_avalon_lcd_slave_end_xfer;
    end if;

  end process;

  --Char_LCD_16x2_avalon_lcd_slave_waits_for_read in a cycle, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_waits_for_read <= Char_LCD_16x2_avalon_lcd_slave_in_a_read_cycle AND internal_Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa;
  --Char_LCD_16x2_avalon_lcd_slave_in_a_read_cycle assignment, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Char_LCD_16x2_avalon_lcd_slave_in_a_read_cycle;
  --Char_LCD_16x2_avalon_lcd_slave_waits_for_write in a cycle, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_waits_for_write <= Char_LCD_16x2_avalon_lcd_slave_in_a_write_cycle AND internal_Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa;
  --Char_LCD_16x2_avalon_lcd_slave_in_a_write_cycle assignment, which is an e_assign
  Char_LCD_16x2_avalon_lcd_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Char_LCD_16x2_avalon_lcd_slave_in_a_write_cycle;
  wait_for_Char_LCD_16x2_avalon_lcd_slave_counter <= std_logic'('0');
  --Char_LCD_16x2_avalon_lcd_slave_pretend_byte_enable byte enable port mux, which is an e_mux
  Char_LCD_16x2_avalon_lcd_slave_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_3, CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_2, CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_1, CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_0) <= CPU_data_master_byteenable;
  internal_CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_2, CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave_segment_3)));
  --vhdl renameroo for output signals
  CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave <= internal_CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave;
  --vhdl renameroo for output signals
  Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa <= internal_Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa;
--synthesis translate_off
    --Char_LCD_16x2/avalon_lcd_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Expansion_JP1_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Expansion_JP1_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Expansion_JP1_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Expansion_JP1_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Expansion_JP1_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Expansion_JP1_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Expansion_JP1_avalon_parallel_port_slave_arbitrator;


architecture europa of Expansion_JP1_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Expansion_JP1_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Expansion_JP1_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Expansion_JP1_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Expansion_JP1_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave);
  --assign Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa = Expansion_JP1_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa <= Expansion_JP1_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000001100000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register_in;
  --Expansion_JP1_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Expansion_JP1_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave;
  --Expansion_JP1_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Expansion_JP1_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Expansion_JP1_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Expansion_JP1_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Expansion_JP1_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Expansion_JP1_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_allgrants <= Expansion_JP1_avalon_parallel_port_slave_grant_vector;
  --Expansion_JP1_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_end_xfer <= NOT ((Expansion_JP1_avalon_parallel_port_slave_waits_for_read OR Expansion_JP1_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave <= Expansion_JP1_avalon_parallel_port_slave_end_xfer AND (((NOT Expansion_JP1_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Expansion_JP1_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave AND Expansion_JP1_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave AND NOT Expansion_JP1_avalon_parallel_port_slave_non_bursting_master_requests));
  --Expansion_JP1_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP1_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Expansion_JP1_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Expansion_JP1_avalon_parallel_port_slave_arb_share_counter <= Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Expansion_JP1_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Expansion_JP1_avalon_parallel_port_slave AND NOT Expansion_JP1_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Expansion_JP1/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Expansion_JP1_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Expansion_JP1/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Expansion_JP1_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Expansion_JP1_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave_shift_register;
  --Expansion_JP1_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Expansion_JP1/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave;
  --allow new arb cycle for Expansion_JP1/avalon_parallel_port_slave, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Expansion_JP1_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Expansion_JP1_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Expansion_JP1_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_reset <= NOT reset_n;
  Expansion_JP1_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave;
  --Expansion_JP1_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Expansion_JP1_avalon_parallel_port_slave_begins_xfer) = '1'), Expansion_JP1_avalon_parallel_port_slave_unreg_firsttransfer, Expansion_JP1_avalon_parallel_port_slave_reg_firsttransfer);
  --Expansion_JP1_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Expansion_JP1_avalon_parallel_port_slave_slavearbiterlockenable AND Expansion_JP1_avalon_parallel_port_slave_any_continuerequest));
  --Expansion_JP1_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP1_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Expansion_JP1_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Expansion_JP1_avalon_parallel_port_slave_reg_firsttransfer <= Expansion_JP1_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Expansion_JP1_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_beginbursttransfer_internal <= Expansion_JP1_avalon_parallel_port_slave_begins_xfer;
  --Expansion_JP1_avalon_parallel_port_slave_read assignment, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_read;
  --Expansion_JP1_avalon_parallel_port_slave_write assignment, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Expansion_JP1_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Expansion_JP1_avalon_parallel_port_slave_address mux, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Expansion_JP1_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer <= Expansion_JP1_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Expansion_JP1_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Expansion_JP1_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Expansion_JP1_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Expansion_JP1_avalon_parallel_port_slave_in_a_read_cycle;
  --Expansion_JP1_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Expansion_JP1_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Expansion_JP1_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Expansion_JP1_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Expansion_JP1_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Expansion_JP1_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Expansion_JP1_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign Expansion_JP1_avalon_parallel_port_slave_irq_from_sa = Expansion_JP1_avalon_parallel_port_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Expansion_JP1_avalon_parallel_port_slave_irq_from_sa <= Expansion_JP1_avalon_parallel_port_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave;
--synthesis translate_off
    --Expansion_JP1/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Expansion_JP2_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Expansion_JP2_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Expansion_JP2_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Expansion_JP2_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Expansion_JP2_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Expansion_JP2_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Expansion_JP2_avalon_parallel_port_slave_arbitrator;


architecture europa of Expansion_JP2_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Expansion_JP2_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Expansion_JP2_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Expansion_JP2_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Expansion_JP2_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave);
  --assign Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa = Expansion_JP2_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa <= Expansion_JP2_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000001110000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register_in;
  --Expansion_JP2_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Expansion_JP2_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave;
  --Expansion_JP2_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Expansion_JP2_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Expansion_JP2_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Expansion_JP2_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Expansion_JP2_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Expansion_JP2_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_allgrants <= Expansion_JP2_avalon_parallel_port_slave_grant_vector;
  --Expansion_JP2_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_end_xfer <= NOT ((Expansion_JP2_avalon_parallel_port_slave_waits_for_read OR Expansion_JP2_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave <= Expansion_JP2_avalon_parallel_port_slave_end_xfer AND (((NOT Expansion_JP2_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Expansion_JP2_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave AND Expansion_JP2_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave AND NOT Expansion_JP2_avalon_parallel_port_slave_non_bursting_master_requests));
  --Expansion_JP2_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP2_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Expansion_JP2_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Expansion_JP2_avalon_parallel_port_slave_arb_share_counter <= Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Expansion_JP2_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Expansion_JP2_avalon_parallel_port_slave AND NOT Expansion_JP2_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Expansion_JP2/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Expansion_JP2_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Expansion_JP2/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Expansion_JP2_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Expansion_JP2_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave_shift_register;
  --Expansion_JP2_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Expansion_JP2/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave;
  --allow new arb cycle for Expansion_JP2/avalon_parallel_port_slave, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Expansion_JP2_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Expansion_JP2_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Expansion_JP2_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_reset <= NOT reset_n;
  Expansion_JP2_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave;
  --Expansion_JP2_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Expansion_JP2_avalon_parallel_port_slave_begins_xfer) = '1'), Expansion_JP2_avalon_parallel_port_slave_unreg_firsttransfer, Expansion_JP2_avalon_parallel_port_slave_reg_firsttransfer);
  --Expansion_JP2_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Expansion_JP2_avalon_parallel_port_slave_slavearbiterlockenable AND Expansion_JP2_avalon_parallel_port_slave_any_continuerequest));
  --Expansion_JP2_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Expansion_JP2_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Expansion_JP2_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Expansion_JP2_avalon_parallel_port_slave_reg_firsttransfer <= Expansion_JP2_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Expansion_JP2_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_beginbursttransfer_internal <= Expansion_JP2_avalon_parallel_port_slave_begins_xfer;
  --Expansion_JP2_avalon_parallel_port_slave_read assignment, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_read;
  --Expansion_JP2_avalon_parallel_port_slave_write assignment, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Expansion_JP2_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Expansion_JP2_avalon_parallel_port_slave_address mux, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Expansion_JP2_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer <= Expansion_JP2_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Expansion_JP2_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Expansion_JP2_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Expansion_JP2_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Expansion_JP2_avalon_parallel_port_slave_in_a_read_cycle;
  --Expansion_JP2_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Expansion_JP2_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Expansion_JP2_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Expansion_JP2_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Expansion_JP2_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Expansion_JP2_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Expansion_JP2_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign Expansion_JP2_avalon_parallel_port_slave_irq_from_sa = Expansion_JP2_avalon_parallel_port_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Expansion_JP2_avalon_parallel_port_slave_irq_from_sa <= Expansion_JP2_avalon_parallel_port_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave;
--synthesis translate_off
    --Expansion_JP2/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity External_Clocks_avalon_clocks_slave_arbitrator is 
        port (
              -- inputs:
                 signal External_Clocks_avalon_clocks_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal nios_system_clock_0_out_address_to_slave : IN STD_LOGIC;
                 signal nios_system_clock_0_out_read : IN STD_LOGIC;
                 signal nios_system_clock_0_out_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal External_Clocks_avalon_clocks_slave_address : OUT STD_LOGIC;
                 signal External_Clocks_avalon_clocks_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal d1_External_Clocks_avalon_clocks_slave_end_xfer : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC
              );
end entity External_Clocks_avalon_clocks_slave_arbitrator;


architecture europa of External_Clocks_avalon_clocks_slave_arbitrator is
                signal External_Clocks_avalon_clocks_slave_allgrants :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_any_continuerequest :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_arb_counter_enable :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_arb_share_counter :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_arb_share_set_values :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_begins_xfer :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_end_xfer :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_firsttransfer :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_grant_vector :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_in_a_read_cycle :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_in_a_write_cycle :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_master_qreq_vector :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_non_bursting_master_requests :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_reg_firsttransfer :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_slavearbiterlockenable :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_unreg_firsttransfer :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_waits_for_read :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal internal_nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_arbiterlock :  STD_LOGIC;
                signal nios_system_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal nios_system_clock_0_out_continuerequest :  STD_LOGIC;
                signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register :  STD_LOGIC;
                signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register_in :  STD_LOGIC;
                signal nios_system_clock_0_out_saved_grant_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal p1_nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register :  STD_LOGIC;
                signal wait_for_External_Clocks_avalon_clocks_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT External_Clocks_avalon_clocks_slave_end_xfer;
    end if;

  end process;

  External_Clocks_avalon_clocks_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave);
  --assign External_Clocks_avalon_clocks_slave_readdata_from_sa = External_Clocks_avalon_clocks_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  External_Clocks_avalon_clocks_slave_readdata_from_sa <= External_Clocks_avalon_clocks_slave_readdata;
  internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios_system_clock_0_out_read OR nios_system_clock_0_out_write))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios_system_clock_0_out_read)))));
  --External_Clocks_avalon_clocks_slave_arb_share_counter set values, which is an e_mux
  External_Clocks_avalon_clocks_slave_arb_share_set_values <= std_logic'('1');
  --External_Clocks_avalon_clocks_slave_non_bursting_master_requests mux, which is an e_mux
  External_Clocks_avalon_clocks_slave_non_bursting_master_requests <= internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave;
  --External_Clocks_avalon_clocks_slave_any_bursting_master_saved_grant mux, which is an e_mux
  External_Clocks_avalon_clocks_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --External_Clocks_avalon_clocks_slave_arb_share_counter_next_value assignment, which is an e_assign
  External_Clocks_avalon_clocks_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(External_Clocks_avalon_clocks_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(External_Clocks_avalon_clocks_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(External_Clocks_avalon_clocks_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(External_Clocks_avalon_clocks_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --External_Clocks_avalon_clocks_slave_allgrants all slave grants, which is an e_mux
  External_Clocks_avalon_clocks_slave_allgrants <= External_Clocks_avalon_clocks_slave_grant_vector;
  --External_Clocks_avalon_clocks_slave_end_xfer assignment, which is an e_assign
  External_Clocks_avalon_clocks_slave_end_xfer <= NOT ((External_Clocks_avalon_clocks_slave_waits_for_read OR External_Clocks_avalon_clocks_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave <= External_Clocks_avalon_clocks_slave_end_xfer AND (((NOT External_Clocks_avalon_clocks_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --External_Clocks_avalon_clocks_slave_arb_share_counter arbitration counter enable, which is an e_assign
  External_Clocks_avalon_clocks_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave AND External_Clocks_avalon_clocks_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave AND NOT External_Clocks_avalon_clocks_slave_non_bursting_master_requests));
  --External_Clocks_avalon_clocks_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      External_Clocks_avalon_clocks_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(External_Clocks_avalon_clocks_slave_arb_counter_enable) = '1' then 
        External_Clocks_avalon_clocks_slave_arb_share_counter <= External_Clocks_avalon_clocks_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --External_Clocks_avalon_clocks_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      External_Clocks_avalon_clocks_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((External_Clocks_avalon_clocks_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave)) OR ((end_xfer_arb_share_counter_term_External_Clocks_avalon_clocks_slave AND NOT External_Clocks_avalon_clocks_slave_non_bursting_master_requests)))) = '1' then 
        External_Clocks_avalon_clocks_slave_slavearbiterlockenable <= External_Clocks_avalon_clocks_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios_system_clock_0/out External_Clocks/avalon_clocks_slave arbiterlock, which is an e_assign
  nios_system_clock_0_out_arbiterlock <= External_Clocks_avalon_clocks_slave_slavearbiterlockenable AND nios_system_clock_0_out_continuerequest;
  --External_Clocks_avalon_clocks_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  External_Clocks_avalon_clocks_slave_slavearbiterlockenable2 <= External_Clocks_avalon_clocks_slave_arb_share_counter_next_value;
  --nios_system_clock_0/out External_Clocks/avalon_clocks_slave arbiterlock2, which is an e_assign
  nios_system_clock_0_out_arbiterlock2 <= External_Clocks_avalon_clocks_slave_slavearbiterlockenable2 AND nios_system_clock_0_out_continuerequest;
  --External_Clocks_avalon_clocks_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  External_Clocks_avalon_clocks_slave_any_continuerequest <= std_logic'('1');
  --nios_system_clock_0_out_continuerequest continued request, which is an e_assign
  nios_system_clock_0_out_continuerequest <= std_logic'('1');
  internal_nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave AND NOT ((nios_system_clock_0_out_read AND (nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register)));
  --nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register_in <= ((internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave AND nios_system_clock_0_out_read) AND NOT External_Clocks_avalon_clocks_slave_waits_for_read) AND NOT (nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register);
  --shift register p1 nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register) & A_ToStdLogicVector(nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register_in)));
  --nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register <= p1_nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register;
    end if;

  end process;

  --local readdatavalid nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave, which is an e_mux
  nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave <= nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave_shift_register;
  --master is always granted when requested
  internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave;
  --nios_system_clock_0/out saved-grant External_Clocks/avalon_clocks_slave, which is an e_assign
  nios_system_clock_0_out_saved_grant_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave;
  --allow new arb cycle for External_Clocks/avalon_clocks_slave, which is an e_assign
  External_Clocks_avalon_clocks_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  External_Clocks_avalon_clocks_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  External_Clocks_avalon_clocks_slave_master_qreq_vector <= std_logic'('1');
  --External_Clocks_avalon_clocks_slave_firsttransfer first transaction, which is an e_assign
  External_Clocks_avalon_clocks_slave_firsttransfer <= A_WE_StdLogic((std_logic'(External_Clocks_avalon_clocks_slave_begins_xfer) = '1'), External_Clocks_avalon_clocks_slave_unreg_firsttransfer, External_Clocks_avalon_clocks_slave_reg_firsttransfer);
  --External_Clocks_avalon_clocks_slave_unreg_firsttransfer first transaction, which is an e_assign
  External_Clocks_avalon_clocks_slave_unreg_firsttransfer <= NOT ((External_Clocks_avalon_clocks_slave_slavearbiterlockenable AND External_Clocks_avalon_clocks_slave_any_continuerequest));
  --External_Clocks_avalon_clocks_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      External_Clocks_avalon_clocks_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(External_Clocks_avalon_clocks_slave_begins_xfer) = '1' then 
        External_Clocks_avalon_clocks_slave_reg_firsttransfer <= External_Clocks_avalon_clocks_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --External_Clocks_avalon_clocks_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  External_Clocks_avalon_clocks_slave_beginbursttransfer_internal <= External_Clocks_avalon_clocks_slave_begins_xfer;
  --External_Clocks_avalon_clocks_slave_address mux, which is an e_mux
  External_Clocks_avalon_clocks_slave_address <= nios_system_clock_0_out_address_to_slave;
  --d1_External_Clocks_avalon_clocks_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_External_Clocks_avalon_clocks_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_External_Clocks_avalon_clocks_slave_end_xfer <= External_Clocks_avalon_clocks_slave_end_xfer;
    end if;

  end process;

  --External_Clocks_avalon_clocks_slave_waits_for_read in a cycle, which is an e_mux
  External_Clocks_avalon_clocks_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(External_Clocks_avalon_clocks_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --External_Clocks_avalon_clocks_slave_in_a_read_cycle assignment, which is an e_assign
  External_Clocks_avalon_clocks_slave_in_a_read_cycle <= internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave AND nios_system_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= External_Clocks_avalon_clocks_slave_in_a_read_cycle;
  --External_Clocks_avalon_clocks_slave_waits_for_write in a cycle, which is an e_mux
  External_Clocks_avalon_clocks_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(External_Clocks_avalon_clocks_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --External_Clocks_avalon_clocks_slave_in_a_write_cycle assignment, which is an e_assign
  External_Clocks_avalon_clocks_slave_in_a_write_cycle <= internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave AND nios_system_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= External_Clocks_avalon_clocks_slave_in_a_write_cycle;
  wait_for_External_Clocks_avalon_clocks_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave;
  --vhdl renameroo for output signals
  nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave;
  --vhdl renameroo for output signals
  nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave <= internal_nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave;
--synthesis translate_off
    --External_Clocks/avalon_clocks_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Green_LEDs_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Green_LEDs_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Green_LEDs_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Green_LEDs_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Green_LEDs_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Green_LEDs_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Green_LEDs_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Green_LEDs_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Green_LEDs_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Green_LEDs_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Green_LEDs_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Green_LEDs_avalon_parallel_port_slave_arbitrator;


architecture europa of Green_LEDs_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Green_LEDs_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Green_LEDs_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Green_LEDs_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Green_LEDs_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave);
  --assign Green_LEDs_avalon_parallel_port_slave_readdata_from_sa = Green_LEDs_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_readdata_from_sa <= Green_LEDs_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000000010000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register_in;
  --Green_LEDs_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Green_LEDs_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave;
  --Green_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Green_LEDs_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Green_LEDs_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Green_LEDs_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Green_LEDs_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Green_LEDs_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_allgrants <= Green_LEDs_avalon_parallel_port_slave_grant_vector;
  --Green_LEDs_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_end_xfer <= NOT ((Green_LEDs_avalon_parallel_port_slave_waits_for_read OR Green_LEDs_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave <= Green_LEDs_avalon_parallel_port_slave_end_xfer AND (((NOT Green_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Green_LEDs_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave AND Green_LEDs_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave AND NOT Green_LEDs_avalon_parallel_port_slave_non_bursting_master_requests));
  --Green_LEDs_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Green_LEDs_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Green_LEDs_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Green_LEDs_avalon_parallel_port_slave_arb_share_counter <= Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Green_LEDs_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Green_LEDs_avalon_parallel_port_slave AND NOT Green_LEDs_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Green_LEDs/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Green_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Green_LEDs/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Green_LEDs_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Green_LEDs_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave_shift_register;
  --Green_LEDs_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Green_LEDs/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave;
  --allow new arb cycle for Green_LEDs/avalon_parallel_port_slave, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Green_LEDs_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Green_LEDs_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Green_LEDs_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_reset <= NOT reset_n;
  Green_LEDs_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave;
  --Green_LEDs_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Green_LEDs_avalon_parallel_port_slave_begins_xfer) = '1'), Green_LEDs_avalon_parallel_port_slave_unreg_firsttransfer, Green_LEDs_avalon_parallel_port_slave_reg_firsttransfer);
  --Green_LEDs_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Green_LEDs_avalon_parallel_port_slave_slavearbiterlockenable AND Green_LEDs_avalon_parallel_port_slave_any_continuerequest));
  --Green_LEDs_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Green_LEDs_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Green_LEDs_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Green_LEDs_avalon_parallel_port_slave_reg_firsttransfer <= Green_LEDs_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Green_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal <= Green_LEDs_avalon_parallel_port_slave_begins_xfer;
  --Green_LEDs_avalon_parallel_port_slave_read assignment, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_read;
  --Green_LEDs_avalon_parallel_port_slave_write assignment, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Green_LEDs_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Green_LEDs_avalon_parallel_port_slave_address mux, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Green_LEDs_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Green_LEDs_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Green_LEDs_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Green_LEDs_avalon_parallel_port_slave_end_xfer <= Green_LEDs_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Green_LEDs_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Green_LEDs_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Green_LEDs_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Green_LEDs_avalon_parallel_port_slave_in_a_read_cycle;
  --Green_LEDs_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Green_LEDs_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Green_LEDs_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Green_LEDs_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Green_LEDs_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Green_LEDs_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Green_LEDs_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Green_LEDs_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave;
--synthesis translate_off
    --Green_LEDs/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity HEX3_HEX0_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX3_HEX0_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal HEX3_HEX0_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal HEX3_HEX0_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal HEX3_HEX0_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal HEX3_HEX0_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX3_HEX0_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal HEX3_HEX0_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal HEX3_HEX0_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity HEX3_HEX0_avalon_parallel_port_slave_arbitrator;


architecture europa of HEX3_HEX0_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_HEX3_HEX0_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_HEX3_HEX0_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT HEX3_HEX0_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  HEX3_HEX0_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave);
  --assign HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa = HEX3_HEX0_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa <= HEX3_HEX0_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000000100000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register_in;
  --HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --HEX3_HEX0_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave;
  --HEX3_HEX0_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(HEX3_HEX0_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (HEX3_HEX0_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --HEX3_HEX0_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_allgrants <= HEX3_HEX0_avalon_parallel_port_slave_grant_vector;
  --HEX3_HEX0_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_end_xfer <= NOT ((HEX3_HEX0_avalon_parallel_port_slave_waits_for_read OR HEX3_HEX0_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave <= HEX3_HEX0_avalon_parallel_port_slave_end_xfer AND (((NOT HEX3_HEX0_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave AND HEX3_HEX0_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave AND NOT HEX3_HEX0_avalon_parallel_port_slave_non_bursting_master_requests));
  --HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(HEX3_HEX0_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter <= HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((HEX3_HEX0_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_HEX3_HEX0_avalon_parallel_port_slave AND NOT HEX3_HEX0_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master HEX3_HEX0/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(HEX3_HEX0_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master HEX3_HEX0/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --HEX3_HEX0_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT HEX3_HEX0_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave_shift_register;
  --HEX3_HEX0_avalon_parallel_port_slave_writedata mux, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave;
  --CPU/data_master saved-grant HEX3_HEX0/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave;
  --allow new arb cycle for HEX3_HEX0/avalon_parallel_port_slave, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  HEX3_HEX0_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  HEX3_HEX0_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~HEX3_HEX0_avalon_parallel_port_slave_reset assignment, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_reset <= NOT reset_n;
  HEX3_HEX0_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave;
  --HEX3_HEX0_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(HEX3_HEX0_avalon_parallel_port_slave_begins_xfer) = '1'), HEX3_HEX0_avalon_parallel_port_slave_unreg_firsttransfer, HEX3_HEX0_avalon_parallel_port_slave_reg_firsttransfer);
  --HEX3_HEX0_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((HEX3_HEX0_avalon_parallel_port_slave_slavearbiterlockenable AND HEX3_HEX0_avalon_parallel_port_slave_any_continuerequest));
  --HEX3_HEX0_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX3_HEX0_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(HEX3_HEX0_avalon_parallel_port_slave_begins_xfer) = '1' then 
        HEX3_HEX0_avalon_parallel_port_slave_reg_firsttransfer <= HEX3_HEX0_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --HEX3_HEX0_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_beginbursttransfer_internal <= HEX3_HEX0_avalon_parallel_port_slave_begins_xfer;
  --HEX3_HEX0_avalon_parallel_port_slave_read assignment, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_read;
  --HEX3_HEX0_avalon_parallel_port_slave_write assignment, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_HEX3_HEX0_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --HEX3_HEX0_avalon_parallel_port_slave_address mux, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_HEX3_HEX0_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer <= HEX3_HEX0_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --HEX3_HEX0_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(HEX3_HEX0_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --HEX3_HEX0_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= HEX3_HEX0_avalon_parallel_port_slave_in_a_read_cycle;
  --HEX3_HEX0_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(HEX3_HEX0_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --HEX3_HEX0_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  HEX3_HEX0_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= HEX3_HEX0_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_HEX3_HEX0_avalon_parallel_port_slave_counter <= std_logic'('0');
  --HEX3_HEX0_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  HEX3_HEX0_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave;
--synthesis translate_off
    --HEX3_HEX0/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity HEX7_HEX4_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX7_HEX4_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal HEX7_HEX4_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal HEX7_HEX4_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal HEX7_HEX4_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal HEX7_HEX4_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal HEX7_HEX4_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal HEX7_HEX4_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal HEX7_HEX4_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity HEX7_HEX4_avalon_parallel_port_slave_arbitrator;


architecture europa of HEX7_HEX4_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_HEX7_HEX4_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_HEX7_HEX4_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT HEX7_HEX4_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  HEX7_HEX4_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave);
  --assign HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa = HEX7_HEX4_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa <= HEX7_HEX4_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000000110000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register_in;
  --HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --HEX7_HEX4_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave;
  --HEX7_HEX4_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(HEX7_HEX4_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (HEX7_HEX4_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --HEX7_HEX4_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_allgrants <= HEX7_HEX4_avalon_parallel_port_slave_grant_vector;
  --HEX7_HEX4_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_end_xfer <= NOT ((HEX7_HEX4_avalon_parallel_port_slave_waits_for_read OR HEX7_HEX4_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave <= HEX7_HEX4_avalon_parallel_port_slave_end_xfer AND (((NOT HEX7_HEX4_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave AND HEX7_HEX4_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave AND NOT HEX7_HEX4_avalon_parallel_port_slave_non_bursting_master_requests));
  --HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(HEX7_HEX4_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter <= HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((HEX7_HEX4_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_HEX7_HEX4_avalon_parallel_port_slave AND NOT HEX7_HEX4_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master HEX7_HEX4/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(HEX7_HEX4_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master HEX7_HEX4/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --HEX7_HEX4_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT HEX7_HEX4_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave_shift_register;
  --HEX7_HEX4_avalon_parallel_port_slave_writedata mux, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave;
  --CPU/data_master saved-grant HEX7_HEX4/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave;
  --allow new arb cycle for HEX7_HEX4/avalon_parallel_port_slave, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  HEX7_HEX4_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  HEX7_HEX4_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~HEX7_HEX4_avalon_parallel_port_slave_reset assignment, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_reset <= NOT reset_n;
  HEX7_HEX4_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave;
  --HEX7_HEX4_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(HEX7_HEX4_avalon_parallel_port_slave_begins_xfer) = '1'), HEX7_HEX4_avalon_parallel_port_slave_unreg_firsttransfer, HEX7_HEX4_avalon_parallel_port_slave_reg_firsttransfer);
  --HEX7_HEX4_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((HEX7_HEX4_avalon_parallel_port_slave_slavearbiterlockenable AND HEX7_HEX4_avalon_parallel_port_slave_any_continuerequest));
  --HEX7_HEX4_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      HEX7_HEX4_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(HEX7_HEX4_avalon_parallel_port_slave_begins_xfer) = '1' then 
        HEX7_HEX4_avalon_parallel_port_slave_reg_firsttransfer <= HEX7_HEX4_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --HEX7_HEX4_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_beginbursttransfer_internal <= HEX7_HEX4_avalon_parallel_port_slave_begins_xfer;
  --HEX7_HEX4_avalon_parallel_port_slave_read assignment, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_read;
  --HEX7_HEX4_avalon_parallel_port_slave_write assignment, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_HEX7_HEX4_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --HEX7_HEX4_avalon_parallel_port_slave_address mux, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_HEX7_HEX4_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer <= HEX7_HEX4_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --HEX7_HEX4_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(HEX7_HEX4_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --HEX7_HEX4_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= HEX7_HEX4_avalon_parallel_port_slave_in_a_read_cycle;
  --HEX7_HEX4_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(HEX7_HEX4_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --HEX7_HEX4_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  HEX7_HEX4_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= HEX7_HEX4_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_HEX7_HEX4_avalon_parallel_port_slave_counter <= std_logic'('0');
  --HEX7_HEX4_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  HEX7_HEX4_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave <= internal_CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave;
--synthesis translate_off
    --HEX7_HEX4/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Interval_Timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Interval_Timer_s1_irq : IN STD_LOGIC;
                 signal Interval_Timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Interval_Timer_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Interval_Timer_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Interval_Timer_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Interval_Timer_s1 : OUT STD_LOGIC;
                 signal Interval_Timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal Interval_Timer_s1_chipselect : OUT STD_LOGIC;
                 signal Interval_Timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal Interval_Timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal Interval_Timer_s1_reset_n : OUT STD_LOGIC;
                 signal Interval_Timer_s1_write_n : OUT STD_LOGIC;
                 signal Interval_Timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_Interval_Timer_s1_end_xfer : OUT STD_LOGIC
              );
end entity Interval_Timer_s1_arbitrator;


architecture europa of Interval_Timer_s1_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Interval_Timer_s1 :  STD_LOGIC;
                signal Interval_Timer_s1_allgrants :  STD_LOGIC;
                signal Interval_Timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal Interval_Timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Interval_Timer_s1_any_continuerequest :  STD_LOGIC;
                signal Interval_Timer_s1_arb_counter_enable :  STD_LOGIC;
                signal Interval_Timer_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Interval_Timer_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Interval_Timer_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Interval_Timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal Interval_Timer_s1_begins_xfer :  STD_LOGIC;
                signal Interval_Timer_s1_end_xfer :  STD_LOGIC;
                signal Interval_Timer_s1_firsttransfer :  STD_LOGIC;
                signal Interval_Timer_s1_grant_vector :  STD_LOGIC;
                signal Interval_Timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal Interval_Timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal Interval_Timer_s1_master_qreq_vector :  STD_LOGIC;
                signal Interval_Timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal Interval_Timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal Interval_Timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal Interval_Timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal Interval_Timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal Interval_Timer_s1_waits_for_read :  STD_LOGIC;
                signal Interval_Timer_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Interval_Timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Interval_Timer_s1 :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Interval_Timer_s1 :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Interval_Timer_s1 :  STD_LOGIC;
                signal shifted_address_to_Interval_Timer_s1_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Interval_Timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Interval_Timer_s1_end_xfer;
    end if;

  end process;

  Interval_Timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Interval_Timer_s1);
  --assign Interval_Timer_s1_readdata_from_sa = Interval_Timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Interval_Timer_s1_readdata_from_sa <= Interval_Timer_s1_readdata;
  internal_CPU_data_master_requests_Interval_Timer_s1 <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("10000000000000010000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --Interval_Timer_s1_arb_share_counter set values, which is an e_mux
  Interval_Timer_s1_arb_share_set_values <= std_logic_vector'("001");
  --Interval_Timer_s1_non_bursting_master_requests mux, which is an e_mux
  Interval_Timer_s1_non_bursting_master_requests <= internal_CPU_data_master_requests_Interval_Timer_s1;
  --Interval_Timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  Interval_Timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --Interval_Timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  Interval_Timer_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Interval_Timer_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Interval_Timer_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Interval_Timer_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Interval_Timer_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Interval_Timer_s1_allgrants all slave grants, which is an e_mux
  Interval_Timer_s1_allgrants <= Interval_Timer_s1_grant_vector;
  --Interval_Timer_s1_end_xfer assignment, which is an e_assign
  Interval_Timer_s1_end_xfer <= NOT ((Interval_Timer_s1_waits_for_read OR Interval_Timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_Interval_Timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Interval_Timer_s1 <= Interval_Timer_s1_end_xfer AND (((NOT Interval_Timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Interval_Timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  Interval_Timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Interval_Timer_s1 AND Interval_Timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_Interval_Timer_s1 AND NOT Interval_Timer_s1_non_bursting_master_requests));
  --Interval_Timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Interval_Timer_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Interval_Timer_s1_arb_counter_enable) = '1' then 
        Interval_Timer_s1_arb_share_counter <= Interval_Timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Interval_Timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Interval_Timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Interval_Timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_Interval_Timer_s1)) OR ((end_xfer_arb_share_counter_term_Interval_Timer_s1 AND NOT Interval_Timer_s1_non_bursting_master_requests)))) = '1' then 
        Interval_Timer_s1_slavearbiterlockenable <= or_reduce(Interval_Timer_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Interval_Timer/s1 arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Interval_Timer_s1_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Interval_Timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Interval_Timer_s1_slavearbiterlockenable2 <= or_reduce(Interval_Timer_s1_arb_share_counter_next_value);
  --CPU/data_master Interval_Timer/s1 arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Interval_Timer_s1_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Interval_Timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  Interval_Timer_s1_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Interval_Timer_s1 <= internal_CPU_data_master_requests_Interval_Timer_s1 AND NOT (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write));
  --Interval_Timer_s1_writedata mux, which is an e_mux
  Interval_Timer_s1_writedata <= CPU_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_CPU_data_master_granted_Interval_Timer_s1 <= internal_CPU_data_master_qualified_request_Interval_Timer_s1;
  --CPU/data_master saved-grant Interval_Timer/s1, which is an e_assign
  CPU_data_master_saved_grant_Interval_Timer_s1 <= internal_CPU_data_master_requests_Interval_Timer_s1;
  --allow new arb cycle for Interval_Timer/s1, which is an e_assign
  Interval_Timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Interval_Timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Interval_Timer_s1_master_qreq_vector <= std_logic'('1');
  --Interval_Timer_s1_reset_n assignment, which is an e_assign
  Interval_Timer_s1_reset_n <= reset_n;
  Interval_Timer_s1_chipselect <= internal_CPU_data_master_granted_Interval_Timer_s1;
  --Interval_Timer_s1_firsttransfer first transaction, which is an e_assign
  Interval_Timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(Interval_Timer_s1_begins_xfer) = '1'), Interval_Timer_s1_unreg_firsttransfer, Interval_Timer_s1_reg_firsttransfer);
  --Interval_Timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  Interval_Timer_s1_unreg_firsttransfer <= NOT ((Interval_Timer_s1_slavearbiterlockenable AND Interval_Timer_s1_any_continuerequest));
  --Interval_Timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Interval_Timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Interval_Timer_s1_begins_xfer) = '1' then 
        Interval_Timer_s1_reg_firsttransfer <= Interval_Timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Interval_Timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Interval_Timer_s1_beginbursttransfer_internal <= Interval_Timer_s1_begins_xfer;
  --~Interval_Timer_s1_write_n assignment, which is an e_mux
  Interval_Timer_s1_write_n <= NOT ((internal_CPU_data_master_granted_Interval_Timer_s1 AND CPU_data_master_write));
  shifted_address_to_Interval_Timer_s1_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Interval_Timer_s1_address mux, which is an e_mux
  Interval_Timer_s1_address <= A_EXT (A_SRL(shifted_address_to_Interval_Timer_s1_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_Interval_Timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Interval_Timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Interval_Timer_s1_end_xfer <= Interval_Timer_s1_end_xfer;
    end if;

  end process;

  --Interval_Timer_s1_waits_for_read in a cycle, which is an e_mux
  Interval_Timer_s1_waits_for_read <= Interval_Timer_s1_in_a_read_cycle AND Interval_Timer_s1_begins_xfer;
  --Interval_Timer_s1_in_a_read_cycle assignment, which is an e_assign
  Interval_Timer_s1_in_a_read_cycle <= internal_CPU_data_master_granted_Interval_Timer_s1 AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Interval_Timer_s1_in_a_read_cycle;
  --Interval_Timer_s1_waits_for_write in a cycle, which is an e_mux
  Interval_Timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Interval_Timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Interval_Timer_s1_in_a_write_cycle assignment, which is an e_assign
  Interval_Timer_s1_in_a_write_cycle <= internal_CPU_data_master_granted_Interval_Timer_s1 AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Interval_Timer_s1_in_a_write_cycle;
  wait_for_Interval_Timer_s1_counter <= std_logic'('0');
  --assign Interval_Timer_s1_irq_from_sa = Interval_Timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Interval_Timer_s1_irq_from_sa <= Interval_Timer_s1_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Interval_Timer_s1 <= internal_CPU_data_master_granted_Interval_Timer_s1;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Interval_Timer_s1 <= internal_CPU_data_master_qualified_request_Interval_Timer_s1;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Interval_Timer_s1 <= internal_CPU_data_master_requests_Interval_Timer_s1;
--synthesis translate_off
    --Interval_Timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity JTAG_UART_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal JTAG_UART_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal JTAG_UART_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal JTAG_UART_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal JTAG_UART_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_JTAG_UART_avalon_jtag_slave_end_xfer : OUT STD_LOGIC
              );
end entity JTAG_UART_avalon_jtag_slave_arbitrator;


architecture europa of JTAG_UART_avalon_jtag_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal internal_JTAG_UART_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal shifted_address_to_JTAG_UART_avalon_jtag_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_JTAG_UART_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT JTAG_UART_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  JTAG_UART_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave);
  --assign JTAG_UART_avalon_jtag_slave_readdata_from_sa = JTAG_UART_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  JTAG_UART_avalon_jtag_slave_readdata_from_sa <= JTAG_UART_avalon_jtag_slave_readdata;
  internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("10000000000000001000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign JTAG_UART_avalon_jtag_slave_dataavailable_from_sa = JTAG_UART_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  JTAG_UART_avalon_jtag_slave_dataavailable_from_sa <= JTAG_UART_avalon_jtag_slave_dataavailable;
  --assign JTAG_UART_avalon_jtag_slave_readyfordata_from_sa = JTAG_UART_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  JTAG_UART_avalon_jtag_slave_readyfordata_from_sa <= JTAG_UART_avalon_jtag_slave_readyfordata;
  --assign JTAG_UART_avalon_jtag_slave_waitrequest_from_sa = JTAG_UART_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_JTAG_UART_avalon_jtag_slave_waitrequest_from_sa <= JTAG_UART_avalon_jtag_slave_waitrequest;
  --JTAG_UART_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  JTAG_UART_avalon_jtag_slave_arb_share_set_values <= std_logic_vector'("001");
  --JTAG_UART_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  JTAG_UART_avalon_jtag_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave;
  --JTAG_UART_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  JTAG_UART_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(JTAG_UART_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (JTAG_UART_avalon_jtag_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(JTAG_UART_avalon_jtag_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (JTAG_UART_avalon_jtag_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --JTAG_UART_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  JTAG_UART_avalon_jtag_slave_allgrants <= JTAG_UART_avalon_jtag_slave_grant_vector;
  --JTAG_UART_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  JTAG_UART_avalon_jtag_slave_end_xfer <= NOT ((JTAG_UART_avalon_jtag_slave_waits_for_read OR JTAG_UART_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave <= JTAG_UART_avalon_jtag_slave_end_xfer AND (((NOT JTAG_UART_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --JTAG_UART_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  JTAG_UART_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave AND JTAG_UART_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave AND NOT JTAG_UART_avalon_jtag_slave_non_bursting_master_requests));
  --JTAG_UART_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      JTAG_UART_avalon_jtag_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(JTAG_UART_avalon_jtag_slave_arb_counter_enable) = '1' then 
        JTAG_UART_avalon_jtag_slave_arb_share_counter <= JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --JTAG_UART_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      JTAG_UART_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((JTAG_UART_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_JTAG_UART_avalon_jtag_slave AND NOT JTAG_UART_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        JTAG_UART_avalon_jtag_slave_slavearbiterlockenable <= or_reduce(JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master JTAG_UART/avalon_jtag_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= JTAG_UART_avalon_jtag_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --JTAG_UART_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  JTAG_UART_avalon_jtag_slave_slavearbiterlockenable2 <= or_reduce(JTAG_UART_avalon_jtag_slave_arb_share_counter_next_value);
  --CPU/data_master JTAG_UART/avalon_jtag_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= JTAG_UART_avalon_jtag_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --JTAG_UART_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  JTAG_UART_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave AND NOT ((((CPU_data_master_read AND (NOT CPU_data_master_waitrequest))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --JTAG_UART_avalon_jtag_slave_writedata mux, which is an e_mux
  JTAG_UART_avalon_jtag_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave;
  --CPU/data_master saved-grant JTAG_UART/avalon_jtag_slave, which is an e_assign
  CPU_data_master_saved_grant_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave;
  --allow new arb cycle for JTAG_UART/avalon_jtag_slave, which is an e_assign
  JTAG_UART_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  JTAG_UART_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  JTAG_UART_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --JTAG_UART_avalon_jtag_slave_reset_n assignment, which is an e_assign
  JTAG_UART_avalon_jtag_slave_reset_n <= reset_n;
  JTAG_UART_avalon_jtag_slave_chipselect <= internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave;
  --JTAG_UART_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  JTAG_UART_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(JTAG_UART_avalon_jtag_slave_begins_xfer) = '1'), JTAG_UART_avalon_jtag_slave_unreg_firsttransfer, JTAG_UART_avalon_jtag_slave_reg_firsttransfer);
  --JTAG_UART_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  JTAG_UART_avalon_jtag_slave_unreg_firsttransfer <= NOT ((JTAG_UART_avalon_jtag_slave_slavearbiterlockenable AND JTAG_UART_avalon_jtag_slave_any_continuerequest));
  --JTAG_UART_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      JTAG_UART_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(JTAG_UART_avalon_jtag_slave_begins_xfer) = '1' then 
        JTAG_UART_avalon_jtag_slave_reg_firsttransfer <= JTAG_UART_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --JTAG_UART_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  JTAG_UART_avalon_jtag_slave_beginbursttransfer_internal <= JTAG_UART_avalon_jtag_slave_begins_xfer;
  --~JTAG_UART_avalon_jtag_slave_read_n assignment, which is an e_mux
  JTAG_UART_avalon_jtag_slave_read_n <= NOT ((internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave AND CPU_data_master_read));
  --~JTAG_UART_avalon_jtag_slave_write_n assignment, which is an e_mux
  JTAG_UART_avalon_jtag_slave_write_n <= NOT ((internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave AND CPU_data_master_write));
  shifted_address_to_JTAG_UART_avalon_jtag_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --JTAG_UART_avalon_jtag_slave_address mux, which is an e_mux
  JTAG_UART_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_JTAG_UART_avalon_jtag_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_JTAG_UART_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_JTAG_UART_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_JTAG_UART_avalon_jtag_slave_end_xfer <= JTAG_UART_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --JTAG_UART_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  JTAG_UART_avalon_jtag_slave_waits_for_read <= JTAG_UART_avalon_jtag_slave_in_a_read_cycle AND internal_JTAG_UART_avalon_jtag_slave_waitrequest_from_sa;
  --JTAG_UART_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  JTAG_UART_avalon_jtag_slave_in_a_read_cycle <= internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= JTAG_UART_avalon_jtag_slave_in_a_read_cycle;
  --JTAG_UART_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  JTAG_UART_avalon_jtag_slave_waits_for_write <= JTAG_UART_avalon_jtag_slave_in_a_write_cycle AND internal_JTAG_UART_avalon_jtag_slave_waitrequest_from_sa;
  --JTAG_UART_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  JTAG_UART_avalon_jtag_slave_in_a_write_cycle <= internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= JTAG_UART_avalon_jtag_slave_in_a_write_cycle;
  wait_for_JTAG_UART_avalon_jtag_slave_counter <= std_logic'('0');
  --assign JTAG_UART_avalon_jtag_slave_irq_from_sa = JTAG_UART_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  JTAG_UART_avalon_jtag_slave_irq_from_sa <= JTAG_UART_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_granted_JTAG_UART_avalon_jtag_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_JTAG_UART_avalon_jtag_slave <= internal_CPU_data_master_requests_JTAG_UART_avalon_jtag_slave;
  --vhdl renameroo for output signals
  JTAG_UART_avalon_jtag_slave_waitrequest_from_sa <= internal_JTAG_UART_avalon_jtag_slave_waitrequest_from_sa;
--synthesis translate_off
    --JTAG_UART/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity PS2_Port_avalon_ps2_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal PS2_Port_avalon_ps2_slave_irq : IN STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal PS2_Port_avalon_ps2_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_address : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal PS2_Port_avalon_ps2_slave_chipselect : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_irq_from_sa : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_read : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal PS2_Port_avalon_ps2_slave_reset : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_write : OUT STD_LOGIC;
                 signal PS2_Port_avalon_ps2_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_PS2_Port_avalon_ps2_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC
              );
end entity PS2_Port_avalon_ps2_slave_arbitrator;


architecture europa of PS2_Port_avalon_ps2_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_allgrants :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_any_continuerequest :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_arb_counter_enable :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_begins_xfer :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_end_xfer :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_firsttransfer :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_grant_vector :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_in_a_read_cycle :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_in_a_write_cycle :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_master_qreq_vector :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_non_bursting_master_requests :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_reg_firsttransfer :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_slavearbiterlockenable :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_unreg_firsttransfer :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_waits_for_read :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal internal_PS2_Port_avalon_ps2_slave_waitrequest_from_sa :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_PS2_Port_avalon_ps2_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_PS2_Port_avalon_ps2_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT PS2_Port_avalon_ps2_slave_end_xfer;
    end if;

  end process;

  PS2_Port_avalon_ps2_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave);
  --assign PS2_Port_avalon_ps2_slave_readdata_from_sa = PS2_Port_avalon_ps2_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  PS2_Port_avalon_ps2_slave_readdata_from_sa <= PS2_Port_avalon_ps2_slave_readdata;
  internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("10000000000000000000100000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign PS2_Port_avalon_ps2_slave_waitrequest_from_sa = PS2_Port_avalon_ps2_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_PS2_Port_avalon_ps2_slave_waitrequest_from_sa <= PS2_Port_avalon_ps2_slave_waitrequest;
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave <= CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register_in;
  --PS2_Port_avalon_ps2_slave_arb_share_counter set values, which is an e_mux
  PS2_Port_avalon_ps2_slave_arb_share_set_values <= std_logic_vector'("001");
  --PS2_Port_avalon_ps2_slave_non_bursting_master_requests mux, which is an e_mux
  PS2_Port_avalon_ps2_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave;
  --PS2_Port_avalon_ps2_slave_any_bursting_master_saved_grant mux, which is an e_mux
  PS2_Port_avalon_ps2_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --PS2_Port_avalon_ps2_slave_arb_share_counter_next_value assignment, which is an e_assign
  PS2_Port_avalon_ps2_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(PS2_Port_avalon_ps2_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (PS2_Port_avalon_ps2_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(PS2_Port_avalon_ps2_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (PS2_Port_avalon_ps2_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --PS2_Port_avalon_ps2_slave_allgrants all slave grants, which is an e_mux
  PS2_Port_avalon_ps2_slave_allgrants <= PS2_Port_avalon_ps2_slave_grant_vector;
  --PS2_Port_avalon_ps2_slave_end_xfer assignment, which is an e_assign
  PS2_Port_avalon_ps2_slave_end_xfer <= NOT ((PS2_Port_avalon_ps2_slave_waits_for_read OR PS2_Port_avalon_ps2_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave <= PS2_Port_avalon_ps2_slave_end_xfer AND (((NOT PS2_Port_avalon_ps2_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --PS2_Port_avalon_ps2_slave_arb_share_counter arbitration counter enable, which is an e_assign
  PS2_Port_avalon_ps2_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave AND PS2_Port_avalon_ps2_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave AND NOT PS2_Port_avalon_ps2_slave_non_bursting_master_requests));
  --PS2_Port_avalon_ps2_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      PS2_Port_avalon_ps2_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(PS2_Port_avalon_ps2_slave_arb_counter_enable) = '1' then 
        PS2_Port_avalon_ps2_slave_arb_share_counter <= PS2_Port_avalon_ps2_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --PS2_Port_avalon_ps2_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      PS2_Port_avalon_ps2_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((PS2_Port_avalon_ps2_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave)) OR ((end_xfer_arb_share_counter_term_PS2_Port_avalon_ps2_slave AND NOT PS2_Port_avalon_ps2_slave_non_bursting_master_requests)))) = '1' then 
        PS2_Port_avalon_ps2_slave_slavearbiterlockenable <= or_reduce(PS2_Port_avalon_ps2_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master PS2_Port/avalon_ps2_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= PS2_Port_avalon_ps2_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --PS2_Port_avalon_ps2_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  PS2_Port_avalon_ps2_slave_slavearbiterlockenable2 <= or_reduce(PS2_Port_avalon_ps2_slave_arb_share_counter_next_value);
  --CPU/data_master PS2_Port/avalon_ps2_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= PS2_Port_avalon_ps2_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --PS2_Port_avalon_ps2_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  PS2_Port_avalon_ps2_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register_in <= ((internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave AND CPU_data_master_read) AND NOT PS2_Port_avalon_ps2_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register <= p1_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave, which is an e_mux
  CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave <= CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave_shift_register;
  --PS2_Port_avalon_ps2_slave_writedata mux, which is an e_mux
  PS2_Port_avalon_ps2_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave;
  --CPU/data_master saved-grant PS2_Port/avalon_ps2_slave, which is an e_assign
  CPU_data_master_saved_grant_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave;
  --allow new arb cycle for PS2_Port/avalon_ps2_slave, which is an e_assign
  PS2_Port_avalon_ps2_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  PS2_Port_avalon_ps2_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  PS2_Port_avalon_ps2_slave_master_qreq_vector <= std_logic'('1');
  --~PS2_Port_avalon_ps2_slave_reset assignment, which is an e_assign
  PS2_Port_avalon_ps2_slave_reset <= NOT reset_n;
  PS2_Port_avalon_ps2_slave_chipselect <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave;
  --PS2_Port_avalon_ps2_slave_firsttransfer first transaction, which is an e_assign
  PS2_Port_avalon_ps2_slave_firsttransfer <= A_WE_StdLogic((std_logic'(PS2_Port_avalon_ps2_slave_begins_xfer) = '1'), PS2_Port_avalon_ps2_slave_unreg_firsttransfer, PS2_Port_avalon_ps2_slave_reg_firsttransfer);
  --PS2_Port_avalon_ps2_slave_unreg_firsttransfer first transaction, which is an e_assign
  PS2_Port_avalon_ps2_slave_unreg_firsttransfer <= NOT ((PS2_Port_avalon_ps2_slave_slavearbiterlockenable AND PS2_Port_avalon_ps2_slave_any_continuerequest));
  --PS2_Port_avalon_ps2_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      PS2_Port_avalon_ps2_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(PS2_Port_avalon_ps2_slave_begins_xfer) = '1' then 
        PS2_Port_avalon_ps2_slave_reg_firsttransfer <= PS2_Port_avalon_ps2_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --PS2_Port_avalon_ps2_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  PS2_Port_avalon_ps2_slave_beginbursttransfer_internal <= PS2_Port_avalon_ps2_slave_begins_xfer;
  --PS2_Port_avalon_ps2_slave_read assignment, which is an e_mux
  PS2_Port_avalon_ps2_slave_read <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave AND CPU_data_master_read;
  --PS2_Port_avalon_ps2_slave_write assignment, which is an e_mux
  PS2_Port_avalon_ps2_slave_write <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave AND CPU_data_master_write;
  shifted_address_to_PS2_Port_avalon_ps2_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --PS2_Port_avalon_ps2_slave_address mux, which is an e_mux
  PS2_Port_avalon_ps2_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_PS2_Port_avalon_ps2_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_PS2_Port_avalon_ps2_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_PS2_Port_avalon_ps2_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_PS2_Port_avalon_ps2_slave_end_xfer <= PS2_Port_avalon_ps2_slave_end_xfer;
    end if;

  end process;

  --PS2_Port_avalon_ps2_slave_waits_for_read in a cycle, which is an e_mux
  PS2_Port_avalon_ps2_slave_waits_for_read <= PS2_Port_avalon_ps2_slave_in_a_read_cycle AND internal_PS2_Port_avalon_ps2_slave_waitrequest_from_sa;
  --PS2_Port_avalon_ps2_slave_in_a_read_cycle assignment, which is an e_assign
  PS2_Port_avalon_ps2_slave_in_a_read_cycle <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= PS2_Port_avalon_ps2_slave_in_a_read_cycle;
  --PS2_Port_avalon_ps2_slave_waits_for_write in a cycle, which is an e_mux
  PS2_Port_avalon_ps2_slave_waits_for_write <= PS2_Port_avalon_ps2_slave_in_a_write_cycle AND internal_PS2_Port_avalon_ps2_slave_waitrequest_from_sa;
  --PS2_Port_avalon_ps2_slave_in_a_write_cycle assignment, which is an e_assign
  PS2_Port_avalon_ps2_slave_in_a_write_cycle <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= PS2_Port_avalon_ps2_slave_in_a_write_cycle;
  wait_for_PS2_Port_avalon_ps2_slave_counter <= std_logic'('0');
  --PS2_Port_avalon_ps2_slave_byteenable byte enable port mux, which is an e_mux
  PS2_Port_avalon_ps2_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign PS2_Port_avalon_ps2_slave_irq_from_sa = PS2_Port_avalon_ps2_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  PS2_Port_avalon_ps2_slave_irq_from_sa <= PS2_Port_avalon_ps2_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_granted_PS2_Port_avalon_ps2_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_PS2_Port_avalon_ps2_slave <= internal_CPU_data_master_requests_PS2_Port_avalon_ps2_slave;
  --vhdl renameroo for output signals
  PS2_Port_avalon_ps2_slave_waitrequest_from_sa <= internal_PS2_Port_avalon_ps2_slave_waitrequest_from_sa;
--synthesis translate_off
    --PS2_Port/avalon_ps2_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Pushbuttons_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Pushbuttons_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Pushbuttons_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Pushbuttons_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Pushbuttons_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Pushbuttons_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Pushbuttons_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Pushbuttons_avalon_parallel_port_slave_arbitrator;


architecture europa of Pushbuttons_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Pushbuttons_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Pushbuttons_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Pushbuttons_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Pushbuttons_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave);
  --assign Pushbuttons_avalon_parallel_port_slave_readdata_from_sa = Pushbuttons_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_readdata_from_sa <= Pushbuttons_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000001010000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register_in;
  --Pushbuttons_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Pushbuttons_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave;
  --Pushbuttons_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Pushbuttons_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Pushbuttons_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Pushbuttons_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Pushbuttons_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Pushbuttons_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_allgrants <= Pushbuttons_avalon_parallel_port_slave_grant_vector;
  --Pushbuttons_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_end_xfer <= NOT ((Pushbuttons_avalon_parallel_port_slave_waits_for_read OR Pushbuttons_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave <= Pushbuttons_avalon_parallel_port_slave_end_xfer AND (((NOT Pushbuttons_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Pushbuttons_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave AND Pushbuttons_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave AND NOT Pushbuttons_avalon_parallel_port_slave_non_bursting_master_requests));
  --Pushbuttons_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Pushbuttons_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Pushbuttons_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Pushbuttons_avalon_parallel_port_slave_arb_share_counter <= Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Pushbuttons_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Pushbuttons_avalon_parallel_port_slave AND NOT Pushbuttons_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Pushbuttons/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Pushbuttons_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Pushbuttons/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Pushbuttons_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Pushbuttons_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave_shift_register;
  --Pushbuttons_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Pushbuttons/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave;
  --allow new arb cycle for Pushbuttons/avalon_parallel_port_slave, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Pushbuttons_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Pushbuttons_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Pushbuttons_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_reset <= NOT reset_n;
  Pushbuttons_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave;
  --Pushbuttons_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Pushbuttons_avalon_parallel_port_slave_begins_xfer) = '1'), Pushbuttons_avalon_parallel_port_slave_unreg_firsttransfer, Pushbuttons_avalon_parallel_port_slave_reg_firsttransfer);
  --Pushbuttons_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Pushbuttons_avalon_parallel_port_slave_slavearbiterlockenable AND Pushbuttons_avalon_parallel_port_slave_any_continuerequest));
  --Pushbuttons_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Pushbuttons_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Pushbuttons_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Pushbuttons_avalon_parallel_port_slave_reg_firsttransfer <= Pushbuttons_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Pushbuttons_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_beginbursttransfer_internal <= Pushbuttons_avalon_parallel_port_slave_begins_xfer;
  --Pushbuttons_avalon_parallel_port_slave_read assignment, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_read;
  --Pushbuttons_avalon_parallel_port_slave_write assignment, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Pushbuttons_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Pushbuttons_avalon_parallel_port_slave_address mux, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Pushbuttons_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Pushbuttons_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Pushbuttons_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Pushbuttons_avalon_parallel_port_slave_end_xfer <= Pushbuttons_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Pushbuttons_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Pushbuttons_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Pushbuttons_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Pushbuttons_avalon_parallel_port_slave_in_a_read_cycle;
  --Pushbuttons_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Pushbuttons_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Pushbuttons_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Pushbuttons_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Pushbuttons_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Pushbuttons_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Pushbuttons_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign Pushbuttons_avalon_parallel_port_slave_irq_from_sa = Pushbuttons_avalon_parallel_port_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Pushbuttons_avalon_parallel_port_slave_irq_from_sa <= Pushbuttons_avalon_parallel_port_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave;
--synthesis translate_off
    --Pushbuttons/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Red_LEDs_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Red_LEDs_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Red_LEDs_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Red_LEDs_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Red_LEDs_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Red_LEDs_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Red_LEDs_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Red_LEDs_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Red_LEDs_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Red_LEDs_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Red_LEDs_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Red_LEDs_avalon_parallel_port_slave_arbitrator;


architecture europa of Red_LEDs_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Red_LEDs_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Red_LEDs_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Red_LEDs_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Red_LEDs_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave);
  --assign Red_LEDs_avalon_parallel_port_slave_readdata_from_sa = Red_LEDs_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_readdata_from_sa <= Red_LEDs_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register_in;
  --Red_LEDs_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Red_LEDs_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave;
  --Red_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Red_LEDs_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Red_LEDs_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Red_LEDs_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Red_LEDs_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Red_LEDs_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_allgrants <= Red_LEDs_avalon_parallel_port_slave_grant_vector;
  --Red_LEDs_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_end_xfer <= NOT ((Red_LEDs_avalon_parallel_port_slave_waits_for_read OR Red_LEDs_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave <= Red_LEDs_avalon_parallel_port_slave_end_xfer AND (((NOT Red_LEDs_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Red_LEDs_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave AND Red_LEDs_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave AND NOT Red_LEDs_avalon_parallel_port_slave_non_bursting_master_requests));
  --Red_LEDs_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Red_LEDs_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Red_LEDs_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Red_LEDs_avalon_parallel_port_slave_arb_share_counter <= Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Red_LEDs_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Red_LEDs_avalon_parallel_port_slave AND NOT Red_LEDs_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Red_LEDs/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Red_LEDs_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Red_LEDs/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Red_LEDs_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Red_LEDs_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave_shift_register;
  --Red_LEDs_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Red_LEDs/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave;
  --allow new arb cycle for Red_LEDs/avalon_parallel_port_slave, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Red_LEDs_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Red_LEDs_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Red_LEDs_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_reset <= NOT reset_n;
  Red_LEDs_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave;
  --Red_LEDs_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Red_LEDs_avalon_parallel_port_slave_begins_xfer) = '1'), Red_LEDs_avalon_parallel_port_slave_unreg_firsttransfer, Red_LEDs_avalon_parallel_port_slave_reg_firsttransfer);
  --Red_LEDs_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Red_LEDs_avalon_parallel_port_slave_slavearbiterlockenable AND Red_LEDs_avalon_parallel_port_slave_any_continuerequest));
  --Red_LEDs_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Red_LEDs_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Red_LEDs_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Red_LEDs_avalon_parallel_port_slave_reg_firsttransfer <= Red_LEDs_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Red_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_beginbursttransfer_internal <= Red_LEDs_avalon_parallel_port_slave_begins_xfer;
  --Red_LEDs_avalon_parallel_port_slave_read assignment, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_read;
  --Red_LEDs_avalon_parallel_port_slave_write assignment, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Red_LEDs_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Red_LEDs_avalon_parallel_port_slave_address mux, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Red_LEDs_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Red_LEDs_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Red_LEDs_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Red_LEDs_avalon_parallel_port_slave_end_xfer <= Red_LEDs_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Red_LEDs_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Red_LEDs_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Red_LEDs_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Red_LEDs_avalon_parallel_port_slave_in_a_read_cycle;
  --Red_LEDs_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Red_LEDs_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Red_LEDs_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Red_LEDs_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Red_LEDs_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Red_LEDs_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Red_LEDs_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Red_LEDs_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave;
--synthesis translate_off
    --Red_LEDs/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module;


architecture europa of rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module;


architecture europa of rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity SDRAM_s1_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal CPU_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_instruction_master_latency_counter : IN STD_LOGIC;
                 signal CPU_instruction_master_read : IN STD_LOGIC;
                 signal SDRAM_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SDRAM_s1_readdatavalid : IN STD_LOGIC;
                 signal SDRAM_s1_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_byteenable_SDRAM_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_granted_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SDRAM_s1_shift_register : OUT STD_LOGIC;
                 signal CPU_data_master_requests_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_instruction_master_granted_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_instruction_master_qualified_request_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_SDRAM_s1 : OUT STD_LOGIC;
                 signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : OUT STD_LOGIC;
                 signal CPU_instruction_master_requests_SDRAM_s1 : OUT STD_LOGIC;
                 signal SDRAM_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal SDRAM_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal SDRAM_s1_chipselect : OUT STD_LOGIC;
                 signal SDRAM_s1_read_n : OUT STD_LOGIC;
                 signal SDRAM_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SDRAM_s1_reset_n : OUT STD_LOGIC;
                 signal SDRAM_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal SDRAM_s1_write_n : OUT STD_LOGIC;
                 signal SDRAM_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_SDRAM_s1_end_xfer : OUT STD_LOGIC
              );
end entity SDRAM_s1_arbitrator;


architecture europa of SDRAM_s1_arbitrator is
component rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module;

component rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module;

                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_SDRAM_s1_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_byteenable_SDRAM_s1_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_rdv_fifo_empty_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_rdv_fifo_output_from_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_saved_grant_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_arbiterlock :  STD_LOGIC;
                signal CPU_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_instruction_master_continuerequest :  STD_LOGIC;
                signal CPU_instruction_master_rdv_fifo_empty_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_rdv_fifo_output_from_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_saved_grant_SDRAM_s1 :  STD_LOGIC;
                signal SDRAM_s1_allgrants :  STD_LOGIC;
                signal SDRAM_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal SDRAM_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal SDRAM_s1_any_continuerequest :  STD_LOGIC;
                signal SDRAM_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_arb_counter_enable :  STD_LOGIC;
                signal SDRAM_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SDRAM_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SDRAM_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SDRAM_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal SDRAM_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal SDRAM_s1_begins_xfer :  STD_LOGIC;
                signal SDRAM_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal SDRAM_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_end_xfer :  STD_LOGIC;
                signal SDRAM_s1_firsttransfer :  STD_LOGIC;
                signal SDRAM_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_in_a_read_cycle :  STD_LOGIC;
                signal SDRAM_s1_in_a_write_cycle :  STD_LOGIC;
                signal SDRAM_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal SDRAM_s1_non_bursting_master_requests :  STD_LOGIC;
                signal SDRAM_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal SDRAM_s1_reg_firsttransfer :  STD_LOGIC;
                signal SDRAM_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_slavearbiterlockenable :  STD_LOGIC;
                signal SDRAM_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal SDRAM_s1_unreg_firsttransfer :  STD_LOGIC;
                signal SDRAM_s1_waits_for_read :  STD_LOGIC;
                signal SDRAM_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_SDRAM_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_byteenable_SDRAM_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_CPU_data_master_granted_SDRAM_s1 :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_SDRAM_s1 :  STD_LOGIC;
                signal internal_CPU_data_master_read_data_valid_SDRAM_s1_shift_register :  STD_LOGIC;
                signal internal_CPU_data_master_requests_SDRAM_s1 :  STD_LOGIC;
                signal internal_CPU_instruction_master_granted_SDRAM_s1 :  STD_LOGIC;
                signal internal_CPU_instruction_master_qualified_request_SDRAM_s1 :  STD_LOGIC;
                signal internal_CPU_instruction_master_requests_SDRAM_s1 :  STD_LOGIC;
                signal internal_SDRAM_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_CPU_data_master_granted_slave_SDRAM_s1 :  STD_LOGIC;
                signal last_cycle_CPU_instruction_master_granted_slave_SDRAM_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal shifted_address_to_SDRAM_s1_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal shifted_address_to_SDRAM_s1_from_CPU_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_SDRAM_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT SDRAM_s1_end_xfer;
    end if;

  end process;

  SDRAM_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_CPU_data_master_qualified_request_SDRAM_s1 OR internal_CPU_instruction_master_qualified_request_SDRAM_s1));
  --assign SDRAM_s1_readdatavalid_from_sa = SDRAM_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  SDRAM_s1_readdatavalid_from_sa <= SDRAM_s1_readdatavalid;
  --assign SDRAM_s1_readdata_from_sa = SDRAM_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  SDRAM_s1_readdata_from_sa <= SDRAM_s1_readdata;
  internal_CPU_data_master_requests_SDRAM_s1 <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("00000000000000000000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign SDRAM_s1_waitrequest_from_sa = SDRAM_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_SDRAM_s1_waitrequest_from_sa <= SDRAM_s1_waitrequest;
  --SDRAM_s1_arb_share_counter set values, which is an e_mux
  SDRAM_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_CPU_instruction_master_granted_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_CPU_instruction_master_granted_SDRAM_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001"))))), 3);
  --SDRAM_s1_non_bursting_master_requests mux, which is an e_mux
  SDRAM_s1_non_bursting_master_requests <= ((internal_CPU_data_master_requests_SDRAM_s1 OR internal_CPU_instruction_master_requests_SDRAM_s1) OR internal_CPU_data_master_requests_SDRAM_s1) OR internal_CPU_instruction_master_requests_SDRAM_s1;
  --SDRAM_s1_any_bursting_master_saved_grant mux, which is an e_mux
  SDRAM_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --SDRAM_s1_arb_share_counter_next_value assignment, which is an e_assign
  SDRAM_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(SDRAM_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (SDRAM_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(SDRAM_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (SDRAM_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --SDRAM_s1_allgrants all slave grants, which is an e_mux
  SDRAM_s1_allgrants <= (((or_reduce(SDRAM_s1_grant_vector)) OR (or_reduce(SDRAM_s1_grant_vector))) OR (or_reduce(SDRAM_s1_grant_vector))) OR (or_reduce(SDRAM_s1_grant_vector));
  --SDRAM_s1_end_xfer assignment, which is an e_assign
  SDRAM_s1_end_xfer <= NOT ((SDRAM_s1_waits_for_read OR SDRAM_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_SDRAM_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_SDRAM_s1 <= SDRAM_s1_end_xfer AND (((NOT SDRAM_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --SDRAM_s1_arb_share_counter arbitration counter enable, which is an e_assign
  SDRAM_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_SDRAM_s1 AND SDRAM_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_SDRAM_s1 AND NOT SDRAM_s1_non_bursting_master_requests));
  --SDRAM_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SDRAM_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(SDRAM_s1_arb_counter_enable) = '1' then 
        SDRAM_s1_arb_share_counter <= SDRAM_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --SDRAM_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SDRAM_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(SDRAM_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_SDRAM_s1)) OR ((end_xfer_arb_share_counter_term_SDRAM_s1 AND NOT SDRAM_s1_non_bursting_master_requests)))) = '1' then 
        SDRAM_s1_slavearbiterlockenable <= or_reduce(SDRAM_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master SDRAM/s1 arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= SDRAM_s1_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --SDRAM_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  SDRAM_s1_slavearbiterlockenable2 <= or_reduce(SDRAM_s1_arb_share_counter_next_value);
  --CPU/data_master SDRAM/s1 arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= SDRAM_s1_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --CPU/instruction_master SDRAM/s1 arbiterlock, which is an e_assign
  CPU_instruction_master_arbiterlock <= SDRAM_s1_slavearbiterlockenable AND CPU_instruction_master_continuerequest;
  --CPU/instruction_master SDRAM/s1 arbiterlock2, which is an e_assign
  CPU_instruction_master_arbiterlock2 <= SDRAM_s1_slavearbiterlockenable2 AND CPU_instruction_master_continuerequest;
  --CPU/instruction_master granted SDRAM/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_CPU_instruction_master_granted_slave_SDRAM_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_CPU_instruction_master_granted_slave_SDRAM_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(CPU_instruction_master_saved_grant_SDRAM_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((SDRAM_s1_arbitration_holdoff_internal OR NOT internal_CPU_instruction_master_requests_SDRAM_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_CPU_instruction_master_granted_slave_SDRAM_s1))))));
    end if;

  end process;

  --CPU_instruction_master_continuerequest continued request, which is an e_mux
  CPU_instruction_master_continuerequest <= last_cycle_CPU_instruction_master_granted_slave_SDRAM_s1 AND internal_CPU_instruction_master_requests_SDRAM_s1;
  --SDRAM_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  SDRAM_s1_any_continuerequest <= CPU_instruction_master_continuerequest OR CPU_data_master_continuerequest;
  internal_CPU_data_master_qualified_request_SDRAM_s1 <= internal_CPU_data_master_requests_SDRAM_s1 AND NOT (((((CPU_data_master_read AND ((NOT CPU_data_master_waitrequest OR (internal_CPU_data_master_read_data_valid_SDRAM_s1_shift_register))))) OR (((((NOT CPU_data_master_waitrequest OR CPU_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_CPU_data_master_byteenable_SDRAM_s1)))) AND CPU_data_master_write))) OR CPU_instruction_master_arbiterlock));
  --unique name for SDRAM_s1_move_on_to_next_transaction, which is an e_assign
  SDRAM_s1_move_on_to_next_transaction <= SDRAM_s1_readdatavalid_from_sa;
  --rdv_fifo_for_CPU_data_master_to_SDRAM_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_CPU_data_master_to_SDRAM_s1 : rdv_fifo_for_CPU_data_master_to_SDRAM_s1_module
    port map(
      data_out => CPU_data_master_rdv_fifo_output_from_SDRAM_s1,
      empty => open,
      fifo_contains_ones_n => CPU_data_master_rdv_fifo_empty_SDRAM_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_CPU_data_master_granted_SDRAM_s1,
      read => SDRAM_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT SDRAM_s1_waits_for_read;

  internal_CPU_data_master_read_data_valid_SDRAM_s1_shift_register <= NOT CPU_data_master_rdv_fifo_empty_SDRAM_s1;
  --local readdatavalid CPU_data_master_read_data_valid_SDRAM_s1, which is an e_mux
  CPU_data_master_read_data_valid_SDRAM_s1 <= ((SDRAM_s1_readdatavalid_from_sa AND CPU_data_master_rdv_fifo_output_from_SDRAM_s1)) AND NOT CPU_data_master_rdv_fifo_empty_SDRAM_s1;
  --SDRAM_s1_writedata mux, which is an e_mux
  SDRAM_s1_writedata <= CPU_data_master_dbs_write_16;
  internal_CPU_instruction_master_requests_SDRAM_s1 <= ((to_std_logic(((Std_Logic_Vector'(CPU_instruction_master_address_to_slave(27 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("0000000000000000000000000000")))) AND (CPU_instruction_master_read))) AND CPU_instruction_master_read;
  --CPU/data_master granted SDRAM/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_CPU_data_master_granted_slave_SDRAM_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_CPU_data_master_granted_slave_SDRAM_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(CPU_data_master_saved_grant_SDRAM_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((SDRAM_s1_arbitration_holdoff_internal OR NOT internal_CPU_data_master_requests_SDRAM_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_CPU_data_master_granted_slave_SDRAM_s1))))));
    end if;

  end process;

  --CPU_data_master_continuerequest continued request, which is an e_mux
  CPU_data_master_continuerequest <= last_cycle_CPU_data_master_granted_slave_SDRAM_s1 AND internal_CPU_data_master_requests_SDRAM_s1;
  internal_CPU_instruction_master_qualified_request_SDRAM_s1 <= internal_CPU_instruction_master_requests_SDRAM_s1 AND NOT ((((CPU_instruction_master_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_latency_counter)))))))))) OR CPU_data_master_arbiterlock));
  --rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1 : rdv_fifo_for_CPU_instruction_master_to_SDRAM_s1_module
    port map(
      data_out => CPU_instruction_master_rdv_fifo_output_from_SDRAM_s1,
      empty => open,
      fifo_contains_ones_n => CPU_instruction_master_rdv_fifo_empty_SDRAM_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_CPU_instruction_master_granted_SDRAM_s1,
      read => SDRAM_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT SDRAM_s1_waits_for_read;

  CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register <= NOT CPU_instruction_master_rdv_fifo_empty_SDRAM_s1;
  --local readdatavalid CPU_instruction_master_read_data_valid_SDRAM_s1, which is an e_mux
  CPU_instruction_master_read_data_valid_SDRAM_s1 <= ((SDRAM_s1_readdatavalid_from_sa AND CPU_instruction_master_rdv_fifo_output_from_SDRAM_s1)) AND NOT CPU_instruction_master_rdv_fifo_empty_SDRAM_s1;
  --allow new arb cycle for SDRAM/s1, which is an e_assign
  SDRAM_s1_allow_new_arb_cycle <= NOT CPU_data_master_arbiterlock AND NOT CPU_instruction_master_arbiterlock;
  --CPU/instruction_master assignment into master qualified-requests vector for SDRAM/s1, which is an e_assign
  SDRAM_s1_master_qreq_vector(0) <= internal_CPU_instruction_master_qualified_request_SDRAM_s1;
  --CPU/instruction_master grant SDRAM/s1, which is an e_assign
  internal_CPU_instruction_master_granted_SDRAM_s1 <= SDRAM_s1_grant_vector(0);
  --CPU/instruction_master saved-grant SDRAM/s1, which is an e_assign
  CPU_instruction_master_saved_grant_SDRAM_s1 <= SDRAM_s1_arb_winner(0) AND internal_CPU_instruction_master_requests_SDRAM_s1;
  --CPU/data_master assignment into master qualified-requests vector for SDRAM/s1, which is an e_assign
  SDRAM_s1_master_qreq_vector(1) <= internal_CPU_data_master_qualified_request_SDRAM_s1;
  --CPU/data_master grant SDRAM/s1, which is an e_assign
  internal_CPU_data_master_granted_SDRAM_s1 <= SDRAM_s1_grant_vector(1);
  --CPU/data_master saved-grant SDRAM/s1, which is an e_assign
  CPU_data_master_saved_grant_SDRAM_s1 <= SDRAM_s1_arb_winner(1) AND internal_CPU_data_master_requests_SDRAM_s1;
  --SDRAM/s1 chosen-master double-vector, which is an e_assign
  SDRAM_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((SDRAM_s1_master_qreq_vector & SDRAM_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT SDRAM_s1_master_qreq_vector & NOT SDRAM_s1_master_qreq_vector))) + (std_logic_vector'("000") & (SDRAM_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  SDRAM_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((SDRAM_s1_allow_new_arb_cycle AND or_reduce(SDRAM_s1_grant_vector)))) = '1'), SDRAM_s1_grant_vector, SDRAM_s1_saved_chosen_master_vector);
  --saved SDRAM_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SDRAM_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(SDRAM_s1_allow_new_arb_cycle) = '1' then 
        SDRAM_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(SDRAM_s1_grant_vector)) = '1'), SDRAM_s1_grant_vector, SDRAM_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  SDRAM_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((SDRAM_s1_chosen_master_double_vector(1) OR SDRAM_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((SDRAM_s1_chosen_master_double_vector(0) OR SDRAM_s1_chosen_master_double_vector(2)))));
  --SDRAM/s1 chosen master rotated left, which is an e_assign
  SDRAM_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(SDRAM_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(SDRAM_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --SDRAM/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SDRAM_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(SDRAM_s1_grant_vector)) = '1' then 
        SDRAM_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(SDRAM_s1_end_xfer) = '1'), SDRAM_s1_chosen_master_rot_left, SDRAM_s1_grant_vector);
      end if;
    end if;

  end process;

  --SDRAM_s1_reset_n assignment, which is an e_assign
  SDRAM_s1_reset_n <= reset_n;
  SDRAM_s1_chipselect <= internal_CPU_data_master_granted_SDRAM_s1 OR internal_CPU_instruction_master_granted_SDRAM_s1;
  --SDRAM_s1_firsttransfer first transaction, which is an e_assign
  SDRAM_s1_firsttransfer <= A_WE_StdLogic((std_logic'(SDRAM_s1_begins_xfer) = '1'), SDRAM_s1_unreg_firsttransfer, SDRAM_s1_reg_firsttransfer);
  --SDRAM_s1_unreg_firsttransfer first transaction, which is an e_assign
  SDRAM_s1_unreg_firsttransfer <= NOT ((SDRAM_s1_slavearbiterlockenable AND SDRAM_s1_any_continuerequest));
  --SDRAM_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SDRAM_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(SDRAM_s1_begins_xfer) = '1' then 
        SDRAM_s1_reg_firsttransfer <= SDRAM_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --SDRAM_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  SDRAM_s1_beginbursttransfer_internal <= SDRAM_s1_begins_xfer;
  --SDRAM_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  SDRAM_s1_arbitration_holdoff_internal <= SDRAM_s1_begins_xfer AND SDRAM_s1_firsttransfer;
  --~SDRAM_s1_read_n assignment, which is an e_mux
  SDRAM_s1_read_n <= NOT ((((internal_CPU_data_master_granted_SDRAM_s1 AND CPU_data_master_read)) OR ((internal_CPU_instruction_master_granted_SDRAM_s1 AND CPU_instruction_master_read))));
  --~SDRAM_s1_write_n assignment, which is an e_mux
  SDRAM_s1_write_n <= NOT ((internal_CPU_data_master_granted_SDRAM_s1 AND CPU_data_master_write));
  shifted_address_to_SDRAM_s1_from_CPU_data_master <= A_EXT (Std_Logic_Vector'(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(CPU_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 29);
  --SDRAM_s1_address mux, which is an e_mux
  SDRAM_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SDRAM_s1)) = '1'), (A_SRL(shifted_address_to_SDRAM_s1_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000001"))), (std_logic_vector'("0") & ((A_SRL(shifted_address_to_SDRAM_s1_from_CPU_instruction_master,std_logic_vector'("00000000000000000000000000000001")))))), 22);
  shifted_address_to_SDRAM_s1_from_CPU_instruction_master <= A_EXT (Std_Logic_Vector'(A_SRL(CPU_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(CPU_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 28);
  --d1_SDRAM_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_SDRAM_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_SDRAM_s1_end_xfer <= SDRAM_s1_end_xfer;
    end if;

  end process;

  --SDRAM_s1_waits_for_read in a cycle, which is an e_mux
  SDRAM_s1_waits_for_read <= SDRAM_s1_in_a_read_cycle AND internal_SDRAM_s1_waitrequest_from_sa;
  --SDRAM_s1_in_a_read_cycle assignment, which is an e_assign
  SDRAM_s1_in_a_read_cycle <= ((internal_CPU_data_master_granted_SDRAM_s1 AND CPU_data_master_read)) OR ((internal_CPU_instruction_master_granted_SDRAM_s1 AND CPU_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= SDRAM_s1_in_a_read_cycle;
  --SDRAM_s1_waits_for_write in a cycle, which is an e_mux
  SDRAM_s1_waits_for_write <= SDRAM_s1_in_a_write_cycle AND internal_SDRAM_s1_waitrequest_from_sa;
  --SDRAM_s1_in_a_write_cycle assignment, which is an e_assign
  SDRAM_s1_in_a_write_cycle <= internal_CPU_data_master_granted_SDRAM_s1 AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= SDRAM_s1_in_a_write_cycle;
  wait_for_SDRAM_s1_counter <= std_logic'('0');
  --~SDRAM_s1_byteenable_n byte enable port mux, which is an e_mux
  SDRAM_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SDRAM_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_byteenable_SDRAM_s1)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 2);
  (CPU_data_master_byteenable_SDRAM_s1_segment_1(1), CPU_data_master_byteenable_SDRAM_s1_segment_1(0), CPU_data_master_byteenable_SDRAM_s1_segment_0(1), CPU_data_master_byteenable_SDRAM_s1_segment_0(0)) <= CPU_data_master_byteenable;
  internal_CPU_data_master_byteenable_SDRAM_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_byteenable_SDRAM_s1_segment_0, CPU_data_master_byteenable_SDRAM_s1_segment_1);
  --vhdl renameroo for output signals
  CPU_data_master_byteenable_SDRAM_s1 <= internal_CPU_data_master_byteenable_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_data_master_granted_SDRAM_s1 <= internal_CPU_data_master_granted_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_SDRAM_s1 <= internal_CPU_data_master_qualified_request_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_data_master_read_data_valid_SDRAM_s1_shift_register <= internal_CPU_data_master_read_data_valid_SDRAM_s1_shift_register;
  --vhdl renameroo for output signals
  CPU_data_master_requests_SDRAM_s1 <= internal_CPU_data_master_requests_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_instruction_master_granted_SDRAM_s1 <= internal_CPU_instruction_master_granted_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_instruction_master_qualified_request_SDRAM_s1 <= internal_CPU_instruction_master_qualified_request_SDRAM_s1;
  --vhdl renameroo for output signals
  CPU_instruction_master_requests_SDRAM_s1 <= internal_CPU_instruction_master_requests_SDRAM_s1;
  --vhdl renameroo for output signals
  SDRAM_s1_waitrequest_from_sa <= internal_SDRAM_s1_waitrequest_from_sa;
--synthesis translate_off
    --SDRAM/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_granted_SDRAM_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_CPU_instruction_master_granted_SDRAM_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(CPU_data_master_saved_grant_SDRAM_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(CPU_instruction_master_saved_grant_SDRAM_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module;


architecture europa of rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module;


architecture europa of rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity SRAM_avalon_sram_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal SRAM_avalon_sram_slave_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SRAM_avalon_sram_slave_readdatavalid : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_byteenable_SRAM_avalon_sram_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_granted_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : OUT STD_LOGIC;
                 signal CPU_data_master_requests_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal SRAM_avalon_sram_slave_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal SRAM_avalon_sram_slave_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal SRAM_avalon_sram_slave_read : OUT STD_LOGIC;
                 signal SRAM_avalon_sram_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SRAM_avalon_sram_slave_reset : OUT STD_LOGIC;
                 signal SRAM_avalon_sram_slave_write : OUT STD_LOGIC;
                 signal SRAM_avalon_sram_slave_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                 signal d1_SRAM_avalon_sram_slave_end_xfer : OUT STD_LOGIC
              );
end entity SRAM_avalon_sram_slave_arbitrator;


architecture europa of SRAM_avalon_sram_slave_arbitrator is
component rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module;

component rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module;

                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_rdv_fifo_empty_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_rdv_fifo_output_from_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_saved_grant_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_allgrants :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_any_continuerequest :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_arb_counter_enable :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SRAM_avalon_sram_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SRAM_avalon_sram_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal SRAM_avalon_sram_slave_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_begins_xfer :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal SRAM_avalon_sram_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_end_xfer :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_firsttransfer :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_in_a_read_cycle :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_in_a_write_cycle :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_move_on_to_next_transaction :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_non_bursting_master_requests :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_readdatavalid_from_sa :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_reg_firsttransfer :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_slavearbiterlockenable :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_unreg_firsttransfer :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_waits_for_read :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_waits_for_write :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock2 :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_continuerequest :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_empty_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_output_from_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_saved_grant_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_byteenable_SRAM_avalon_sram_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_CPU_data_master_granted_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal internal_CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register :  STD_LOGIC;
                signal internal_CPU_data_master_requests_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal last_cycle_CPU_data_master_granted_slave_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal last_cycle_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_slave_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal saved_chosen_master_btw_VGA_Pixel_Buffer_avalon_pixel_dma_master_and_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal shifted_address_to_SRAM_avalon_sram_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal shifted_address_to_SRAM_avalon_sram_slave_from_VGA_Pixel_Buffer_avalon_pixel_dma_master :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_SRAM_avalon_sram_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT SRAM_avalon_sram_slave_end_xfer;
    end if;

  end process;

  SRAM_avalon_sram_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_CPU_data_master_qualified_request_SRAM_avalon_sram_slave OR internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave));
  --assign SRAM_avalon_sram_slave_readdata_from_sa = SRAM_avalon_sram_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  SRAM_avalon_sram_slave_readdata_from_sa <= SRAM_avalon_sram_slave_readdata;
  internal_CPU_data_master_requests_SRAM_avalon_sram_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("01000000000000000000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign SRAM_avalon_sram_slave_readdatavalid_from_sa = SRAM_avalon_sram_slave_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  SRAM_avalon_sram_slave_readdatavalid_from_sa <= SRAM_avalon_sram_slave_readdatavalid;
  --SRAM_avalon_sram_slave_arb_share_counter set values, which is an e_mux
  SRAM_avalon_sram_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SRAM_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SRAM_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001"))), 3);
  --SRAM_avalon_sram_slave_non_bursting_master_requests mux, which is an e_mux
  SRAM_avalon_sram_slave_non_bursting_master_requests <= ((internal_CPU_data_master_requests_SRAM_avalon_sram_slave OR internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave) OR internal_CPU_data_master_requests_SRAM_avalon_sram_slave) OR internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave;
  --SRAM_avalon_sram_slave_any_bursting_master_saved_grant mux, which is an e_mux
  SRAM_avalon_sram_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --SRAM_avalon_sram_slave_arb_share_counter_next_value assignment, which is an e_assign
  SRAM_avalon_sram_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(SRAM_avalon_sram_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (SRAM_avalon_sram_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(SRAM_avalon_sram_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (SRAM_avalon_sram_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --SRAM_avalon_sram_slave_allgrants all slave grants, which is an e_mux
  SRAM_avalon_sram_slave_allgrants <= (((or_reduce(SRAM_avalon_sram_slave_grant_vector)) OR (or_reduce(SRAM_avalon_sram_slave_grant_vector))) OR (or_reduce(SRAM_avalon_sram_slave_grant_vector))) OR (or_reduce(SRAM_avalon_sram_slave_grant_vector));
  --SRAM_avalon_sram_slave_end_xfer assignment, which is an e_assign
  SRAM_avalon_sram_slave_end_xfer <= NOT ((SRAM_avalon_sram_slave_waits_for_read OR SRAM_avalon_sram_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_end_xfer AND (((NOT SRAM_avalon_sram_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --SRAM_avalon_sram_slave_arb_share_counter arbitration counter enable, which is an e_assign
  SRAM_avalon_sram_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave AND SRAM_avalon_sram_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave AND NOT SRAM_avalon_sram_slave_non_bursting_master_requests));
  --SRAM_avalon_sram_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SRAM_avalon_sram_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(SRAM_avalon_sram_slave_arb_counter_enable) = '1' then 
        SRAM_avalon_sram_slave_arb_share_counter <= SRAM_avalon_sram_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --SRAM_avalon_sram_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SRAM_avalon_sram_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(SRAM_avalon_sram_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave)) OR ((end_xfer_arb_share_counter_term_SRAM_avalon_sram_slave AND NOT SRAM_avalon_sram_slave_non_bursting_master_requests)))) = '1' then 
        SRAM_avalon_sram_slave_slavearbiterlockenable <= or_reduce(SRAM_avalon_sram_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master SRAM/avalon_sram_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= SRAM_avalon_sram_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --SRAM_avalon_sram_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  SRAM_avalon_sram_slave_slavearbiterlockenable2 <= or_reduce(SRAM_avalon_sram_slave_arb_share_counter_next_value);
  --CPU/data_master SRAM/avalon_sram_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= SRAM_avalon_sram_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --VGA_Pixel_Buffer/avalon_pixel_dma_master SRAM/avalon_sram_slave arbiterlock2, which is an e_assign
  VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock2 <= SRAM_avalon_sram_slave_slavearbiterlockenable2 AND VGA_Pixel_Buffer_avalon_pixel_dma_master_continuerequest;
  --VGA_Pixel_Buffer/avalon_pixel_dma_master granted SRAM/avalon_sram_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_slave_SRAM_avalon_sram_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_slave_SRAM_avalon_sram_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(VGA_Pixel_Buffer_avalon_pixel_dma_master_saved_grant_SRAM_avalon_sram_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((SRAM_avalon_sram_slave_arbitration_holdoff_internal OR NOT internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_slave_SRAM_avalon_sram_slave))))));
    end if;

  end process;

  --VGA_Pixel_Buffer_avalon_pixel_dma_master_continuerequest continued request, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_dma_master_continuerequest <= last_cycle_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_slave_SRAM_avalon_sram_slave AND internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave;
  --SRAM_avalon_sram_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  SRAM_avalon_sram_slave_any_continuerequest <= VGA_Pixel_Buffer_avalon_pixel_dma_master_continuerequest OR CPU_data_master_continuerequest;
  internal_CPU_data_master_qualified_request_SRAM_avalon_sram_slave <= internal_CPU_data_master_requests_SRAM_avalon_sram_slave AND NOT (((((CPU_data_master_read AND ((NOT CPU_data_master_waitrequest OR (internal_CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register))))) OR (((((NOT CPU_data_master_waitrequest OR CPU_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_CPU_data_master_byteenable_SRAM_avalon_sram_slave)))) AND CPU_data_master_write))) OR ((VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock AND (saved_chosen_master_btw_VGA_Pixel_Buffer_avalon_pixel_dma_master_and_SRAM_avalon_sram_slave)))));
  --unique name for SRAM_avalon_sram_slave_move_on_to_next_transaction, which is an e_assign
  SRAM_avalon_sram_slave_move_on_to_next_transaction <= SRAM_avalon_sram_slave_readdatavalid_from_sa;
  --rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave : rdv_fifo_for_CPU_data_master_to_SRAM_avalon_sram_slave_module
    port map(
      data_out => CPU_data_master_rdv_fifo_output_from_SRAM_avalon_sram_slave,
      empty => open,
      fifo_contains_ones_n => CPU_data_master_rdv_fifo_empty_SRAM_avalon_sram_slave,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_CPU_data_master_granted_SRAM_avalon_sram_slave,
      read => SRAM_avalon_sram_slave_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT SRAM_avalon_sram_slave_waits_for_read;

  internal_CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register <= NOT CPU_data_master_rdv_fifo_empty_SRAM_avalon_sram_slave;
  --local readdatavalid CPU_data_master_read_data_valid_SRAM_avalon_sram_slave, which is an e_mux
  CPU_data_master_read_data_valid_SRAM_avalon_sram_slave <= ((SRAM_avalon_sram_slave_readdatavalid_from_sa AND CPU_data_master_rdv_fifo_output_from_SRAM_avalon_sram_slave)) AND NOT CPU_data_master_rdv_fifo_empty_SRAM_avalon_sram_slave;
  --SRAM_avalon_sram_slave_writedata mux, which is an e_mux
  SRAM_avalon_sram_slave_writedata <= CPU_data_master_dbs_write_16;
  internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave <= ((to_std_logic(((Std_Logic_Vector'(VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave(31 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("00001000000000000000000000000000")))) AND (VGA_Pixel_Buffer_avalon_pixel_dma_master_read))) AND VGA_Pixel_Buffer_avalon_pixel_dma_master_read;
  --CPU/data_master granted SRAM/avalon_sram_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_CPU_data_master_granted_slave_SRAM_avalon_sram_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_CPU_data_master_granted_slave_SRAM_avalon_sram_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(CPU_data_master_saved_grant_SRAM_avalon_sram_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((SRAM_avalon_sram_slave_arbitration_holdoff_internal OR NOT internal_CPU_data_master_requests_SRAM_avalon_sram_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_CPU_data_master_granted_slave_SRAM_avalon_sram_slave))))));
    end if;

  end process;

  --CPU_data_master_continuerequest continued request, which is an e_mux
  CPU_data_master_continuerequest <= last_cycle_CPU_data_master_granted_slave_SRAM_avalon_sram_slave AND internal_CPU_data_master_requests_SRAM_avalon_sram_slave;
  internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave AND NOT ((((VGA_Pixel_Buffer_avalon_pixel_dma_master_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter)))))))))) OR CPU_data_master_arbiterlock));
  --rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave : rdv_fifo_for_VGA_Pixel_Buffer_avalon_pixel_dma_master_to_SRAM_avalon_sram_slave_module
    port map(
      data_out => VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_output_from_SRAM_avalon_sram_slave,
      empty => open,
      fifo_contains_ones_n => VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_empty_SRAM_avalon_sram_slave,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave,
      read => SRAM_avalon_sram_slave_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT SRAM_avalon_sram_slave_waits_for_read;

  VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register <= NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_empty_SRAM_avalon_sram_slave;
  --local readdatavalid VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave <= ((SRAM_avalon_sram_slave_readdatavalid_from_sa AND VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_output_from_SRAM_avalon_sram_slave)) AND NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_rdv_fifo_empty_SRAM_avalon_sram_slave;
  --allow new arb cycle for SRAM/avalon_sram_slave, which is an e_assign
  SRAM_avalon_sram_slave_allow_new_arb_cycle <= NOT CPU_data_master_arbiterlock AND NOT ((VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock AND (saved_chosen_master_btw_VGA_Pixel_Buffer_avalon_pixel_dma_master_and_SRAM_avalon_sram_slave)));
  --VGA_Pixel_Buffer/avalon_pixel_dma_master assignment into master qualified-requests vector for SRAM/avalon_sram_slave, which is an e_assign
  SRAM_avalon_sram_slave_master_qreq_vector(0) <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave;
  --VGA_Pixel_Buffer/avalon_pixel_dma_master grant SRAM/avalon_sram_slave, which is an e_assign
  internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_grant_vector(0);
  --VGA_Pixel_Buffer/avalon_pixel_dma_master saved-grant SRAM/avalon_sram_slave, which is an e_assign
  VGA_Pixel_Buffer_avalon_pixel_dma_master_saved_grant_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_arb_winner(0) AND internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave;
  --saved chosen master btw VGA_Pixel_Buffer/avalon_pixel_dma_master and SRAM/avalon_sram_slave, which is an e_assign
  saved_chosen_master_btw_VGA_Pixel_Buffer_avalon_pixel_dma_master_and_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_saved_chosen_master_vector(0);
  --CPU/data_master assignment into master qualified-requests vector for SRAM/avalon_sram_slave, which is an e_assign
  SRAM_avalon_sram_slave_master_qreq_vector(1) <= internal_CPU_data_master_qualified_request_SRAM_avalon_sram_slave;
  --CPU/data_master grant SRAM/avalon_sram_slave, which is an e_assign
  internal_CPU_data_master_granted_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_grant_vector(1);
  --CPU/data_master saved-grant SRAM/avalon_sram_slave, which is an e_assign
  CPU_data_master_saved_grant_SRAM_avalon_sram_slave <= SRAM_avalon_sram_slave_arb_winner(1) AND internal_CPU_data_master_requests_SRAM_avalon_sram_slave;
  --SRAM/avalon_sram_slave chosen-master double-vector, which is an e_assign
  SRAM_avalon_sram_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((SRAM_avalon_sram_slave_master_qreq_vector & SRAM_avalon_sram_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT SRAM_avalon_sram_slave_master_qreq_vector & NOT SRAM_avalon_sram_slave_master_qreq_vector))) + (std_logic_vector'("000") & (SRAM_avalon_sram_slave_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  SRAM_avalon_sram_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((SRAM_avalon_sram_slave_allow_new_arb_cycle AND or_reduce(SRAM_avalon_sram_slave_grant_vector)))) = '1'), SRAM_avalon_sram_slave_grant_vector, SRAM_avalon_sram_slave_saved_chosen_master_vector);
  --saved SRAM_avalon_sram_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SRAM_avalon_sram_slave_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(SRAM_avalon_sram_slave_allow_new_arb_cycle) = '1' then 
        SRAM_avalon_sram_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(SRAM_avalon_sram_slave_grant_vector)) = '1'), SRAM_avalon_sram_slave_grant_vector, SRAM_avalon_sram_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  SRAM_avalon_sram_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((SRAM_avalon_sram_slave_chosen_master_double_vector(1) OR SRAM_avalon_sram_slave_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((SRAM_avalon_sram_slave_chosen_master_double_vector(0) OR SRAM_avalon_sram_slave_chosen_master_double_vector(2)))));
  --SRAM/avalon_sram_slave chosen master rotated left, which is an e_assign
  SRAM_avalon_sram_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(SRAM_avalon_sram_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(SRAM_avalon_sram_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --SRAM/avalon_sram_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SRAM_avalon_sram_slave_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(SRAM_avalon_sram_slave_grant_vector)) = '1' then 
        SRAM_avalon_sram_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(SRAM_avalon_sram_slave_end_xfer) = '1'), SRAM_avalon_sram_slave_chosen_master_rot_left, SRAM_avalon_sram_slave_grant_vector);
      end if;
    end if;

  end process;

  --~SRAM_avalon_sram_slave_reset assignment, which is an e_assign
  SRAM_avalon_sram_slave_reset <= NOT reset_n;
  --SRAM_avalon_sram_slave_firsttransfer first transaction, which is an e_assign
  SRAM_avalon_sram_slave_firsttransfer <= A_WE_StdLogic((std_logic'(SRAM_avalon_sram_slave_begins_xfer) = '1'), SRAM_avalon_sram_slave_unreg_firsttransfer, SRAM_avalon_sram_slave_reg_firsttransfer);
  --SRAM_avalon_sram_slave_unreg_firsttransfer first transaction, which is an e_assign
  SRAM_avalon_sram_slave_unreg_firsttransfer <= NOT ((SRAM_avalon_sram_slave_slavearbiterlockenable AND SRAM_avalon_sram_slave_any_continuerequest));
  --SRAM_avalon_sram_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      SRAM_avalon_sram_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(SRAM_avalon_sram_slave_begins_xfer) = '1' then 
        SRAM_avalon_sram_slave_reg_firsttransfer <= SRAM_avalon_sram_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --SRAM_avalon_sram_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  SRAM_avalon_sram_slave_beginbursttransfer_internal <= SRAM_avalon_sram_slave_begins_xfer;
  --SRAM_avalon_sram_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  SRAM_avalon_sram_slave_arbitration_holdoff_internal <= SRAM_avalon_sram_slave_begins_xfer AND SRAM_avalon_sram_slave_firsttransfer;
  --SRAM_avalon_sram_slave_read assignment, which is an e_mux
  SRAM_avalon_sram_slave_read <= ((internal_CPU_data_master_granted_SRAM_avalon_sram_slave AND CPU_data_master_read)) OR ((internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave AND VGA_Pixel_Buffer_avalon_pixel_dma_master_read));
  --SRAM_avalon_sram_slave_write assignment, which is an e_mux
  SRAM_avalon_sram_slave_write <= internal_CPU_data_master_granted_SRAM_avalon_sram_slave AND CPU_data_master_write;
  shifted_address_to_SRAM_avalon_sram_slave_from_CPU_data_master <= A_EXT (Std_Logic_Vector'(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(CPU_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 29);
  --SRAM_avalon_sram_slave_address mux, which is an e_mux
  SRAM_avalon_sram_slave_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SRAM_avalon_sram_slave)) = '1'), (std_logic_vector'("000") & ((A_SRL(shifted_address_to_SRAM_avalon_sram_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000001"))))), (A_SRL(shifted_address_to_SRAM_avalon_sram_slave_from_VGA_Pixel_Buffer_avalon_pixel_dma_master,std_logic_vector'("00000000000000000000000000000001")))), 18);
  shifted_address_to_SRAM_avalon_sram_slave_from_VGA_Pixel_Buffer_avalon_pixel_dma_master <= VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave;
  --d1_SRAM_avalon_sram_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_SRAM_avalon_sram_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_SRAM_avalon_sram_slave_end_xfer <= SRAM_avalon_sram_slave_end_xfer;
    end if;

  end process;

  --SRAM_avalon_sram_slave_waits_for_read in a cycle, which is an e_mux
  SRAM_avalon_sram_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(SRAM_avalon_sram_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --SRAM_avalon_sram_slave_in_a_read_cycle assignment, which is an e_assign
  SRAM_avalon_sram_slave_in_a_read_cycle <= ((internal_CPU_data_master_granted_SRAM_avalon_sram_slave AND CPU_data_master_read)) OR ((internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave AND VGA_Pixel_Buffer_avalon_pixel_dma_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= SRAM_avalon_sram_slave_in_a_read_cycle;
  --SRAM_avalon_sram_slave_waits_for_write in a cycle, which is an e_mux
  SRAM_avalon_sram_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(SRAM_avalon_sram_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --SRAM_avalon_sram_slave_in_a_write_cycle assignment, which is an e_assign
  SRAM_avalon_sram_slave_in_a_write_cycle <= internal_CPU_data_master_granted_SRAM_avalon_sram_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= SRAM_avalon_sram_slave_in_a_write_cycle;
  wait_for_SRAM_avalon_sram_slave_counter <= std_logic'('0');
  --SRAM_avalon_sram_slave_byteenable byte enable port mux, which is an e_mux
  SRAM_avalon_sram_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_SRAM_avalon_sram_slave)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_CPU_data_master_byteenable_SRAM_avalon_sram_slave)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_1(1), CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_1(0), CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_0(1), CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_0(0)) <= CPU_data_master_byteenable;
  internal_CPU_data_master_byteenable_SRAM_avalon_sram_slave <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_0, CPU_data_master_byteenable_SRAM_avalon_sram_slave_segment_1);
  --vhdl renameroo for output signals
  CPU_data_master_byteenable_SRAM_avalon_sram_slave <= internal_CPU_data_master_byteenable_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  CPU_data_master_granted_SRAM_avalon_sram_slave <= internal_CPU_data_master_granted_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_SRAM_avalon_sram_slave <= internal_CPU_data_master_qualified_request_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register <= internal_CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register;
  --vhdl renameroo for output signals
  CPU_data_master_requests_SRAM_avalon_sram_slave <= internal_CPU_data_master_requests_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave;
--synthesis translate_off
    --SRAM/avalon_sram_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_granted_SRAM_avalon_sram_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(CPU_data_master_saved_grant_SRAM_avalon_sram_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_pixel_dma_master_saved_grant_SRAM_avalon_sram_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Serial_Port_avalon_rs232_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Serial_Port_avalon_rs232_slave_irq : IN STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_address : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Serial_Port_avalon_rs232_slave_chipselect : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_irq_from_sa : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_read : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Serial_Port_avalon_rs232_slave_reset : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_write : OUT STD_LOGIC;
                 signal Serial_Port_avalon_rs232_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Serial_Port_avalon_rs232_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC
              );
end entity Serial_Port_avalon_rs232_slave_arbitrator;


architecture europa of Serial_Port_avalon_rs232_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_allgrants :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_any_continuerequest :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_arb_counter_enable :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_begins_xfer :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_end_xfer :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_firsttransfer :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_grant_vector :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_in_a_read_cycle :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_in_a_write_cycle :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_master_qreq_vector :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_reg_firsttransfer :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_waits_for_read :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Serial_Port_avalon_rs232_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Serial_Port_avalon_rs232_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Serial_Port_avalon_rs232_slave_end_xfer;
    end if;

  end process;

  Serial_Port_avalon_rs232_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave);
  --assign Serial_Port_avalon_rs232_slave_readdata_from_sa = Serial_Port_avalon_rs232_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Serial_Port_avalon_rs232_slave_readdata_from_sa <= Serial_Port_avalon_rs232_slave_readdata;
  internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("10000000000000001000000010000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave <= CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register_in;
  --Serial_Port_avalon_rs232_slave_arb_share_counter set values, which is an e_mux
  Serial_Port_avalon_rs232_slave_arb_share_set_values <= std_logic_vector'("001");
  --Serial_Port_avalon_rs232_slave_non_bursting_master_requests mux, which is an e_mux
  Serial_Port_avalon_rs232_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave;
  --Serial_Port_avalon_rs232_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Serial_Port_avalon_rs232_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Serial_Port_avalon_rs232_slave_arb_share_counter_next_value assignment, which is an e_assign
  Serial_Port_avalon_rs232_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Serial_Port_avalon_rs232_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Serial_Port_avalon_rs232_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Serial_Port_avalon_rs232_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Serial_Port_avalon_rs232_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Serial_Port_avalon_rs232_slave_allgrants all slave grants, which is an e_mux
  Serial_Port_avalon_rs232_slave_allgrants <= Serial_Port_avalon_rs232_slave_grant_vector;
  --Serial_Port_avalon_rs232_slave_end_xfer assignment, which is an e_assign
  Serial_Port_avalon_rs232_slave_end_xfer <= NOT ((Serial_Port_avalon_rs232_slave_waits_for_read OR Serial_Port_avalon_rs232_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave <= Serial_Port_avalon_rs232_slave_end_xfer AND (((NOT Serial_Port_avalon_rs232_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Serial_Port_avalon_rs232_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Serial_Port_avalon_rs232_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave AND Serial_Port_avalon_rs232_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave AND NOT Serial_Port_avalon_rs232_slave_non_bursting_master_requests));
  --Serial_Port_avalon_rs232_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Serial_Port_avalon_rs232_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Serial_Port_avalon_rs232_slave_arb_counter_enable) = '1' then 
        Serial_Port_avalon_rs232_slave_arb_share_counter <= Serial_Port_avalon_rs232_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Serial_Port_avalon_rs232_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Serial_Port_avalon_rs232_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Serial_Port_avalon_rs232_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave)) OR ((end_xfer_arb_share_counter_term_Serial_Port_avalon_rs232_slave AND NOT Serial_Port_avalon_rs232_slave_non_bursting_master_requests)))) = '1' then 
        Serial_Port_avalon_rs232_slave_slavearbiterlockenable <= or_reduce(Serial_Port_avalon_rs232_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Serial_Port/avalon_rs232_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Serial_Port_avalon_rs232_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Serial_Port_avalon_rs232_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Serial_Port_avalon_rs232_slave_slavearbiterlockenable2 <= or_reduce(Serial_Port_avalon_rs232_slave_arb_share_counter_next_value);
  --CPU/data_master Serial_Port/avalon_rs232_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Serial_Port_avalon_rs232_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Serial_Port_avalon_rs232_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Serial_Port_avalon_rs232_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register_in <= ((internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave AND CPU_data_master_read) AND NOT Serial_Port_avalon_rs232_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register <= p1_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave, which is an e_mux
  CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave <= CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave_shift_register;
  --Serial_Port_avalon_rs232_slave_writedata mux, which is an e_mux
  Serial_Port_avalon_rs232_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave;
  --CPU/data_master saved-grant Serial_Port/avalon_rs232_slave, which is an e_assign
  CPU_data_master_saved_grant_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave;
  --allow new arb cycle for Serial_Port/avalon_rs232_slave, which is an e_assign
  Serial_Port_avalon_rs232_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Serial_Port_avalon_rs232_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Serial_Port_avalon_rs232_slave_master_qreq_vector <= std_logic'('1');
  --~Serial_Port_avalon_rs232_slave_reset assignment, which is an e_assign
  Serial_Port_avalon_rs232_slave_reset <= NOT reset_n;
  Serial_Port_avalon_rs232_slave_chipselect <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave;
  --Serial_Port_avalon_rs232_slave_firsttransfer first transaction, which is an e_assign
  Serial_Port_avalon_rs232_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Serial_Port_avalon_rs232_slave_begins_xfer) = '1'), Serial_Port_avalon_rs232_slave_unreg_firsttransfer, Serial_Port_avalon_rs232_slave_reg_firsttransfer);
  --Serial_Port_avalon_rs232_slave_unreg_firsttransfer first transaction, which is an e_assign
  Serial_Port_avalon_rs232_slave_unreg_firsttransfer <= NOT ((Serial_Port_avalon_rs232_slave_slavearbiterlockenable AND Serial_Port_avalon_rs232_slave_any_continuerequest));
  --Serial_Port_avalon_rs232_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Serial_Port_avalon_rs232_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Serial_Port_avalon_rs232_slave_begins_xfer) = '1' then 
        Serial_Port_avalon_rs232_slave_reg_firsttransfer <= Serial_Port_avalon_rs232_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Serial_Port_avalon_rs232_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Serial_Port_avalon_rs232_slave_beginbursttransfer_internal <= Serial_Port_avalon_rs232_slave_begins_xfer;
  --Serial_Port_avalon_rs232_slave_read assignment, which is an e_mux
  Serial_Port_avalon_rs232_slave_read <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave AND CPU_data_master_read;
  --Serial_Port_avalon_rs232_slave_write assignment, which is an e_mux
  Serial_Port_avalon_rs232_slave_write <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave AND CPU_data_master_write;
  shifted_address_to_Serial_Port_avalon_rs232_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Serial_Port_avalon_rs232_slave_address mux, which is an e_mux
  Serial_Port_avalon_rs232_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_Serial_Port_avalon_rs232_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_Serial_Port_avalon_rs232_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Serial_Port_avalon_rs232_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Serial_Port_avalon_rs232_slave_end_xfer <= Serial_Port_avalon_rs232_slave_end_xfer;
    end if;

  end process;

  --Serial_Port_avalon_rs232_slave_waits_for_read in a cycle, which is an e_mux
  Serial_Port_avalon_rs232_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Serial_Port_avalon_rs232_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Serial_Port_avalon_rs232_slave_in_a_read_cycle assignment, which is an e_assign
  Serial_Port_avalon_rs232_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Serial_Port_avalon_rs232_slave_in_a_read_cycle;
  --Serial_Port_avalon_rs232_slave_waits_for_write in a cycle, which is an e_mux
  Serial_Port_avalon_rs232_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Serial_Port_avalon_rs232_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Serial_Port_avalon_rs232_slave_in_a_write_cycle assignment, which is an e_assign
  Serial_Port_avalon_rs232_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Serial_Port_avalon_rs232_slave_in_a_write_cycle;
  wait_for_Serial_Port_avalon_rs232_slave_counter <= std_logic'('0');
  --Serial_Port_avalon_rs232_slave_byteenable byte enable port mux, which is an e_mux
  Serial_Port_avalon_rs232_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign Serial_Port_avalon_rs232_slave_irq_from_sa = Serial_Port_avalon_rs232_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  Serial_Port_avalon_rs232_slave_irq_from_sa <= Serial_Port_avalon_rs232_slave_irq;
  --vhdl renameroo for output signals
  CPU_data_master_granted_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_granted_Serial_Port_avalon_rs232_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Serial_Port_avalon_rs232_slave <= internal_CPU_data_master_requests_Serial_Port_avalon_rs232_slave;
--synthesis translate_off
    --Serial_Port/avalon_rs232_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Slider_Switches_avalon_parallel_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Slider_Switches_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                 signal Slider_Switches_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal Slider_Switches_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Slider_Switches_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                 signal Slider_Switches_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                 signal Slider_Switches_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Slider_Switches_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                 signal Slider_Switches_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                 signal Slider_Switches_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Slider_Switches_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC
              );
end entity Slider_Switches_avalon_parallel_port_slave_arbitrator;


architecture europa of Slider_Switches_avalon_parallel_port_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_allgrants :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_any_continuerequest :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_arb_counter_enable :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_begins_xfer :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_firsttransfer :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_grant_vector :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_master_qreq_vector :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_waits_for_read :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_Slider_Switches_avalon_parallel_port_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_Slider_Switches_avalon_parallel_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Slider_Switches_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  Slider_Switches_avalon_parallel_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave);
  --assign Slider_Switches_avalon_parallel_port_slave_readdata_from_sa = Slider_Switches_avalon_parallel_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_readdata_from_sa <= Slider_Switches_avalon_parallel_port_slave_readdata;
  internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000000000001000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register_in;
  --Slider_Switches_avalon_parallel_port_slave_arb_share_counter set values, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_arb_share_set_values <= std_logic_vector'("001");
  --Slider_Switches_avalon_parallel_port_slave_non_bursting_master_requests mux, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave;
  --Slider_Switches_avalon_parallel_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Slider_Switches_avalon_parallel_port_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Slider_Switches_avalon_parallel_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Slider_Switches_avalon_parallel_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Slider_Switches_avalon_parallel_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Slider_Switches_avalon_parallel_port_slave_allgrants all slave grants, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_allgrants <= Slider_Switches_avalon_parallel_port_slave_grant_vector;
  --Slider_Switches_avalon_parallel_port_slave_end_xfer assignment, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_end_xfer <= NOT ((Slider_Switches_avalon_parallel_port_slave_waits_for_read OR Slider_Switches_avalon_parallel_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave <= Slider_Switches_avalon_parallel_port_slave_end_xfer AND (((NOT Slider_Switches_avalon_parallel_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Slider_Switches_avalon_parallel_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave AND Slider_Switches_avalon_parallel_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave AND NOT Slider_Switches_avalon_parallel_port_slave_non_bursting_master_requests));
  --Slider_Switches_avalon_parallel_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Slider_Switches_avalon_parallel_port_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Slider_Switches_avalon_parallel_port_slave_arb_counter_enable) = '1' then 
        Slider_Switches_avalon_parallel_port_slave_arb_share_counter <= Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Slider_Switches_avalon_parallel_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave)) OR ((end_xfer_arb_share_counter_term_Slider_Switches_avalon_parallel_port_slave AND NOT Slider_Switches_avalon_parallel_port_slave_non_bursting_master_requests)))) = '1' then 
        Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable <= or_reduce(Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master Slider_Switches/avalon_parallel_port_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable2 <= or_reduce(Slider_Switches_avalon_parallel_port_slave_arb_share_counter_next_value);
  --CPU/data_master Slider_Switches/avalon_parallel_port_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --Slider_Switches_avalon_parallel_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register_in <= ((internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_read) AND NOT Slider_Switches_avalon_parallel_port_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register <= p1_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave, which is an e_mux
  CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave <= CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave_shift_register;
  --Slider_Switches_avalon_parallel_port_slave_writedata mux, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave;
  --CPU/data_master saved-grant Slider_Switches/avalon_parallel_port_slave, which is an e_assign
  CPU_data_master_saved_grant_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave;
  --allow new arb cycle for Slider_Switches/avalon_parallel_port_slave, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Slider_Switches_avalon_parallel_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Slider_Switches_avalon_parallel_port_slave_master_qreq_vector <= std_logic'('1');
  --~Slider_Switches_avalon_parallel_port_slave_reset assignment, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_reset <= NOT reset_n;
  Slider_Switches_avalon_parallel_port_slave_chipselect <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave;
  --Slider_Switches_avalon_parallel_port_slave_firsttransfer first transaction, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(Slider_Switches_avalon_parallel_port_slave_begins_xfer) = '1'), Slider_Switches_avalon_parallel_port_slave_unreg_firsttransfer, Slider_Switches_avalon_parallel_port_slave_reg_firsttransfer);
  --Slider_Switches_avalon_parallel_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_unreg_firsttransfer <= NOT ((Slider_Switches_avalon_parallel_port_slave_slavearbiterlockenable AND Slider_Switches_avalon_parallel_port_slave_any_continuerequest));
  --Slider_Switches_avalon_parallel_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Slider_Switches_avalon_parallel_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Slider_Switches_avalon_parallel_port_slave_begins_xfer) = '1' then 
        Slider_Switches_avalon_parallel_port_slave_reg_firsttransfer <= Slider_Switches_avalon_parallel_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Slider_Switches_avalon_parallel_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_beginbursttransfer_internal <= Slider_Switches_avalon_parallel_port_slave_begins_xfer;
  --Slider_Switches_avalon_parallel_port_slave_read assignment, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_read <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_read;
  --Slider_Switches_avalon_parallel_port_slave_write assignment, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_write <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_write;
  shifted_address_to_Slider_Switches_avalon_parallel_port_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --Slider_Switches_avalon_parallel_port_slave_address mux, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_address <= A_EXT (A_SRL(shifted_address_to_Slider_Switches_avalon_parallel_port_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_Slider_Switches_avalon_parallel_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Slider_Switches_avalon_parallel_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Slider_Switches_avalon_parallel_port_slave_end_xfer <= Slider_Switches_avalon_parallel_port_slave_end_xfer;
    end if;

  end process;

  --Slider_Switches_avalon_parallel_port_slave_waits_for_read in a cycle, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Slider_Switches_avalon_parallel_port_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Slider_Switches_avalon_parallel_port_slave_in_a_read_cycle assignment, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_in_a_read_cycle <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Slider_Switches_avalon_parallel_port_slave_in_a_read_cycle;
  --Slider_Switches_avalon_parallel_port_slave_waits_for_write in a cycle, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(Slider_Switches_avalon_parallel_port_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --Slider_Switches_avalon_parallel_port_slave_in_a_write_cycle assignment, which is an e_assign
  Slider_Switches_avalon_parallel_port_slave_in_a_write_cycle <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Slider_Switches_avalon_parallel_port_slave_in_a_write_cycle;
  wait_for_Slider_Switches_avalon_parallel_port_slave_counter <= std_logic'('0');
  --Slider_Switches_avalon_parallel_port_slave_byteenable byte enable port mux, which is an e_mux
  Slider_Switches_avalon_parallel_port_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave <= internal_CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave;
--synthesis translate_off
    --Slider_Switches/avalon_parallel_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_byteenable : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_chipselect : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_read : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_write : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC
              );
end entity VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator;


architecture europa of VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_0 :  STD_LOGIC;
                signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_1 :  STD_LOGIC;
                signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_3 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_allgrants :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_any_continuerequest :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_arb_counter_enable :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_begins_xfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_grant_vector :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_in_a_read_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_in_a_write_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_master_qreq_vector :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_non_bursting_master_requests :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_reg_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_unreg_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_read :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register :  STD_LOGIC;
                signal wait_for_VGA_Char_Buffer_avalon_char_buffer_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer;
    end if;

  end process;

  VGA_Char_Buffer_avalon_char_buffer_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave);
  --assign VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa = VGA_Char_Buffer_avalon_char_buffer_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa <= VGA_Char_Buffer_avalon_char_buffer_slave_readdata;
  internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("01001000000000000000000000000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa = VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa <= VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest;
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave <= CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register_in;
  --VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter set values, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000001")), 3);
  --VGA_Char_Buffer_avalon_char_buffer_slave_non_bursting_master_requests mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave;
  --VGA_Char_Buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(VGA_Char_Buffer_avalon_char_buffer_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --VGA_Char_Buffer_avalon_char_buffer_slave_allgrants all slave grants, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_allgrants <= VGA_Char_Buffer_avalon_char_buffer_slave_grant_vector;
  --VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer <= NOT ((VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_read OR VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave <= VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer AND (((NOT VGA_Char_Buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter arbitration counter enable, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave AND VGA_Char_Buffer_avalon_char_buffer_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave AND NOT VGA_Char_Buffer_avalon_char_buffer_slave_non_bursting_master_requests));
  --VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Char_Buffer_avalon_char_buffer_slave_arb_counter_enable) = '1' then 
        VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter <= VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((VGA_Char_Buffer_avalon_char_buffer_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave)) OR ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_buffer_slave AND NOT VGA_Char_Buffer_avalon_char_buffer_slave_non_bursting_master_requests)))) = '1' then 
        VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable <= or_reduce(VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master VGA_Char_Buffer/avalon_char_buffer_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable2 <= or_reduce(VGA_Char_Buffer_avalon_char_buffer_slave_arb_share_counter_next_value);
  --CPU/data_master VGA_Char_Buffer/avalon_char_buffer_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --VGA_Char_Buffer_avalon_char_buffer_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register))) OR (((((NOT CPU_data_master_waitrequest OR CPU_data_master_no_byte_enables_and_last_term) OR NOT(internal_CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave))) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register_in <= ((internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_read) AND NOT VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register <= p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave <= CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave_shift_register;
  --VGA_Char_Buffer_avalon_char_buffer_slave_writedata mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_writedata <= CPU_data_master_dbs_write_8;
  --master is always granted when requested
  internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave;
  --CPU/data_master saved-grant VGA_Char_Buffer/avalon_char_buffer_slave, which is an e_assign
  CPU_data_master_saved_grant_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave;
  --allow new arb cycle for VGA_Char_Buffer/avalon_char_buffer_slave, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  VGA_Char_Buffer_avalon_char_buffer_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  VGA_Char_Buffer_avalon_char_buffer_slave_master_qreq_vector <= std_logic'('1');
  VGA_Char_Buffer_avalon_char_buffer_slave_chipselect <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave;
  --VGA_Char_Buffer_avalon_char_buffer_slave_firsttransfer first transaction, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_firsttransfer <= A_WE_StdLogic((std_logic'(VGA_Char_Buffer_avalon_char_buffer_slave_begins_xfer) = '1'), VGA_Char_Buffer_avalon_char_buffer_slave_unreg_firsttransfer, VGA_Char_Buffer_avalon_char_buffer_slave_reg_firsttransfer);
  --VGA_Char_Buffer_avalon_char_buffer_slave_unreg_firsttransfer first transaction, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_unreg_firsttransfer <= NOT ((VGA_Char_Buffer_avalon_char_buffer_slave_slavearbiterlockenable AND VGA_Char_Buffer_avalon_char_buffer_slave_any_continuerequest));
  --VGA_Char_Buffer_avalon_char_buffer_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_buffer_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Char_Buffer_avalon_char_buffer_slave_begins_xfer) = '1' then 
        VGA_Char_Buffer_avalon_char_buffer_slave_reg_firsttransfer <= VGA_Char_Buffer_avalon_char_buffer_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_buffer_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_beginbursttransfer_internal <= VGA_Char_Buffer_avalon_char_buffer_slave_begins_xfer;
  --VGA_Char_Buffer_avalon_char_buffer_slave_read assignment, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_read <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_read;
  --VGA_Char_Buffer_avalon_char_buffer_slave_write assignment, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_write <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_write;
  --VGA_Char_Buffer_avalon_char_buffer_slave_address mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_address <= A_EXT (Std_Logic_Vector'(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & CPU_data_master_dbs_address(1 DOWNTO 0)), 13);
  --d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer <= VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_read in a cycle, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_read <= VGA_Char_Buffer_avalon_char_buffer_slave_in_a_read_cycle AND internal_VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa;
  --VGA_Char_Buffer_avalon_char_buffer_slave_in_a_read_cycle assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_in_a_read_cycle <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= VGA_Char_Buffer_avalon_char_buffer_slave_in_a_read_cycle;
  --VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_write in a cycle, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_waits_for_write <= VGA_Char_Buffer_avalon_char_buffer_slave_in_a_write_cycle AND internal_VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa;
  --VGA_Char_Buffer_avalon_char_buffer_slave_in_a_write_cycle assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_buffer_slave_in_a_write_cycle <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= VGA_Char_Buffer_avalon_char_buffer_slave_in_a_write_cycle;
  wait_for_VGA_Char_Buffer_avalon_char_buffer_slave_counter <= std_logic'('0');
  --VGA_Char_Buffer_avalon_char_buffer_slave_byteenable byte enable port mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_buffer_slave_byteenable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_3, CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_2, CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_1, CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_0) <= CPU_data_master_byteenable;
  internal_CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_2, CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave_segment_3)));
  --vhdl renameroo for output signals
  CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa <= internal_VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa;
--synthesis translate_off
    --VGA_Char_Buffer/avalon_char_buffer_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Char_Buffer_avalon_char_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_address : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_control_slave_chipselect : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_read : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_control_slave_reset : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_write : OUT STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC
              );
end entity VGA_Char_Buffer_avalon_char_control_slave_arbitrator;


architecture europa of VGA_Char_Buffer_avalon_char_control_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_allgrants :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_any_continuerequest :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_arb_counter_enable :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_begins_xfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_end_xfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_grant_vector :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_master_qreq_vector :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_waits_for_read :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_VGA_Char_Buffer_avalon_char_control_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_VGA_Char_Buffer_avalon_char_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT VGA_Char_Buffer_avalon_char_control_slave_end_xfer;
    end if;

  end process;

  VGA_Char_Buffer_avalon_char_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave);
  --assign VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa = VGA_Char_Buffer_avalon_char_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa <= VGA_Char_Buffer_avalon_char_control_slave_readdata;
  internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("10000000000000011000000110000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave <= CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register_in;
  --VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter set values, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_arb_share_set_values <= std_logic_vector'("001");
  --VGA_Char_Buffer_avalon_char_control_slave_non_bursting_master_requests mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave;
  --VGA_Char_Buffer_avalon_char_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(VGA_Char_Buffer_avalon_char_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Char_Buffer_avalon_char_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --VGA_Char_Buffer_avalon_char_control_slave_allgrants all slave grants, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_allgrants <= VGA_Char_Buffer_avalon_char_control_slave_grant_vector;
  --VGA_Char_Buffer_avalon_char_control_slave_end_xfer assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_end_xfer <= NOT ((VGA_Char_Buffer_avalon_char_control_slave_waits_for_read OR VGA_Char_Buffer_avalon_char_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave <= VGA_Char_Buffer_avalon_char_control_slave_end_xfer AND (((NOT VGA_Char_Buffer_avalon_char_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave AND VGA_Char_Buffer_avalon_char_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave AND NOT VGA_Char_Buffer_avalon_char_control_slave_non_bursting_master_requests));
  --VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Char_Buffer_avalon_char_control_slave_arb_counter_enable) = '1' then 
        VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter <= VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((VGA_Char_Buffer_avalon_char_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave)) OR ((end_xfer_arb_share_counter_term_VGA_Char_Buffer_avalon_char_control_slave AND NOT VGA_Char_Buffer_avalon_char_control_slave_non_bursting_master_requests)))) = '1' then 
        VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable <= or_reduce(VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master VGA_Char_Buffer/avalon_char_control_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable2 <= or_reduce(VGA_Char_Buffer_avalon_char_control_slave_arb_share_counter_next_value);
  --CPU/data_master VGA_Char_Buffer/avalon_char_control_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --VGA_Char_Buffer_avalon_char_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register_in <= ((internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_read) AND NOT VGA_Char_Buffer_avalon_char_control_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register <= p1_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave <= CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave_shift_register;
  --VGA_Char_Buffer_avalon_char_control_slave_writedata mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave;
  --CPU/data_master saved-grant VGA_Char_Buffer/avalon_char_control_slave, which is an e_assign
  CPU_data_master_saved_grant_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave;
  --allow new arb cycle for VGA_Char_Buffer/avalon_char_control_slave, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  VGA_Char_Buffer_avalon_char_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  VGA_Char_Buffer_avalon_char_control_slave_master_qreq_vector <= std_logic'('1');
  --~VGA_Char_Buffer_avalon_char_control_slave_reset assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_reset <= NOT reset_n;
  VGA_Char_Buffer_avalon_char_control_slave_chipselect <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave;
  --VGA_Char_Buffer_avalon_char_control_slave_firsttransfer first transaction, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(VGA_Char_Buffer_avalon_char_control_slave_begins_xfer) = '1'), VGA_Char_Buffer_avalon_char_control_slave_unreg_firsttransfer, VGA_Char_Buffer_avalon_char_control_slave_reg_firsttransfer);
  --VGA_Char_Buffer_avalon_char_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_unreg_firsttransfer <= NOT ((VGA_Char_Buffer_avalon_char_control_slave_slavearbiterlockenable AND VGA_Char_Buffer_avalon_char_control_slave_any_continuerequest));
  --VGA_Char_Buffer_avalon_char_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Char_Buffer_avalon_char_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Char_Buffer_avalon_char_control_slave_begins_xfer) = '1' then 
        VGA_Char_Buffer_avalon_char_control_slave_reg_firsttransfer <= VGA_Char_Buffer_avalon_char_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_beginbursttransfer_internal <= VGA_Char_Buffer_avalon_char_control_slave_begins_xfer;
  --VGA_Char_Buffer_avalon_char_control_slave_read assignment, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_read <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_read;
  --VGA_Char_Buffer_avalon_char_control_slave_write assignment, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_write <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_write;
  shifted_address_to_VGA_Char_Buffer_avalon_char_control_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --VGA_Char_Buffer_avalon_char_control_slave_address mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_VGA_Char_Buffer_avalon_char_control_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer <= VGA_Char_Buffer_avalon_char_control_slave_end_xfer;
    end if;

  end process;

  --VGA_Char_Buffer_avalon_char_control_slave_waits_for_read in a cycle, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Char_Buffer_avalon_char_control_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --VGA_Char_Buffer_avalon_char_control_slave_in_a_read_cycle assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_in_a_read_cycle <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= VGA_Char_Buffer_avalon_char_control_slave_in_a_read_cycle;
  --VGA_Char_Buffer_avalon_char_control_slave_waits_for_write in a cycle, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Char_Buffer_avalon_char_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --VGA_Char_Buffer_avalon_char_control_slave_in_a_write_cycle assignment, which is an e_assign
  VGA_Char_Buffer_avalon_char_control_slave_in_a_write_cycle <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= VGA_Char_Buffer_avalon_char_control_slave_in_a_write_cycle;
  wait_for_VGA_Char_Buffer_avalon_char_control_slave_counter <= std_logic'('0');
  --VGA_Char_Buffer_avalon_char_control_slave_byteenable byte enable port mux, which is an e_mux
  VGA_Char_Buffer_avalon_char_control_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave <= internal_CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave;
--synthesis translate_off
    --VGA_Char_Buffer/avalon_char_control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Char_Buffer_avalon_char_source_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_foreground_sink_ready_from_sa : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal VGA_Char_Buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Char_Buffer_avalon_char_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Char_Buffer_avalon_char_source_ready : OUT STD_LOGIC
              );
end entity VGA_Char_Buffer_avalon_char_source_arbitrator;


architecture europa of VGA_Char_Buffer_avalon_char_source_arbitrator is

begin

  --mux VGA_Char_Buffer_avalon_char_source_ready, which is an e_mux
  VGA_Char_Buffer_avalon_char_source_ready <= Alpha_Blending_avalon_foreground_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Controller_avalon_vga_sink_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Controller_avalon_vga_sink_ready : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Controller_avalon_vga_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Controller_avalon_vga_sink_endofpacket : OUT STD_LOGIC;
                 signal VGA_Controller_avalon_vga_sink_ready_from_sa : OUT STD_LOGIC;
                 signal VGA_Controller_avalon_vga_sink_reset : OUT STD_LOGIC;
                 signal VGA_Controller_avalon_vga_sink_startofpacket : OUT STD_LOGIC;
                 signal VGA_Controller_avalon_vga_sink_valid : OUT STD_LOGIC
              );
end entity VGA_Controller_avalon_vga_sink_arbitrator;


architecture europa of VGA_Controller_avalon_vga_sink_arbitrator is

begin

  --mux VGA_Controller_avalon_vga_sink_data, which is an e_mux
  VGA_Controller_avalon_vga_sink_data <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data;
  --mux VGA_Controller_avalon_vga_sink_endofpacket, which is an e_mux
  VGA_Controller_avalon_vga_sink_endofpacket <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket;
  --assign VGA_Controller_avalon_vga_sink_ready_from_sa = VGA_Controller_avalon_vga_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Controller_avalon_vga_sink_ready_from_sa <= VGA_Controller_avalon_vga_sink_ready;
  --mux VGA_Controller_avalon_vga_sink_startofpacket, which is an e_mux
  VGA_Controller_avalon_vga_sink_startofpacket <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket;
  --mux VGA_Controller_avalon_vga_sink_valid, which is an e_mux
  VGA_Controller_avalon_vga_sink_valid <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid;
  --~VGA_Controller_avalon_vga_sink_reset assignment, which is an e_assign
  VGA_Controller_avalon_vga_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal Alpha_Blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                 signal Alpha_Blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                 signal Alpha_Blending_avalon_blended_source_valid : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket : OUT STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa : OUT STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket : OUT STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid : OUT STD_LOGIC
              );
end entity VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator;


architecture europa of VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator is

begin

  --mux VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data, which is an e_mux
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data <= Alpha_Blending_avalon_blended_source_data;
  --mux VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket, which is an e_mux
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket <= Alpha_Blending_avalon_blended_source_endofpacket;
  --assign VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa = VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa <= VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready;
  --mux VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket, which is an e_mux
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket <= Alpha_Blending_avalon_blended_source_startofpacket;
  --mux VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid, which is an e_mux
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid <= Alpha_Blending_avalon_blended_source_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Controller_avalon_vga_sink_ready_from_sa : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready : OUT STD_LOGIC
              );
end entity VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator;


architecture europa of VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator is

begin

  --mux VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready, which is an e_mux
  VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready <= VGA_Controller_avalon_vga_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_Buffer_avalon_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_control_slave_read : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_control_slave_write : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC
              );
end entity VGA_Pixel_Buffer_avalon_control_slave_arbitrator;


architecture europa of VGA_Pixel_Buffer_avalon_control_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register_in :  STD_LOGIC;
                signal CPU_data_master_saved_grant_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_allgrants :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_any_continuerequest :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_arb_counter_enable :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_begins_xfer :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_end_xfer :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_firsttransfer :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_grant_vector :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_master_qreq_vector :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_waits_for_read :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal p1_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_VGA_Pixel_Buffer_avalon_control_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal wait_for_VGA_Pixel_Buffer_avalon_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT VGA_Pixel_Buffer_avalon_control_slave_end_xfer;
    end if;

  end process;

  VGA_Pixel_Buffer_avalon_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave);
  --assign VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa = VGA_Pixel_Buffer_avalon_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa <= VGA_Pixel_Buffer_avalon_control_slave_readdata;
  internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10000000000000011000000100000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --registered rdv signal_name registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave assignment, which is an e_assign
  registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave <= CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register_in;
  --VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter set values, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_arb_share_set_values <= std_logic_vector'("001");
  --VGA_Pixel_Buffer_avalon_control_slave_non_bursting_master_requests mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave;
  --VGA_Pixel_Buffer_avalon_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(VGA_Pixel_Buffer_avalon_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Pixel_Buffer_avalon_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --VGA_Pixel_Buffer_avalon_control_slave_allgrants all slave grants, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_allgrants <= VGA_Pixel_Buffer_avalon_control_slave_grant_vector;
  --VGA_Pixel_Buffer_avalon_control_slave_end_xfer assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_end_xfer <= NOT ((VGA_Pixel_Buffer_avalon_control_slave_waits_for_read OR VGA_Pixel_Buffer_avalon_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave <= VGA_Pixel_Buffer_avalon_control_slave_end_xfer AND (((NOT VGA_Pixel_Buffer_avalon_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave AND VGA_Pixel_Buffer_avalon_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave AND NOT VGA_Pixel_Buffer_avalon_control_slave_non_bursting_master_requests));
  --VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Pixel_Buffer_avalon_control_slave_arb_counter_enable) = '1' then 
        VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter <= VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((VGA_Pixel_Buffer_avalon_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave)) OR ((end_xfer_arb_share_counter_term_VGA_Pixel_Buffer_avalon_control_slave AND NOT VGA_Pixel_Buffer_avalon_control_slave_non_bursting_master_requests)))) = '1' then 
        VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable <= or_reduce(VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master VGA_Pixel_Buffer/avalon_control_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable2 <= or_reduce(VGA_Pixel_Buffer_avalon_control_slave_arb_share_counter_next_value);
  --CPU/data_master VGA_Pixel_Buffer/avalon_control_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --VGA_Pixel_Buffer_avalon_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave AND NOT ((((CPU_data_master_read AND (CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register))) OR (((NOT CPU_data_master_waitrequest) AND CPU_data_master_write))));
  --CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register_in <= ((internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_read) AND NOT VGA_Pixel_Buffer_avalon_control_slave_waits_for_read) AND NOT (CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register);
  --shift register p1 CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register) & A_ToStdLogicVector(CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register_in)));
  --CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register <= p1_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register;
    end if;

  end process;

  --local readdatavalid CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave, which is an e_mux
  CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave <= CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave_shift_register;
  --VGA_Pixel_Buffer_avalon_control_slave_writedata mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_writedata <= CPU_data_master_writedata;
  --master is always granted when requested
  internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave;
  --CPU/data_master saved-grant VGA_Pixel_Buffer/avalon_control_slave, which is an e_assign
  CPU_data_master_saved_grant_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave;
  --allow new arb cycle for VGA_Pixel_Buffer/avalon_control_slave, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  VGA_Pixel_Buffer_avalon_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  VGA_Pixel_Buffer_avalon_control_slave_master_qreq_vector <= std_logic'('1');
  --VGA_Pixel_Buffer_avalon_control_slave_firsttransfer first transaction, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(VGA_Pixel_Buffer_avalon_control_slave_begins_xfer) = '1'), VGA_Pixel_Buffer_avalon_control_slave_unreg_firsttransfer, VGA_Pixel_Buffer_avalon_control_slave_reg_firsttransfer);
  --VGA_Pixel_Buffer_avalon_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_unreg_firsttransfer <= NOT ((VGA_Pixel_Buffer_avalon_control_slave_slavearbiterlockenable AND VGA_Pixel_Buffer_avalon_control_slave_any_continuerequest));
  --VGA_Pixel_Buffer_avalon_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Pixel_Buffer_avalon_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(VGA_Pixel_Buffer_avalon_control_slave_begins_xfer) = '1' then 
        VGA_Pixel_Buffer_avalon_control_slave_reg_firsttransfer <= VGA_Pixel_Buffer_avalon_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --VGA_Pixel_Buffer_avalon_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_beginbursttransfer_internal <= VGA_Pixel_Buffer_avalon_control_slave_begins_xfer;
  --VGA_Pixel_Buffer_avalon_control_slave_read assignment, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_read <= internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_read;
  --VGA_Pixel_Buffer_avalon_control_slave_write assignment, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_write <= internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_write;
  shifted_address_to_VGA_Pixel_Buffer_avalon_control_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --VGA_Pixel_Buffer_avalon_control_slave_address mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_address <= A_EXT (A_SRL(shifted_address_to_VGA_Pixel_Buffer_avalon_control_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer <= VGA_Pixel_Buffer_avalon_control_slave_end_xfer;
    end if;

  end process;

  --VGA_Pixel_Buffer_avalon_control_slave_waits_for_read in a cycle, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_control_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --VGA_Pixel_Buffer_avalon_control_slave_in_a_read_cycle assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_in_a_read_cycle <= internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= VGA_Pixel_Buffer_avalon_control_slave_in_a_read_cycle;
  --VGA_Pixel_Buffer_avalon_control_slave_waits_for_write in a cycle, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --VGA_Pixel_Buffer_avalon_control_slave_in_a_write_cycle assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_control_slave_in_a_write_cycle <= internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= VGA_Pixel_Buffer_avalon_control_slave_in_a_write_cycle;
  wait_for_VGA_Pixel_Buffer_avalon_control_slave_counter <= std_logic'('0');
  --VGA_Pixel_Buffer_avalon_control_slave_byteenable byte enable port mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_control_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (CPU_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave <= internal_CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave;
--synthesis translate_off
    --VGA_Pixel_Buffer/avalon_control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator is 
        port (
              -- inputs:
                 signal SRAM_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal d1_SRAM_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_reset : OUT STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest : OUT STD_LOGIC
              );
end entity VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator;


architecture europa of VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator is
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_is_granted_some_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_but_no_slave_selected :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_last_time :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_run :  STD_LOGIC;
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter :  STD_LOGIC;
                signal internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter :  STD_LOGIC;
                signal pre_flush_VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave OR NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave OR NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave OR NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_read)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(VGA_Pixel_Buffer_avalon_pixel_dma_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_pixel_dma_master_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000100000000") & VGA_Pixel_Buffer_avalon_pixel_dma_master_address(18 DOWNTO 0));
  --VGA_Pixel_Buffer_avalon_pixel_dma_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_but_no_slave_selected <= (VGA_Pixel_Buffer_avalon_pixel_dma_master_read AND VGA_Pixel_Buffer_avalon_pixel_dma_master_run) AND NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_dma_master_is_granted_some_slave <= VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid <= VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave;
  --latent slave read data valid which is not flushed, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid <= VGA_Pixel_Buffer_avalon_pixel_dma_master_read_but_no_slave_selected OR pre_flush_VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid;
  --VGA_Pixel_Buffer/avalon_pixel_dma_master readdata mux, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata <= SRAM_avalon_sram_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest <= NOT VGA_Pixel_Buffer_avalon_pixel_dma_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter <= p1_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((VGA_Pixel_Buffer_avalon_pixel_dma_master_run AND VGA_Pixel_Buffer_avalon_pixel_dma_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --~VGA_Pixel_Buffer_avalon_pixel_dma_master_reset assignment, which is an e_assign
  VGA_Pixel_Buffer_avalon_pixel_dma_master_reset <= NOT reset_n;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter;
  --vhdl renameroo for output signals
  VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest;
--synthesis translate_off
    --VGA_Pixel_Buffer_avalon_pixel_dma_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        VGA_Pixel_Buffer_avalon_pixel_dma_master_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        VGA_Pixel_Buffer_avalon_pixel_dma_master_address_last_time <= VGA_Pixel_Buffer_avalon_pixel_dma_master_address;
      end if;

    end process;

    --VGA_Pixel_Buffer/avalon_pixel_dma_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest AND (VGA_Pixel_Buffer_avalon_pixel_dma_master_read);
      end if;

    end process;

    --VGA_Pixel_Buffer_avalon_pixel_dma_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((VGA_Pixel_Buffer_avalon_pixel_dma_master_address /= VGA_Pixel_Buffer_avalon_pixel_dma_master_address_last_time))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("VGA_Pixel_Buffer_avalon_pixel_dma_master_address did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --VGA_Pixel_Buffer_avalon_pixel_dma_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        VGA_Pixel_Buffer_avalon_pixel_dma_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        VGA_Pixel_Buffer_avalon_pixel_dma_master_read_last_time <= VGA_Pixel_Buffer_avalon_pixel_dma_master_read;
      end if;

    end process;

    --VGA_Pixel_Buffer_avalon_pixel_dma_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(VGA_Pixel_Buffer_avalon_pixel_dma_master_read) /= std_logic'(VGA_Pixel_Buffer_avalon_pixel_dma_master_read_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("VGA_Pixel_Buffer_avalon_pixel_dma_master_read did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_Buffer_avalon_pixel_source_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Pixel_Buffer_avalon_pixel_source_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_source_valid : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_Buffer_avalon_pixel_source_ready : OUT STD_LOGIC
              );
end entity VGA_Pixel_Buffer_avalon_pixel_source_arbitrator;


architecture europa of VGA_Pixel_Buffer_avalon_pixel_source_arbitrator is

begin

  --mux VGA_Pixel_Buffer_avalon_pixel_source_ready, which is an e_mux
  VGA_Pixel_Buffer_avalon_pixel_source_ready <= VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Pixel_Buffer_avalon_pixel_source_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_Buffer_avalon_pixel_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Buffer_avalon_pixel_source_valid : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket : OUT STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa : OUT STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset : OUT STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket : OUT STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid : OUT STD_LOGIC
              );
end entity VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator;


architecture europa of VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator is

begin

  --mux VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data, which is an e_mux
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data <= VGA_Pixel_Buffer_avalon_pixel_source_data;
  --mux VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket, which is an e_mux
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket <= VGA_Pixel_Buffer_avalon_pixel_source_endofpacket;
  --assign VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa = VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa <= VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready;
  --mux VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket, which is an e_mux
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket <= VGA_Pixel_Buffer_avalon_pixel_source_startofpacket;
  --mux VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid, which is an e_mux
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid <= VGA_Pixel_Buffer_avalon_pixel_source_valid;
  --~VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset assignment, which is an e_assign
  VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready : OUT STD_LOGIC
              );
end entity VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator;


architecture europa of VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator is

begin

  --mux VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready, which is an e_mux
  VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready <= VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator is 
        port (
              -- inputs:
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_ready : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket : OUT STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa : OUT STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_reset : OUT STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket : OUT STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_sink_valid : OUT STD_LOGIC
              );
end entity VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator;


architecture europa of VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator is

begin

  --mux VGA_Pixel_Scaler_avalon_scaler_sink_data, which is an e_mux
  VGA_Pixel_Scaler_avalon_scaler_sink_data <= VGA_Pixel_RGB_Resampler_avalon_rgb_source_data;
  --mux VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket, which is an e_mux
  VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket <= VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket;
  --assign VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa = VGA_Pixel_Scaler_avalon_scaler_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa <= VGA_Pixel_Scaler_avalon_scaler_sink_ready;
  --mux VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket, which is an e_mux
  VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket <= VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket;
  --mux VGA_Pixel_Scaler_avalon_scaler_sink_valid, which is an e_mux
  VGA_Pixel_Scaler_avalon_scaler_sink_valid <= VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid;
  --~VGA_Pixel_Scaler_avalon_scaler_sink_reset assignment, which is an e_assign
  VGA_Pixel_Scaler_avalon_scaler_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGA_Pixel_Scaler_avalon_scaler_source_arbitrator is 
        port (
              -- inputs:
                 signal Alpha_Blending_avalon_background_sink_ready_from_sa : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal VGA_Pixel_Scaler_avalon_scaler_source_endofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_startofpacket : IN STD_LOGIC;
                 signal VGA_Pixel_Scaler_avalon_scaler_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal VGA_Pixel_Scaler_avalon_scaler_source_ready : OUT STD_LOGIC
              );
end entity VGA_Pixel_Scaler_avalon_scaler_source_arbitrator;


architecture europa of VGA_Pixel_Scaler_avalon_scaler_source_arbitrator is

begin

  --mux VGA_Pixel_Scaler_avalon_scaler_source_ready, which is an e_mux
  VGA_Pixel_Scaler_avalon_scaler_source_ready <= Alpha_Blending_avalon_background_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios_system_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_waitrequest : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal nios_system_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal nios_system_clock_0_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios_system_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal CPU_data_master_byteenable_nios_system_clock_0_in : OUT STD_LOGIC;
                 signal CPU_data_master_granted_nios_system_clock_0_in : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_nios_system_clock_0_in : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_nios_system_clock_0_in : OUT STD_LOGIC;
                 signal CPU_data_master_requests_nios_system_clock_0_in : OUT STD_LOGIC;
                 signal d1_nios_system_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_address : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_nativeaddress : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_read : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios_system_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_write : OUT STD_LOGIC;
                 signal nios_system_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios_system_clock_0_in_arbitrator;


architecture europa of nios_system_clock_0_in_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_nios_system_clock_0_in_segment_0 :  STD_LOGIC;
                signal CPU_data_master_byteenable_nios_system_clock_0_in_segment_1 :  STD_LOGIC;
                signal CPU_data_master_byteenable_nios_system_clock_0_in_segment_2 :  STD_LOGIC;
                signal CPU_data_master_byteenable_nios_system_clock_0_in_segment_3 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_nios_system_clock_0_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios_system_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_byteenable_nios_system_clock_0_in :  STD_LOGIC;
                signal internal_CPU_data_master_granted_nios_system_clock_0_in :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_nios_system_clock_0_in :  STD_LOGIC;
                signal internal_CPU_data_master_requests_nios_system_clock_0_in :  STD_LOGIC;
                signal internal_nios_system_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios_system_clock_0_in_allgrants :  STD_LOGIC;
                signal nios_system_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios_system_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios_system_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal nios_system_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal nios_system_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios_system_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios_system_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios_system_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios_system_clock_0_in_begins_xfer :  STD_LOGIC;
                signal nios_system_clock_0_in_end_xfer :  STD_LOGIC;
                signal nios_system_clock_0_in_firsttransfer :  STD_LOGIC;
                signal nios_system_clock_0_in_grant_vector :  STD_LOGIC;
                signal nios_system_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal nios_system_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal nios_system_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal nios_system_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios_system_clock_0_in_pretend_byte_enable :  STD_LOGIC;
                signal nios_system_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal nios_system_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios_system_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios_system_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios_system_clock_0_in_waits_for_read :  STD_LOGIC;
                signal nios_system_clock_0_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios_system_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios_system_clock_0_in_end_xfer;
    end if;

  end process;

  nios_system_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_nios_system_clock_0_in);
  --assign nios_system_clock_0_in_readdata_from_sa = nios_system_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios_system_clock_0_in_readdata_from_sa <= nios_system_clock_0_in_readdata;
  internal_CPU_data_master_requests_nios_system_clock_0_in <= to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 1) & A_ToStdLogicVector(std_logic'('0'))) = std_logic_vector'("10000000000000010000000110000")))) AND ((CPU_data_master_read OR CPU_data_master_write));
  --assign nios_system_clock_0_in_waitrequest_from_sa = nios_system_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios_system_clock_0_in_waitrequest_from_sa <= nios_system_clock_0_in_waitrequest;
  --nios_system_clock_0_in_arb_share_counter set values, which is an e_mux
  nios_system_clock_0_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_nios_system_clock_0_in)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000001")), 3);
  --nios_system_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  nios_system_clock_0_in_non_bursting_master_requests <= internal_CPU_data_master_requests_nios_system_clock_0_in;
  --nios_system_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios_system_clock_0_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios_system_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  nios_system_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios_system_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (nios_system_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios_system_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (nios_system_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --nios_system_clock_0_in_allgrants all slave grants, which is an e_mux
  nios_system_clock_0_in_allgrants <= nios_system_clock_0_in_grant_vector;
  --nios_system_clock_0_in_end_xfer assignment, which is an e_assign
  nios_system_clock_0_in_end_xfer <= NOT ((nios_system_clock_0_in_waits_for_read OR nios_system_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios_system_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios_system_clock_0_in <= nios_system_clock_0_in_end_xfer AND (((NOT nios_system_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios_system_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios_system_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios_system_clock_0_in AND nios_system_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios_system_clock_0_in AND NOT nios_system_clock_0_in_non_bursting_master_requests));
  --nios_system_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios_system_clock_0_in_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios_system_clock_0_in_arb_counter_enable) = '1' then 
        nios_system_clock_0_in_arb_share_counter <= nios_system_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios_system_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios_system_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios_system_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios_system_clock_0_in)) OR ((end_xfer_arb_share_counter_term_nios_system_clock_0_in AND NOT nios_system_clock_0_in_non_bursting_master_requests)))) = '1' then 
        nios_system_clock_0_in_slavearbiterlockenable <= or_reduce(nios_system_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master nios_system_clock_0/in arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= nios_system_clock_0_in_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --nios_system_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios_system_clock_0_in_slavearbiterlockenable2 <= or_reduce(nios_system_clock_0_in_arb_share_counter_next_value);
  --CPU/data_master nios_system_clock_0/in arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= nios_system_clock_0_in_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --nios_system_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios_system_clock_0_in_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_nios_system_clock_0_in <= internal_CPU_data_master_requests_nios_system_clock_0_in AND NOT ((((CPU_data_master_read AND (NOT CPU_data_master_waitrequest))) OR (((((NOT CPU_data_master_waitrequest OR CPU_data_master_no_byte_enables_and_last_term) OR NOT(internal_CPU_data_master_byteenable_nios_system_clock_0_in))) AND CPU_data_master_write))));
  --nios_system_clock_0_in_writedata mux, which is an e_mux
  nios_system_clock_0_in_writedata <= CPU_data_master_dbs_write_8;
  --assign nios_system_clock_0_in_endofpacket_from_sa = nios_system_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios_system_clock_0_in_endofpacket_from_sa <= nios_system_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_CPU_data_master_granted_nios_system_clock_0_in <= internal_CPU_data_master_qualified_request_nios_system_clock_0_in;
  --CPU/data_master saved-grant nios_system_clock_0/in, which is an e_assign
  CPU_data_master_saved_grant_nios_system_clock_0_in <= internal_CPU_data_master_requests_nios_system_clock_0_in;
  --allow new arb cycle for nios_system_clock_0/in, which is an e_assign
  nios_system_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios_system_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios_system_clock_0_in_master_qreq_vector <= std_logic'('1');
  --nios_system_clock_0_in_reset_n assignment, which is an e_assign
  nios_system_clock_0_in_reset_n <= reset_n;
  --nios_system_clock_0_in_firsttransfer first transaction, which is an e_assign
  nios_system_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios_system_clock_0_in_begins_xfer) = '1'), nios_system_clock_0_in_unreg_firsttransfer, nios_system_clock_0_in_reg_firsttransfer);
  --nios_system_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  nios_system_clock_0_in_unreg_firsttransfer <= NOT ((nios_system_clock_0_in_slavearbiterlockenable AND nios_system_clock_0_in_any_continuerequest));
  --nios_system_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios_system_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios_system_clock_0_in_begins_xfer) = '1' then 
        nios_system_clock_0_in_reg_firsttransfer <= nios_system_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios_system_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios_system_clock_0_in_beginbursttransfer_internal <= nios_system_clock_0_in_begins_xfer;
  --nios_system_clock_0_in_read assignment, which is an e_mux
  nios_system_clock_0_in_read <= internal_CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_read;
  --nios_system_clock_0_in_write assignment, which is an e_mux
  nios_system_clock_0_in_write <= ((internal_CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_write)) AND nios_system_clock_0_in_pretend_byte_enable;
  --nios_system_clock_0_in_address mux, which is an e_mux
  nios_system_clock_0_in_address <= Vector_To_Std_Logic(Std_Logic_Vector'(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & CPU_data_master_dbs_address(1 DOWNTO 0)));
  --slaveid nios_system_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  nios_system_clock_0_in_nativeaddress <= Vector_To_Std_Logic(A_SRL(CPU_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")));
  --d1_nios_system_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios_system_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios_system_clock_0_in_end_xfer <= nios_system_clock_0_in_end_xfer;
    end if;

  end process;

  --nios_system_clock_0_in_waits_for_read in a cycle, which is an e_mux
  nios_system_clock_0_in_waits_for_read <= nios_system_clock_0_in_in_a_read_cycle AND internal_nios_system_clock_0_in_waitrequest_from_sa;
  --nios_system_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  nios_system_clock_0_in_in_a_read_cycle <= internal_CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios_system_clock_0_in_in_a_read_cycle;
  --nios_system_clock_0_in_waits_for_write in a cycle, which is an e_mux
  nios_system_clock_0_in_waits_for_write <= nios_system_clock_0_in_in_a_write_cycle AND internal_nios_system_clock_0_in_waitrequest_from_sa;
  --nios_system_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  nios_system_clock_0_in_in_a_write_cycle <= internal_CPU_data_master_granted_nios_system_clock_0_in AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios_system_clock_0_in_in_a_write_cycle;
  wait_for_nios_system_clock_0_in_counter <= std_logic'('0');
  --nios_system_clock_0_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios_system_clock_0_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_CPU_data_master_granted_nios_system_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_CPU_data_master_byteenable_nios_system_clock_0_in))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (CPU_data_master_byteenable_nios_system_clock_0_in_segment_3, CPU_data_master_byteenable_nios_system_clock_0_in_segment_2, CPU_data_master_byteenable_nios_system_clock_0_in_segment_1, CPU_data_master_byteenable_nios_system_clock_0_in_segment_0) <= CPU_data_master_byteenable;
  internal_CPU_data_master_byteenable_nios_system_clock_0_in <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), CPU_data_master_byteenable_nios_system_clock_0_in_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), CPU_data_master_byteenable_nios_system_clock_0_in_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (CPU_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), CPU_data_master_byteenable_nios_system_clock_0_in_segment_2, CPU_data_master_byteenable_nios_system_clock_0_in_segment_3)));
  --vhdl renameroo for output signals
  CPU_data_master_byteenable_nios_system_clock_0_in <= internal_CPU_data_master_byteenable_nios_system_clock_0_in;
  --vhdl renameroo for output signals
  CPU_data_master_granted_nios_system_clock_0_in <= internal_CPU_data_master_granted_nios_system_clock_0_in;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_nios_system_clock_0_in <= internal_CPU_data_master_qualified_request_nios_system_clock_0_in;
  --vhdl renameroo for output signals
  CPU_data_master_requests_nios_system_clock_0_in <= internal_CPU_data_master_requests_nios_system_clock_0_in;
  --vhdl renameroo for output signals
  nios_system_clock_0_in_waitrequest_from_sa <= internal_nios_system_clock_0_in_waitrequest_from_sa;
--synthesis translate_off
    --nios_system_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios_system_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal External_Clocks_avalon_clocks_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_External_Clocks_avalon_clocks_slave_end_xfer : IN STD_LOGIC;
                 signal nios_system_clock_0_out_address : IN STD_LOGIC;
                 signal nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                 signal nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                 signal nios_system_clock_0_out_read : IN STD_LOGIC;
                 signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                 signal nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                 signal nios_system_clock_0_out_write : IN STD_LOGIC;
                 signal nios_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios_system_clock_0_out_address_to_slave : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios_system_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal nios_system_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity nios_system_clock_0_out_arbitrator;


architecture europa of nios_system_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios_system_clock_0_out_address_to_slave :  STD_LOGIC;
                signal internal_nios_system_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios_system_clock_0_out_address_last_time :  STD_LOGIC;
                signal nios_system_clock_0_out_read_last_time :  STD_LOGIC;
                signal nios_system_clock_0_out_run :  STD_LOGIC;
                signal nios_system_clock_0_out_write_last_time :  STD_LOGIC;
                signal nios_system_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave OR nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave) OR NOT nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave OR NOT nios_system_clock_0_out_read) OR ((nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave AND nios_system_clock_0_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave OR NOT ((nios_system_clock_0_out_read OR nios_system_clock_0_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios_system_clock_0_out_read OR nios_system_clock_0_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios_system_clock_0_out_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios_system_clock_0_out_address_to_slave <= nios_system_clock_0_out_address;
  --nios_system_clock_0/out readdata mux, which is an e_mux
  nios_system_clock_0_out_readdata <= External_Clocks_avalon_clocks_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios_system_clock_0_out_waitrequest <= NOT nios_system_clock_0_out_run;
  --nios_system_clock_0_out_reset_n assignment, which is an e_assign
  nios_system_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios_system_clock_0_out_address_to_slave <= internal_nios_system_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  nios_system_clock_0_out_waitrequest <= internal_nios_system_clock_0_out_waitrequest;
--synthesis translate_off
    --nios_system_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios_system_clock_0_out_address_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios_system_clock_0_out_address_last_time <= nios_system_clock_0_out_address;
      end if;

    end process;

    --nios_system_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios_system_clock_0_out_waitrequest AND ((nios_system_clock_0_out_read OR nios_system_clock_0_out_write));
      end if;

    end process;

    --nios_system_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios_system_clock_0_out_address) /= std_logic'(nios_system_clock_0_out_address_last_time)))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("nios_system_clock_0_out_address did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios_system_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios_system_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios_system_clock_0_out_read_last_time <= nios_system_clock_0_out_read;
      end if;

    end process;

    --nios_system_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios_system_clock_0_out_read) /= std_logic'(nios_system_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("nios_system_clock_0_out_read did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios_system_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios_system_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios_system_clock_0_out_write_last_time <= nios_system_clock_0_out_write;
      end if;

    end process;

    --nios_system_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios_system_clock_0_out_write) /= std_logic'(nios_system_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("nios_system_clock_0_out_write did not heed wait!!!"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios_system_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios_system_clock_0_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios_system_clock_0_out_writedata_last_time <= nios_system_clock_0_out_writedata;
      end if;

    end process;

    --nios_system_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios_system_clock_0_out_writedata /= nios_system_clock_0_out_writedata_last_time)))) AND nios_system_clock_0_out_write)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("nios_system_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal CPU_data_master_read : IN STD_LOGIC;
                 signal CPU_data_master_write : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal CPU_data_master_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal CPU_data_master_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal CPU_data_master_arbiterlock :  STD_LOGIC;
                signal CPU_data_master_arbiterlock2 :  STD_LOGIC;
                signal CPU_data_master_continuerequest :  STD_LOGIC;
                signal CPU_data_master_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_CPU_data_master_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_CPU_data_master_requests_sysid_control_slave :  STD_LOGIC;
                signal shifted_address_to_sysid_control_slave_from_CPU_data_master :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC;
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC;
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_CPU_data_master_qualified_request_sysid_control_slave);
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_CPU_data_master_requests_sysid_control_slave <= ((to_std_logic(((Std_Logic_Vector'(CPU_data_master_address_to_slave(28 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("10000000000000010000000100000")))) AND ((CPU_data_master_read OR CPU_data_master_write)))) AND CPU_data_master_read;
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= std_logic_vector'("001");
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= internal_CPU_data_master_requests_sysid_control_slave;
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sysid_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sysid_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sysid_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= sysid_control_slave_grant_vector;
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysid_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= or_reduce(sysid_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --CPU/data_master sysid/control_slave arbiterlock, which is an e_assign
  CPU_data_master_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND CPU_data_master_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= or_reduce(sysid_control_slave_arb_share_counter_next_value);
  --CPU/data_master sysid/control_slave arbiterlock2, which is an e_assign
  CPU_data_master_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND CPU_data_master_continuerequest;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  sysid_control_slave_any_continuerequest <= std_logic'('1');
  --CPU_data_master_continuerequest continued request, which is an e_assign
  CPU_data_master_continuerequest <= std_logic'('1');
  internal_CPU_data_master_qualified_request_sysid_control_slave <= internal_CPU_data_master_requests_sysid_control_slave;
  --master is always granted when requested
  internal_CPU_data_master_granted_sysid_control_slave <= internal_CPU_data_master_qualified_request_sysid_control_slave;
  --CPU/data_master saved-grant sysid/control_slave, which is an e_assign
  CPU_data_master_saved_grant_sysid_control_slave <= internal_CPU_data_master_requests_sysid_control_slave;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysid_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysid_control_slave_master_qreq_vector <= std_logic'('1');
  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  shifted_address_to_sysid_control_slave_from_CPU_data_master <= CPU_data_master_address_to_slave;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_sysid_control_slave_from_CPU_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= internal_CPU_data_master_granted_sysid_control_slave AND CPU_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= internal_CPU_data_master_granted_sysid_control_slave AND CPU_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  CPU_data_master_granted_sysid_control_slave <= internal_CPU_data_master_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_qualified_request_sysid_control_slave <= internal_CPU_data_master_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  CPU_data_master_requests_sysid_control_slave <= internal_CPU_data_master_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios_system_reset_sys_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios_system_reset_sys_clk_domain_synch_module;


architecture europa of nios_system_reset_sys_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios_system_reset_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios_system_reset_clk_domain_synch_module;


architecture europa of nios_system_reset_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios_system_reset_vga_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios_system_reset_vga_clk_domain_synch_module;


architecture europa of nios_system_reset_vga_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios_system is 
        port (
              -- 1) global signals:
                 signal audio_clk : OUT STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal clk_27 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_clk : OUT STD_LOGIC;
                 signal sys_clk : OUT STD_LOGIC;
                 signal vga_clk : OUT STD_LOGIC;

              -- the_AV_Config
                 signal I2C_SCLK_from_the_AV_Config : OUT STD_LOGIC;
                 signal I2C_SDAT_to_and_from_the_AV_Config : INOUT STD_LOGIC;

              -- the_Audio
                 signal AUD_ADCDAT_to_the_Audio : IN STD_LOGIC;
                 signal AUD_ADCLRCK_to_and_from_the_Audio : INOUT STD_LOGIC;
                 signal AUD_BCLK_to_and_from_the_Audio : INOUT STD_LOGIC;
                 signal AUD_DACDAT_from_the_Audio : OUT STD_LOGIC;
                 signal AUD_DACLRCK_to_and_from_the_Audio : INOUT STD_LOGIC;

              -- the_Char_LCD_16x2
                 signal LCD_BLON_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                 signal LCD_DATA_to_and_from_the_Char_LCD_16x2 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal LCD_EN_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                 signal LCD_ON_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                 signal LCD_RS_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                 signal LCD_RW_from_the_Char_LCD_16x2 : OUT STD_LOGIC;

              -- the_Expansion_JP1
                 signal GPIO_0_to_and_from_the_Expansion_JP1 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- the_Expansion_JP2
                 signal GPIO_1_to_and_from_the_Expansion_JP2 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- the_Green_LEDs
                 signal LEDG_from_the_Green_LEDs : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);

              -- the_HEX3_HEX0
                 signal HEX0_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX1_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX2_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX3_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);

              -- the_HEX7_HEX4
                 signal HEX4_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX5_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX6_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal HEX7_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);

              -- the_PS2_Port
                 signal PS2_CLK_to_and_from_the_PS2_Port : INOUT STD_LOGIC;
                 signal PS2_DAT_to_and_from_the_PS2_Port : INOUT STD_LOGIC;

              -- the_Pushbuttons
                 signal KEY_to_the_Pushbuttons : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_Red_LEDs
                 signal LEDR_from_the_Red_LEDs : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);

              -- the_SDRAM
                 signal zs_addr_from_the_SDRAM : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_SDRAM : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_SDRAM : OUT STD_LOGIC;
                 signal zs_cke_from_the_SDRAM : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_SDRAM : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_SDRAM : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_SDRAM : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_SDRAM : OUT STD_LOGIC;
                 signal zs_we_n_from_the_SDRAM : OUT STD_LOGIC;

              -- the_SRAM
                 signal SRAM_ADDR_from_the_SRAM : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal SRAM_CE_N_from_the_SRAM : OUT STD_LOGIC;
                 signal SRAM_DQ_to_and_from_the_SRAM : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SRAM_LB_N_from_the_SRAM : OUT STD_LOGIC;
                 signal SRAM_OE_N_from_the_SRAM : OUT STD_LOGIC;
                 signal SRAM_UB_N_from_the_SRAM : OUT STD_LOGIC;
                 signal SRAM_WE_N_from_the_SRAM : OUT STD_LOGIC;

              -- the_Serial_Port
                 signal UART_RXD_to_the_Serial_Port : IN STD_LOGIC;
                 signal UART_TXD_from_the_Serial_Port : OUT STD_LOGIC;

              -- the_Slider_Switches
                 signal SW_to_the_Slider_Switches : IN STD_LOGIC_VECTOR (17 DOWNTO 0);

              -- the_VGA_Controller
                 signal VGA_BLANK_from_the_VGA_Controller : OUT STD_LOGIC;
                 signal VGA_B_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_CLK_from_the_VGA_Controller : OUT STD_LOGIC;
                 signal VGA_G_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_HS_from_the_VGA_Controller : OUT STD_LOGIC;
                 signal VGA_R_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_SYNC_from_the_VGA_Controller : OUT STD_LOGIC;
                 signal VGA_VS_from_the_VGA_Controller : OUT STD_LOGIC
              );
end entity nios_system;


architecture europa of nios_system is
component AV_Config_avalon_av_config_slave_arbitrator is 
           port (
                 -- inputs:
                    signal AV_Config_avalon_av_config_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal AV_Config_avalon_av_config_slave_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal AV_Config_avalon_av_config_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal AV_Config_avalon_av_config_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal AV_Config_avalon_av_config_slave_read : OUT STD_LOGIC;
                    signal AV_Config_avalon_av_config_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal AV_Config_avalon_av_config_slave_reset : OUT STD_LOGIC;
                    signal AV_Config_avalon_av_config_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal AV_Config_avalon_av_config_slave_write : OUT STD_LOGIC;
                    signal AV_Config_avalon_av_config_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_granted_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_AV_Config_avalon_av_config_slave : OUT STD_LOGIC;
                    signal d1_AV_Config_avalon_av_config_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : OUT STD_LOGIC
                 );
end component AV_Config_avalon_av_config_slave_arbitrator;

component AV_Config is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal I2C_SCLK : OUT STD_LOGIC;
                    signal I2C_SDAT : INOUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component AV_Config;

component Alpha_Blending_avalon_background_sink_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_background_sink_ready : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Pixel_Scaler_avalon_scaler_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Alpha_Blending_avalon_background_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal Alpha_Blending_avalon_background_sink_endofpacket : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_background_sink_ready_from_sa : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_background_sink_startofpacket : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_background_sink_valid : OUT STD_LOGIC
                 );
end component Alpha_Blending_avalon_background_sink_arbitrator;

component Alpha_Blending_avalon_foreground_sink_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_foreground_sink_ready : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Alpha_Blending_avalon_foreground_sink_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal Alpha_Blending_avalon_foreground_sink_endofpacket : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_foreground_sink_ready_from_sa : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_foreground_sink_reset : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_foreground_sink_startofpacket : OUT STD_LOGIC;
                    signal Alpha_Blending_avalon_foreground_sink_valid : OUT STD_LOGIC
                 );
end component Alpha_Blending_avalon_foreground_sink_arbitrator;

component Alpha_Blending_avalon_blended_source_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal Alpha_Blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                    signal Alpha_Blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                    signal Alpha_Blending_avalon_blended_source_valid : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Alpha_Blending_avalon_blended_source_ready : OUT STD_LOGIC
                 );
end component Alpha_Blending_avalon_blended_source_arbitrator;

component Alpha_Blending is 
           port (
                 -- inputs:
                    signal background_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal background_endofpacket : IN STD_LOGIC;
                    signal background_startofpacket : IN STD_LOGIC;
                    signal background_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal foreground_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal foreground_endofpacket : IN STD_LOGIC;
                    signal foreground_startofpacket : IN STD_LOGIC;
                    signal foreground_valid : IN STD_LOGIC;
                    signal output_ready : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;

                 -- outputs:
                    signal background_ready : OUT STD_LOGIC;
                    signal foreground_ready : OUT STD_LOGIC;
                    signal output_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal output_endofpacket : OUT STD_LOGIC;
                    signal output_startofpacket : OUT STD_LOGIC;
                    signal output_valid : OUT STD_LOGIC
                 );
end component Alpha_Blending;

component Audio_avalon_audio_slave_arbitrator is 
           port (
                 -- inputs:
                    signal Audio_avalon_audio_slave_irq : IN STD_LOGIC;
                    signal Audio_avalon_audio_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Audio_avalon_audio_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Audio_avalon_audio_slave_chipselect : OUT STD_LOGIC;
                    signal Audio_avalon_audio_slave_irq_from_sa : OUT STD_LOGIC;
                    signal Audio_avalon_audio_slave_read : OUT STD_LOGIC;
                    signal Audio_avalon_audio_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Audio_avalon_audio_slave_reset : OUT STD_LOGIC;
                    signal Audio_avalon_audio_slave_write : OUT STD_LOGIC;
                    signal Audio_avalon_audio_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_granted_Audio_avalon_audio_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Audio_avalon_audio_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Audio_avalon_audio_slave : OUT STD_LOGIC;
                    signal d1_Audio_avalon_audio_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave : OUT STD_LOGIC
                 );
end component Audio_avalon_audio_slave_arbitrator;

component Audio is 
           port (
                 -- inputs:
                    signal AUD_ADCDAT : IN STD_LOGIC;
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal AUD_ADCLRCK : INOUT STD_LOGIC;
                    signal AUD_BCLK : INOUT STD_LOGIC;
                    signal AUD_DACDAT : OUT STD_LOGIC;
                    signal AUD_DACLRCK : INOUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Audio;

component CPU_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_debugaccess : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal CPU_instruction_master_latency_counter : IN STD_LOGIC;
                    signal CPU_instruction_master_read : IN STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                    signal CPU_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_data_master_requests_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_instruction_master_granted_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_instruction_master_qualified_request_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_instruction_master_requests_CPU_jtag_debug_module : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal CPU_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_write : OUT STD_LOGIC;
                    signal CPU_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_CPU_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component CPU_jtag_debug_module_arbitrator;

component CPU_custom_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_custom_instruction_master_multi_start : IN STD_LOGIC;
                    signal CPU_fpoint_s1_done_from_sa : IN STD_LOGIC;
                    signal CPU_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_custom_instruction_master_multi_done : OUT STD_LOGIC;
                    signal CPU_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_custom_instruction_master_reset_n : OUT STD_LOGIC;
                    signal CPU_custom_instruction_master_start_CPU_fpoint_s1 : OUT STD_LOGIC;
                    signal CPU_fpoint_s1_select : OUT STD_LOGIC
                 );
end component CPU_custom_instruction_master_arbitrator;

component CPU_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal AV_Config_avalon_av_config_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal AV_Config_avalon_av_config_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal Audio_avalon_audio_slave_irq_from_sa : IN STD_LOGIC;
                    signal Audio_avalon_audio_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_address : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                    signal CPU_data_master_byteenable_SDRAM_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_byteenable_SRAM_avalon_sram_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal CPU_data_master_byteenable_nios_system_clock_0_in : IN STD_LOGIC;
                    signal CPU_data_master_granted_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Audio_avalon_audio_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Interval_Timer_s1 : IN STD_LOGIC;
                    signal CPU_data_master_granted_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_data_master_granted_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_granted_nios_system_clock_0_in : IN STD_LOGIC;
                    signal CPU_data_master_granted_sysid_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Audio_avalon_audio_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Interval_Timer_s1 : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_nios_system_clock_0_in : IN STD_LOGIC;
                    signal CPU_data_master_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Interval_Timer_s1 : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_nios_system_clock_0_in : IN STD_LOGIC;
                    signal CPU_data_master_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Audio_avalon_audio_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Interval_Timer_s1 : IN STD_LOGIC;
                    signal CPU_data_master_requests_JTAG_UART_avalon_jtag_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_data_master_requests_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_requests_nios_system_clock_0_in : IN STD_LOGIC;
                    signal CPU_data_master_requests_sysid_control_slave : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Expansion_JP2_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Green_LEDs_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Interval_Timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal Interval_Timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal JTAG_UART_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal JTAG_UART_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_irq_from_sa : IN STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal PS2_Port_avalon_ps2_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_irq_from_sa : IN STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Red_LEDs_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal SDRAM_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SDRAM_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal SRAM_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal Serial_Port_avalon_rs232_slave_irq_from_sa : IN STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Slider_Switches_avalon_parallel_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_AV_Config_avalon_av_config_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Audio_avalon_audio_slave_end_xfer : IN STD_LOGIC;
                    signal d1_CPU_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Green_LEDs_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Interval_Timer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_JTAG_UART_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_PS2_Port_avalon_ps2_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Pushbuttons_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Red_LEDs_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_SDRAM_s1_end_xfer : IN STD_LOGIC;
                    signal d1_SRAM_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Serial_Port_avalon_rs232_slave_end_xfer : IN STD_LOGIC;
                    signal d1_Slider_Switches_avalon_parallel_port_slave_end_xfer : IN STD_LOGIC;
                    signal d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer : IN STD_LOGIC;
                    signal d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_nios_system_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal nios_system_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios_system_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal CPU_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal CPU_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal CPU_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                    signal CPU_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_data_master_waitrequest : OUT STD_LOGIC
                 );
end component CPU_data_master_arbitrator;

component CPU_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal CPU_instruction_master_granted_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_instruction_master_granted_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_instruction_master_qualified_request_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_instruction_master_qualified_request_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_instruction_master_read : IN STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : IN STD_LOGIC;
                    signal CPU_instruction_master_requests_CPU_jtag_debug_module : IN STD_LOGIC;
                    signal CPU_instruction_master_requests_SDRAM_s1 : IN STD_LOGIC;
                    signal CPU_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal SDRAM_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SDRAM_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal d1_CPU_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_SDRAM_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal CPU_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_instruction_master_latency_counter : OUT STD_LOGIC;
                    signal CPU_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal CPU_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component CPU_instruction_master_arbitrator;

component CPU is 
           port (
                 -- inputs:
                    signal M_ci_multi_done : IN STD_LOGIC;
                    signal M_ci_multi_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal M_ci_multi_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal M_ci_multi_b : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal M_ci_multi_c : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal M_ci_multi_clk_en : OUT STD_LOGIC;
                    signal M_ci_multi_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal M_ci_multi_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal M_ci_multi_estatus : OUT STD_LOGIC;
                    signal M_ci_multi_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal M_ci_multi_n : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal M_ci_multi_readra : OUT STD_LOGIC;
                    signal M_ci_multi_readrb : OUT STD_LOGIC;
                    signal M_ci_multi_start : OUT STD_LOGIC;
                    signal M_ci_multi_status : OUT STD_LOGIC;
                    signal M_ci_multi_writerc : OUT STD_LOGIC;
                    signal d_address : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component CPU;

component CPU_fpoint_s1_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                    signal CPU_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal CPU_custom_instruction_master_start_CPU_fpoint_s1 : IN STD_LOGIC;
                    signal CPU_fpoint_s1_done : IN STD_LOGIC;
                    signal CPU_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_fpoint_s1_select : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_fpoint_s1_clk_en : OUT STD_LOGIC;
                    signal CPU_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                    signal CPU_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_fpoint_s1_reset : OUT STD_LOGIC;
                    signal CPU_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CPU_fpoint_s1_start : OUT STD_LOGIC
                 );
end component CPU_fpoint_s1_arbitrator;

component CPU_fpoint is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clk_en : IN STD_LOGIC;
                    signal dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal start : IN STD_LOGIC;

                 -- outputs:
                    signal done : OUT STD_LOGIC;
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component CPU_fpoint;

component Char_LCD_16x2_avalon_lcd_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal Char_LCD_16x2_avalon_lcd_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                    signal CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_address : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_chipselect : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_read : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal Char_LCD_16x2_avalon_lcd_slave_reset : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_write : OUT STD_LOGIC;
                    signal Char_LCD_16x2_avalon_lcd_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer : OUT STD_LOGIC
                 );
end component Char_LCD_16x2_avalon_lcd_slave_arbitrator;

component Char_LCD_16x2 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal LCD_BLON : OUT STD_LOGIC;
                    signal LCD_DATA : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal LCD_EN : OUT STD_LOGIC;
                    signal LCD_ON : OUT STD_LOGIC;
                    signal LCD_RS : OUT STD_LOGIC;
                    signal LCD_RW : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component Char_LCD_16x2;

component Expansion_JP1_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Expansion_JP1_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Expansion_JP1_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Expansion_JP1_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Expansion_JP1_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Expansion_JP1_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Expansion_JP1_avalon_parallel_port_slave_arbitrator;

component Expansion_JP1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal GPIO_0 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Expansion_JP1;

component Expansion_JP2_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Expansion_JP2_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Expansion_JP2_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Expansion_JP2_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Expansion_JP2_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Expansion_JP2_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Expansion_JP2_avalon_parallel_port_slave_arbitrator;

component Expansion_JP2 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal GPIO_1 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Expansion_JP2;

component External_Clocks_avalon_clocks_slave_arbitrator is 
           port (
                 -- inputs:
                    signal External_Clocks_avalon_clocks_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal nios_system_clock_0_out_address_to_slave : IN STD_LOGIC;
                    signal nios_system_clock_0_out_read : IN STD_LOGIC;
                    signal nios_system_clock_0_out_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal External_Clocks_avalon_clocks_slave_address : OUT STD_LOGIC;
                    signal External_Clocks_avalon_clocks_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal d1_External_Clocks_avalon_clocks_slave_end_xfer : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave : OUT STD_LOGIC
                 );
end component External_Clocks_avalon_clocks_slave_arbitrator;

component External_Clocks is 
           port (
                 -- inputs:
                    signal CLOCK_27 : IN STD_LOGIC;
                    signal CLOCK_50 : IN STD_LOGIC;
                    signal address : IN STD_LOGIC;

                 -- outputs:
                    signal AUD_CLK : OUT STD_LOGIC;
                    signal SDRAM_CLK : OUT STD_LOGIC;
                    signal VGA_CLK : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal sys_clk : OUT STD_LOGIC
                 );
end component External_Clocks;

component Green_LEDs_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Green_LEDs_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Green_LEDs_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Green_LEDs_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Green_LEDs_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Green_LEDs_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Green_LEDs_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Green_LEDs_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Green_LEDs_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Green_LEDs_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Green_LEDs_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Green_LEDs_avalon_parallel_port_slave_arbitrator;

component Green_LEDs is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal LEDG : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Green_LEDs;

component HEX3_HEX0_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX3_HEX0_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal HEX3_HEX0_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal HEX3_HEX0_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal HEX3_HEX0_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal HEX3_HEX0_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX3_HEX0_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal HEX3_HEX0_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal HEX3_HEX0_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component HEX3_HEX0_avalon_parallel_port_slave_arbitrator;

component HEX3_HEX0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX1 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX2 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX3 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component HEX3_HEX0;

component HEX7_HEX4_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX7_HEX4_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal HEX7_HEX4_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal HEX7_HEX4_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal HEX7_HEX4_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal HEX7_HEX4_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal HEX7_HEX4_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal HEX7_HEX4_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal HEX7_HEX4_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component HEX7_HEX4_avalon_parallel_port_slave_arbitrator;

component HEX7_HEX4 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX5 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX6 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX7 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component HEX7_HEX4;

component Interval_Timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Interval_Timer_s1_irq : IN STD_LOGIC;
                    signal Interval_Timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Interval_Timer_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Interval_Timer_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Interval_Timer_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Interval_Timer_s1 : OUT STD_LOGIC;
                    signal Interval_Timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal Interval_Timer_s1_chipselect : OUT STD_LOGIC;
                    signal Interval_Timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal Interval_Timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal Interval_Timer_s1_reset_n : OUT STD_LOGIC;
                    signal Interval_Timer_s1_write_n : OUT STD_LOGIC;
                    signal Interval_Timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_Interval_Timer_s1_end_xfer : OUT STD_LOGIC
                 );
end component Interval_Timer_s1_arbitrator;

component Interval_Timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component Interval_Timer;

component JTAG_UART_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal JTAG_UART_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal JTAG_UART_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_JTAG_UART_avalon_jtag_slave : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal JTAG_UART_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal JTAG_UART_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_JTAG_UART_avalon_jtag_slave_end_xfer : OUT STD_LOGIC
                 );
end component JTAG_UART_avalon_jtag_slave_arbitrator;

component JTAG_UART is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component JTAG_UART;

component PS2_Port_avalon_ps2_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal PS2_Port_avalon_ps2_slave_irq : IN STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal PS2_Port_avalon_ps2_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_address : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal PS2_Port_avalon_ps2_slave_chipselect : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_irq_from_sa : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_read : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal PS2_Port_avalon_ps2_slave_reset : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_write : OUT STD_LOGIC;
                    signal PS2_Port_avalon_ps2_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_PS2_Port_avalon_ps2_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave : OUT STD_LOGIC
                 );
end component PS2_Port_avalon_ps2_slave_arbitrator;

component PS2_Port is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal PS2_CLK : INOUT STD_LOGIC;
                    signal PS2_DAT : INOUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component PS2_Port;

component Pushbuttons_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Pushbuttons_avalon_parallel_port_slave_irq : IN STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Pushbuttons_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Pushbuttons_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_irq_from_sa : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Pushbuttons_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Pushbuttons_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Pushbuttons_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Pushbuttons_avalon_parallel_port_slave_arbitrator;

component Pushbuttons is 
           port (
                 -- inputs:
                    signal KEY : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Pushbuttons;

component Red_LEDs_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Red_LEDs_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Red_LEDs_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Red_LEDs_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Red_LEDs_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Red_LEDs_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Red_LEDs_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Red_LEDs_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Red_LEDs_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Red_LEDs_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Red_LEDs_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Red_LEDs_avalon_parallel_port_slave_arbitrator;

component Red_LEDs is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal LEDR : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Red_LEDs;

component SDRAM_s1_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal CPU_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_instruction_master_latency_counter : IN STD_LOGIC;
                    signal CPU_instruction_master_read : IN STD_LOGIC;
                    signal SDRAM_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SDRAM_s1_readdatavalid : IN STD_LOGIC;
                    signal SDRAM_s1_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_byteenable_SDRAM_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_granted_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SDRAM_s1_shift_register : OUT STD_LOGIC;
                    signal CPU_data_master_requests_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_instruction_master_granted_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_instruction_master_qualified_request_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_SDRAM_s1 : OUT STD_LOGIC;
                    signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register : OUT STD_LOGIC;
                    signal CPU_instruction_master_requests_SDRAM_s1 : OUT STD_LOGIC;
                    signal SDRAM_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal SDRAM_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal SDRAM_s1_chipselect : OUT STD_LOGIC;
                    signal SDRAM_s1_read_n : OUT STD_LOGIC;
                    signal SDRAM_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SDRAM_s1_reset_n : OUT STD_LOGIC;
                    signal SDRAM_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal SDRAM_s1_write_n : OUT STD_LOGIC;
                    signal SDRAM_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_SDRAM_s1_end_xfer : OUT STD_LOGIC
                 );
end component SDRAM_s1_arbitrator;

component SDRAM is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component SDRAM;

component SRAM_avalon_sram_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal SRAM_avalon_sram_slave_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_avalon_sram_slave_readdatavalid : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_byteenable_SRAM_avalon_sram_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_granted_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : OUT STD_LOGIC;
                    signal CPU_data_master_requests_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal SRAM_avalon_sram_slave_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal SRAM_avalon_sram_slave_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal SRAM_avalon_sram_slave_read : OUT STD_LOGIC;
                    signal SRAM_avalon_sram_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_avalon_sram_slave_reset : OUT STD_LOGIC;
                    signal SRAM_avalon_sram_slave_write : OUT STD_LOGIC;
                    signal SRAM_avalon_sram_slave_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave : OUT STD_LOGIC;
                    signal d1_SRAM_avalon_sram_slave_end_xfer : OUT STD_LOGIC
                 );
end component SRAM_avalon_sram_slave_arbitrator;

component SRAM is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal SRAM_ADDR : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal SRAM_CE_N : OUT STD_LOGIC;
                    signal SRAM_DQ : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_LB_N : OUT STD_LOGIC;
                    signal SRAM_OE_N : OUT STD_LOGIC;
                    signal SRAM_UB_N : OUT STD_LOGIC;
                    signal SRAM_WE_N : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdatavalid : OUT STD_LOGIC
                 );
end component SRAM;

component Serial_Port_avalon_rs232_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Serial_Port_avalon_rs232_slave_irq : IN STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_address : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Serial_Port_avalon_rs232_slave_chipselect : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_irq_from_sa : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_read : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Serial_Port_avalon_rs232_slave_reset : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_write : OUT STD_LOGIC;
                    signal Serial_Port_avalon_rs232_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Serial_Port_avalon_rs232_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave : OUT STD_LOGIC
                 );
end component Serial_Port_avalon_rs232_slave_arbitrator;

component Serial_Port is 
           port (
                 -- inputs:
                    signal UART_RXD : IN STD_LOGIC;
                    signal address : IN STD_LOGIC;
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal UART_TXD : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Serial_Port;

component Slider_Switches_avalon_parallel_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Slider_Switches_avalon_parallel_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC;
                    signal Slider_Switches_avalon_parallel_port_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal Slider_Switches_avalon_parallel_port_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Slider_Switches_avalon_parallel_port_slave_chipselect : OUT STD_LOGIC;
                    signal Slider_Switches_avalon_parallel_port_slave_read : OUT STD_LOGIC;
                    signal Slider_Switches_avalon_parallel_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Slider_Switches_avalon_parallel_port_slave_reset : OUT STD_LOGIC;
                    signal Slider_Switches_avalon_parallel_port_slave_write : OUT STD_LOGIC;
                    signal Slider_Switches_avalon_parallel_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Slider_Switches_avalon_parallel_port_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave : OUT STD_LOGIC
                 );
end component Slider_Switches_avalon_parallel_port_slave_arbitrator;

component Slider_Switches is 
           port (
                 -- inputs:
                    signal SW : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component Slider_Switches;

component VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_byteenable : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_chipselect : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_read : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_write : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave : OUT STD_LOGIC
                 );
end component VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator;

component VGA_Char_Buffer_avalon_char_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_address : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_control_slave_chipselect : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_read : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_control_slave_reset : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_write : OUT STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave : OUT STD_LOGIC
                 );
end component VGA_Char_Buffer_avalon_char_control_slave_arbitrator;

component VGA_Char_Buffer_avalon_char_source_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_foreground_sink_ready_from_sa : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal VGA_Char_Buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Char_Buffer_avalon_char_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Char_Buffer_avalon_char_source_ready : OUT STD_LOGIC
                 );
end component VGA_Char_Buffer_avalon_char_source_arbitrator;

component VGA_Char_Buffer is 
           port (
                 -- inputs:
                    signal buf_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal buf_byteenable : IN STD_LOGIC;
                    signal buf_chipselect : IN STD_LOGIC;
                    signal buf_read : IN STD_LOGIC;
                    signal buf_write : IN STD_LOGIC;
                    signal buf_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal ctrl_address : IN STD_LOGIC;
                    signal ctrl_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ctrl_chipselect : IN STD_LOGIC;
                    signal ctrl_read : IN STD_LOGIC;
                    signal ctrl_write : IN STD_LOGIC;
                    signal ctrl_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal stream_ready : IN STD_LOGIC;

                 -- outputs:
                    signal buf_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal buf_waitrequest : OUT STD_LOGIC;
                    signal ctrl_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal stream_endofpacket : OUT STD_LOGIC;
                    signal stream_startofpacket : OUT STD_LOGIC;
                    signal stream_valid : OUT STD_LOGIC
                 );
end component VGA_Char_Buffer;

component VGA_Controller_avalon_vga_sink_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Controller_avalon_vga_sink_ready : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Controller_avalon_vga_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Controller_avalon_vga_sink_endofpacket : OUT STD_LOGIC;
                    signal VGA_Controller_avalon_vga_sink_ready_from_sa : OUT STD_LOGIC;
                    signal VGA_Controller_avalon_vga_sink_reset : OUT STD_LOGIC;
                    signal VGA_Controller_avalon_vga_sink_startofpacket : OUT STD_LOGIC;
                    signal VGA_Controller_avalon_vga_sink_valid : OUT STD_LOGIC
                 );
end component VGA_Controller_avalon_vga_sink_arbitrator;

component VGA_Controller is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal endofpacket : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal startofpacket : IN STD_LOGIC;
                    signal valid : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_B : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_BLANK : OUT STD_LOGIC;
                    signal VGA_CLK : OUT STD_LOGIC;
                    signal VGA_G : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_HS : OUT STD_LOGIC;
                    signal VGA_R : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_SYNC : OUT STD_LOGIC;
                    signal VGA_VS : OUT STD_LOGIC;
                    signal ready : OUT STD_LOGIC
                 );
end component VGA_Controller;

component VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal Alpha_Blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                    signal Alpha_Blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                    signal Alpha_Blending_avalon_blended_source_valid : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket : OUT STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa : OUT STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket : OUT STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid : OUT STD_LOGIC
                 );
end component VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator;

component VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Controller_avalon_vga_sink_ready_from_sa : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready : OUT STD_LOGIC
                 );
end component VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator;

component VGA_Dual_Clock_FIFO is 
           port (
                 -- inputs:
                    signal clk_stream_in : IN STD_LOGIC;
                    signal clk_stream_out : IN STD_LOGIC;
                    signal stream_in_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_in_endofpacket : IN STD_LOGIC;
                    signal stream_in_startofpacket : IN STD_LOGIC;
                    signal stream_in_valid : IN STD_LOGIC;
                    signal stream_out_ready : IN STD_LOGIC;

                 -- outputs:
                    signal stream_in_ready : OUT STD_LOGIC;
                    signal stream_out_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_out_endofpacket : OUT STD_LOGIC;
                    signal stream_out_startofpacket : OUT STD_LOGIC;
                    signal stream_out_valid : OUT STD_LOGIC
                 );
end component VGA_Dual_Clock_FIFO;

component VGA_Pixel_Buffer_avalon_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal CPU_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_control_slave_read : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_control_slave_write : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave : OUT STD_LOGIC
                 );
end component VGA_Pixel_Buffer_avalon_control_slave_arbitrator;

component VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator is 
           port (
                 -- inputs:
                    signal SRAM_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal d1_SRAM_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_reset : OUT STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest : OUT STD_LOGIC
                 );
end component VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator;

component VGA_Pixel_Buffer_avalon_pixel_source_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Pixel_Buffer_avalon_pixel_source_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_source_valid : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_Buffer_avalon_pixel_source_ready : OUT STD_LOGIC
                 );
end component VGA_Pixel_Buffer_avalon_pixel_source_arbitrator;

component VGA_Pixel_Buffer is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_ready : IN STD_LOGIC;

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_arbiterlock : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal stream_endofpacket : OUT STD_LOGIC;
                    signal stream_startofpacket : OUT STD_LOGIC;
                    signal stream_valid : OUT STD_LOGIC
                 );
end component VGA_Pixel_Buffer;

component VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Pixel_Buffer_avalon_pixel_source_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_Buffer_avalon_pixel_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Buffer_avalon_pixel_source_valid : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket : OUT STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa : OUT STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset : OUT STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket : OUT STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid : OUT STD_LOGIC
                 );
end component VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator;

component VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready : OUT STD_LOGIC
                 );
end component VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator;

component VGA_Pixel_RGB_Resampler is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal stream_in_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal stream_in_endofpacket : IN STD_LOGIC;
                    signal stream_in_startofpacket : IN STD_LOGIC;
                    signal stream_in_valid : IN STD_LOGIC;
                    signal stream_out_ready : IN STD_LOGIC;

                 -- outputs:
                    signal stream_in_ready : OUT STD_LOGIC;
                    signal stream_out_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_out_endofpacket : OUT STD_LOGIC;
                    signal stream_out_startofpacket : OUT STD_LOGIC;
                    signal stream_out_valid : OUT STD_LOGIC
                 );
end component VGA_Pixel_RGB_Resampler;

component VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator is 
           port (
                 -- inputs:
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_ready : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket : OUT STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa : OUT STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_reset : OUT STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket : OUT STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_sink_valid : OUT STD_LOGIC
                 );
end component VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator;

component VGA_Pixel_Scaler_avalon_scaler_source_arbitrator is 
           port (
                 -- inputs:
                    signal Alpha_Blending_avalon_background_sink_ready_from_sa : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal VGA_Pixel_Scaler_avalon_scaler_source_endofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_startofpacket : IN STD_LOGIC;
                    signal VGA_Pixel_Scaler_avalon_scaler_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_Pixel_Scaler_avalon_scaler_source_ready : OUT STD_LOGIC
                 );
end component VGA_Pixel_Scaler_avalon_scaler_source_arbitrator;

component VGA_Pixel_Scaler is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal stream_in_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_in_endofpacket : IN STD_LOGIC;
                    signal stream_in_startofpacket : IN STD_LOGIC;
                    signal stream_in_valid : IN STD_LOGIC;
                    signal stream_out_ready : IN STD_LOGIC;

                 -- outputs:
                    signal stream_in_ready : OUT STD_LOGIC;
                    signal stream_out_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_out_endofpacket : OUT STD_LOGIC;
                    signal stream_out_startofpacket : OUT STD_LOGIC;
                    signal stream_out_valid : OUT STD_LOGIC
                 );
end component VGA_Pixel_Scaler;

component nios_system_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CPU_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal CPU_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal CPU_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_waitrequest : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal nios_system_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal nios_system_clock_0_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios_system_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal CPU_data_master_byteenable_nios_system_clock_0_in : OUT STD_LOGIC;
                    signal CPU_data_master_granted_nios_system_clock_0_in : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_nios_system_clock_0_in : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_nios_system_clock_0_in : OUT STD_LOGIC;
                    signal CPU_data_master_requests_nios_system_clock_0_in : OUT STD_LOGIC;
                    signal d1_nios_system_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_address : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_nativeaddress : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_read : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios_system_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_write : OUT STD_LOGIC;
                    signal nios_system_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios_system_clock_0_in_arbitrator;

component nios_system_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal External_Clocks_avalon_clocks_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_External_Clocks_avalon_clocks_slave_end_xfer : IN STD_LOGIC;
                    signal nios_system_clock_0_out_address : IN STD_LOGIC;
                    signal nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                    signal nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                    signal nios_system_clock_0_out_read : IN STD_LOGIC;
                    signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                    signal nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave : IN STD_LOGIC;
                    signal nios_system_clock_0_out_write : IN STD_LOGIC;
                    signal nios_system_clock_0_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios_system_clock_0_out_address_to_slave : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios_system_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal nios_system_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component nios_system_clock_0_out_arbitrator;

component nios_system_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC;
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC;
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC;
                    signal master_nativeaddress : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios_system_clock_0;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal CPU_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal CPU_data_master_read : IN STD_LOGIC;
                    signal CPU_data_master_write : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal CPU_data_master_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal CPU_data_master_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component nios_system_reset_sys_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios_system_reset_sys_clk_domain_synch_module;

component nios_system_reset_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios_system_reset_clk_domain_synch_module;

component nios_system_reset_vga_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios_system_reset_vga_clk_domain_synch_module;

                signal AV_Config_avalon_av_config_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_read :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal AV_Config_avalon_av_config_slave_reset :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_waitrequest :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_waitrequest_from_sa :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_write :  STD_LOGIC;
                signal AV_Config_avalon_av_config_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Alpha_Blending_avalon_background_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal Alpha_Blending_avalon_background_sink_endofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_background_sink_ready :  STD_LOGIC;
                signal Alpha_Blending_avalon_background_sink_ready_from_sa :  STD_LOGIC;
                signal Alpha_Blending_avalon_background_sink_startofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_background_sink_valid :  STD_LOGIC;
                signal Alpha_Blending_avalon_blended_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal Alpha_Blending_avalon_blended_source_endofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_blended_source_ready :  STD_LOGIC;
                signal Alpha_Blending_avalon_blended_source_startofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_blended_source_valid :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_data :  STD_LOGIC_VECTOR (39 DOWNTO 0);
                signal Alpha_Blending_avalon_foreground_sink_endofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_ready :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_ready_from_sa :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_reset :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_startofpacket :  STD_LOGIC;
                signal Alpha_Blending_avalon_foreground_sink_valid :  STD_LOGIC;
                signal Audio_avalon_audio_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Audio_avalon_audio_slave_chipselect :  STD_LOGIC;
                signal Audio_avalon_audio_slave_irq :  STD_LOGIC;
                signal Audio_avalon_audio_slave_irq_from_sa :  STD_LOGIC;
                signal Audio_avalon_audio_slave_read :  STD_LOGIC;
                signal Audio_avalon_audio_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Audio_avalon_audio_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Audio_avalon_audio_slave_reset :  STD_LOGIC;
                signal Audio_avalon_audio_slave_write :  STD_LOGIC;
                signal Audio_avalon_audio_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_clk_en :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_done :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_n :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_start :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_status :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal CPU_custom_instruction_master_reset_n :  STD_LOGIC;
                signal CPU_custom_instruction_master_start_CPU_fpoint_s1 :  STD_LOGIC;
                signal CPU_data_master_address :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal CPU_data_master_address_to_slave :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal CPU_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal CPU_data_master_byteenable_SDRAM_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_byteenable_SRAM_avalon_sram_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal CPU_data_master_byteenable_nios_system_clock_0_in :  STD_LOGIC;
                signal CPU_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal CPU_data_master_dbs_write_8 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal CPU_data_master_debugaccess :  STD_LOGIC;
                signal CPU_data_master_granted_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Audio_avalon_audio_slave :  STD_LOGIC;
                signal CPU_data_master_granted_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Interval_Timer_s1 :  STD_LOGIC;
                signal CPU_data_master_granted_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal CPU_data_master_granted_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_granted_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal CPU_data_master_granted_nios_system_clock_0_in :  STD_LOGIC;
                signal CPU_data_master_granted_sysid_control_slave :  STD_LOGIC;
                signal CPU_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Audio_avalon_audio_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Interval_Timer_s1 :  STD_LOGIC;
                signal CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_qualified_request_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal CPU_data_master_qualified_request_nios_system_clock_0_in :  STD_LOGIC;
                signal CPU_data_master_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal CPU_data_master_read :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Audio_avalon_audio_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Interval_Timer_s1 :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_SDRAM_s1_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_nios_system_clock_0_in :  STD_LOGIC;
                signal CPU_data_master_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal CPU_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_data_master_requests_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Audio_avalon_audio_slave :  STD_LOGIC;
                signal CPU_data_master_requests_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Interval_Timer_s1 :  STD_LOGIC;
                signal CPU_data_master_requests_JTAG_UART_avalon_jtag_slave :  STD_LOGIC;
                signal CPU_data_master_requests_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_SDRAM_s1 :  STD_LOGIC;
                signal CPU_data_master_requests_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal CPU_data_master_requests_nios_system_clock_0_in :  STD_LOGIC;
                signal CPU_data_master_requests_sysid_control_slave :  STD_LOGIC;
                signal CPU_data_master_waitrequest :  STD_LOGIC;
                signal CPU_data_master_write :  STD_LOGIC;
                signal CPU_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_fpoint_s1_clk_en :  STD_LOGIC;
                signal CPU_fpoint_s1_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_fpoint_s1_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_fpoint_s1_done :  STD_LOGIC;
                signal CPU_fpoint_s1_done_from_sa :  STD_LOGIC;
                signal CPU_fpoint_s1_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_fpoint_s1_reset :  STD_LOGIC;
                signal CPU_fpoint_s1_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_fpoint_s1_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_fpoint_s1_select :  STD_LOGIC;
                signal CPU_fpoint_s1_start :  STD_LOGIC;
                signal CPU_instruction_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal CPU_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal CPU_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal CPU_instruction_master_granted_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_instruction_master_granted_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_latency_counter :  STD_LOGIC;
                signal CPU_instruction_master_qualified_request_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_instruction_master_qualified_request_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_read :  STD_LOGIC;
                signal CPU_instruction_master_read_data_valid_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_instruction_master_read_data_valid_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register :  STD_LOGIC;
                signal CPU_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_instruction_master_readdatavalid :  STD_LOGIC;
                signal CPU_instruction_master_requests_CPU_jtag_debug_module :  STD_LOGIC;
                signal CPU_instruction_master_requests_SDRAM_s1 :  STD_LOGIC;
                signal CPU_instruction_master_waitrequest :  STD_LOGIC;
                signal CPU_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal CPU_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal CPU_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal CPU_jtag_debug_module_chipselect :  STD_LOGIC;
                signal CPU_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal CPU_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal CPU_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal CPU_jtag_debug_module_write :  STD_LOGIC;
                signal CPU_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_address :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_chipselect :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_read :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal Char_LCD_16x2_avalon_lcd_slave_reset :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_waitrequest :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_write :  STD_LOGIC;
                signal Char_LCD_16x2_avalon_lcd_slave_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_irq :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_irq_from_sa :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Expansion_JP1_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Expansion_JP1_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_irq :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_irq_from_sa :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Expansion_JP2_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Expansion_JP2_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal External_Clocks_avalon_clocks_slave_address :  STD_LOGIC;
                signal External_Clocks_avalon_clocks_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal External_Clocks_avalon_clocks_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Green_LEDs_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Green_LEDs_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX3_HEX0_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal HEX3_HEX0_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX7_HEX4_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal HEX7_HEX4_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Interval_Timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Interval_Timer_s1_chipselect :  STD_LOGIC;
                signal Interval_Timer_s1_irq :  STD_LOGIC;
                signal Interval_Timer_s1_irq_from_sa :  STD_LOGIC;
                signal Interval_Timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal Interval_Timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal Interval_Timer_s1_reset_n :  STD_LOGIC;
                signal Interval_Timer_s1_write_n :  STD_LOGIC;
                signal Interval_Timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_address :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_irq :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal JTAG_UART_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_address :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_chipselect :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_irq :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_irq_from_sa :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_read :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal PS2_Port_avalon_ps2_slave_reset :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_waitrequest :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_waitrequest_from_sa :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_write :  STD_LOGIC;
                signal PS2_Port_avalon_ps2_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_irq :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_irq_from_sa :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Pushbuttons_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Pushbuttons_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Red_LEDs_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Red_LEDs_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal SDRAM_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal SDRAM_s1_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SDRAM_s1_chipselect :  STD_LOGIC;
                signal SDRAM_s1_read_n :  STD_LOGIC;
                signal SDRAM_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SDRAM_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SDRAM_s1_readdatavalid :  STD_LOGIC;
                signal SDRAM_s1_reset_n :  STD_LOGIC;
                signal SDRAM_s1_waitrequest :  STD_LOGIC;
                signal SDRAM_s1_waitrequest_from_sa :  STD_LOGIC;
                signal SDRAM_s1_write_n :  STD_LOGIC;
                signal SDRAM_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SRAM_avalon_sram_slave_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal SRAM_avalon_sram_slave_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal SRAM_avalon_sram_slave_read :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SRAM_avalon_sram_slave_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SRAM_avalon_sram_slave_readdatavalid :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_reset :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_write :  STD_LOGIC;
                signal SRAM_avalon_sram_slave_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_address :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_chipselect :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_irq :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_irq_from_sa :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_read :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Serial_Port_avalon_rs232_slave_reset :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_write :  STD_LOGIC;
                signal Serial_Port_avalon_rs232_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_chipselect :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_read :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Slider_Switches_avalon_parallel_port_slave_reset :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_write :  STD_LOGIC;
                signal Slider_Switches_avalon_parallel_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_byteenable :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_chipselect :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_read :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_write :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_buffer_slave_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_address :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_chipselect :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_read :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_control_slave_reset :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_write :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_control_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_source_data :  STD_LOGIC_VECTOR (39 DOWNTO 0);
                signal VGA_Char_Buffer_avalon_char_source_endofpacket :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_source_ready :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_source_startofpacket :  STD_LOGIC;
                signal VGA_Char_Buffer_avalon_char_source_valid :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Controller_avalon_vga_sink_endofpacket :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_ready :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_ready_from_sa :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_reset :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_startofpacket :  STD_LOGIC;
                signal VGA_Controller_avalon_vga_sink_valid :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket :  STD_LOGIC;
                signal VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_read :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_control_slave_write :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_control_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_reset :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_source_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal VGA_Pixel_Buffer_avalon_pixel_source_endofpacket :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_source_ready :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_source_startofpacket :  STD_LOGIC;
                signal VGA_Pixel_Buffer_avalon_pixel_source_valid :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket :  STD_LOGIC;
                signal VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_ready :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_reset :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_sink_valid :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal VGA_Pixel_Scaler_avalon_scaler_source_endofpacket :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_source_ready :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_source_startofpacket :  STD_LOGIC;
                signal VGA_Pixel_Scaler_avalon_scaler_source_valid :  STD_LOGIC;
                signal clk_reset_n :  STD_LOGIC;
                signal d1_AV_Config_avalon_av_config_slave_end_xfer :  STD_LOGIC;
                signal d1_Audio_avalon_audio_slave_end_xfer :  STD_LOGIC;
                signal d1_CPU_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer :  STD_LOGIC;
                signal d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_External_Clocks_avalon_clocks_slave_end_xfer :  STD_LOGIC;
                signal d1_Green_LEDs_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_Interval_Timer_s1_end_xfer :  STD_LOGIC;
                signal d1_JTAG_UART_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_PS2_Port_avalon_ps2_slave_end_xfer :  STD_LOGIC;
                signal d1_Pushbuttons_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_Red_LEDs_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_SDRAM_s1_end_xfer :  STD_LOGIC;
                signal d1_SRAM_avalon_sram_slave_end_xfer :  STD_LOGIC;
                signal d1_Serial_Port_avalon_rs232_slave_end_xfer :  STD_LOGIC;
                signal d1_Slider_Switches_avalon_parallel_port_slave_end_xfer :  STD_LOGIC;
                signal d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer :  STD_LOGIC;
                signal d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer :  STD_LOGIC;
                signal d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer :  STD_LOGIC;
                signal d1_nios_system_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal internal_AUD_DACDAT_from_the_Audio :  STD_LOGIC;
                signal internal_HEX0_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX1_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX2_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX3_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX4_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX5_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX6_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_HEX7_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_I2C_SCLK_from_the_AV_Config :  STD_LOGIC;
                signal internal_LCD_BLON_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal internal_LCD_EN_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal internal_LCD_ON_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal internal_LCD_RS_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal internal_LCD_RW_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal internal_LEDG_from_the_Green_LEDs :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal internal_LEDR_from_the_Red_LEDs :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal internal_SRAM_ADDR_from_the_SRAM :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal internal_SRAM_CE_N_from_the_SRAM :  STD_LOGIC;
                signal internal_SRAM_LB_N_from_the_SRAM :  STD_LOGIC;
                signal internal_SRAM_OE_N_from_the_SRAM :  STD_LOGIC;
                signal internal_SRAM_UB_N_from_the_SRAM :  STD_LOGIC;
                signal internal_SRAM_WE_N_from_the_SRAM :  STD_LOGIC;
                signal internal_UART_TXD_from_the_Serial_Port :  STD_LOGIC;
                signal internal_VGA_BLANK_from_the_VGA_Controller :  STD_LOGIC;
                signal internal_VGA_B_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_CLK_from_the_VGA_Controller :  STD_LOGIC;
                signal internal_VGA_G_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_HS_from_the_VGA_Controller :  STD_LOGIC;
                signal internal_VGA_R_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_SYNC_from_the_VGA_Controller :  STD_LOGIC;
                signal internal_VGA_VS_from_the_VGA_Controller :  STD_LOGIC;
                signal internal_sys_clk :  STD_LOGIC;
                signal internal_vga_clk :  STD_LOGIC;
                signal internal_zs_addr_from_the_SDRAM :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal internal_zs_ba_from_the_SDRAM :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_SDRAM :  STD_LOGIC;
                signal internal_zs_cke_from_the_SDRAM :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_SDRAM :  STD_LOGIC;
                signal internal_zs_dqm_from_the_SDRAM :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_ras_n_from_the_SDRAM :  STD_LOGIC;
                signal internal_zs_we_n_from_the_SDRAM :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal nios_system_clock_0_in_address :  STD_LOGIC;
                signal nios_system_clock_0_in_endofpacket :  STD_LOGIC;
                signal nios_system_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios_system_clock_0_in_nativeaddress :  STD_LOGIC;
                signal nios_system_clock_0_in_read :  STD_LOGIC;
                signal nios_system_clock_0_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios_system_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios_system_clock_0_in_reset_n :  STD_LOGIC;
                signal nios_system_clock_0_in_waitrequest :  STD_LOGIC;
                signal nios_system_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios_system_clock_0_in_write :  STD_LOGIC;
                signal nios_system_clock_0_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios_system_clock_0_out_address :  STD_LOGIC;
                signal nios_system_clock_0_out_address_to_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_endofpacket :  STD_LOGIC;
                signal nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_nativeaddress :  STD_LOGIC;
                signal nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_read :  STD_LOGIC;
                signal nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave :  STD_LOGIC;
                signal nios_system_clock_0_out_reset_n :  STD_LOGIC;
                signal nios_system_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios_system_clock_0_out_write :  STD_LOGIC;
                signal nios_system_clock_0_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_clk_External_Clocks_AUD_CLK :  STD_LOGIC;
                signal out_clk_External_Clocks_SDRAM_CLK :  STD_LOGIC;
                signal out_clk_External_Clocks_VGA_CLK :  STD_LOGIC;
                signal out_clk_External_Clocks_sys_clk :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave :  STD_LOGIC;
                signal registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal sys_clk_reset_n :  STD_LOGIC;
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_clk_reset_n :  STD_LOGIC;

begin

  --the_AV_Config_avalon_av_config_slave, which is an e_instance
  the_AV_Config_avalon_av_config_slave : AV_Config_avalon_av_config_slave_arbitrator
    port map(
      AV_Config_avalon_av_config_slave_address => AV_Config_avalon_av_config_slave_address,
      AV_Config_avalon_av_config_slave_byteenable => AV_Config_avalon_av_config_slave_byteenable,
      AV_Config_avalon_av_config_slave_read => AV_Config_avalon_av_config_slave_read,
      AV_Config_avalon_av_config_slave_readdata_from_sa => AV_Config_avalon_av_config_slave_readdata_from_sa,
      AV_Config_avalon_av_config_slave_reset => AV_Config_avalon_av_config_slave_reset,
      AV_Config_avalon_av_config_slave_waitrequest_from_sa => AV_Config_avalon_av_config_slave_waitrequest_from_sa,
      AV_Config_avalon_av_config_slave_write => AV_Config_avalon_av_config_slave_write,
      AV_Config_avalon_av_config_slave_writedata => AV_Config_avalon_av_config_slave_writedata,
      CPU_data_master_granted_AV_Config_avalon_av_config_slave => CPU_data_master_granted_AV_Config_avalon_av_config_slave,
      CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave => CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave,
      CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave => CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave,
      CPU_data_master_requests_AV_Config_avalon_av_config_slave => CPU_data_master_requests_AV_Config_avalon_av_config_slave,
      d1_AV_Config_avalon_av_config_slave_end_xfer => d1_AV_Config_avalon_av_config_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave => registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave,
      AV_Config_avalon_av_config_slave_readdata => AV_Config_avalon_av_config_slave_readdata,
      AV_Config_avalon_av_config_slave_waitrequest => AV_Config_avalon_av_config_slave_waitrequest,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_AV_Config, which is an e_ptf_instance
  the_AV_Config : AV_Config
    port map(
      I2C_SCLK => internal_I2C_SCLK_from_the_AV_Config,
      I2C_SDAT => I2C_SDAT_to_and_from_the_AV_Config,
      readdata => AV_Config_avalon_av_config_slave_readdata,
      waitrequest => AV_Config_avalon_av_config_slave_waitrequest,
      address => AV_Config_avalon_av_config_slave_address,
      byteenable => AV_Config_avalon_av_config_slave_byteenable,
      clk => internal_sys_clk,
      read => AV_Config_avalon_av_config_slave_read,
      reset => AV_Config_avalon_av_config_slave_reset,
      write => AV_Config_avalon_av_config_slave_write,
      writedata => AV_Config_avalon_av_config_slave_writedata
    );


  --the_Alpha_Blending_avalon_background_sink, which is an e_instance
  the_Alpha_Blending_avalon_background_sink : Alpha_Blending_avalon_background_sink_arbitrator
    port map(
      Alpha_Blending_avalon_background_sink_data => Alpha_Blending_avalon_background_sink_data,
      Alpha_Blending_avalon_background_sink_endofpacket => Alpha_Blending_avalon_background_sink_endofpacket,
      Alpha_Blending_avalon_background_sink_ready_from_sa => Alpha_Blending_avalon_background_sink_ready_from_sa,
      Alpha_Blending_avalon_background_sink_startofpacket => Alpha_Blending_avalon_background_sink_startofpacket,
      Alpha_Blending_avalon_background_sink_valid => Alpha_Blending_avalon_background_sink_valid,
      Alpha_Blending_avalon_background_sink_ready => Alpha_Blending_avalon_background_sink_ready,
      VGA_Pixel_Scaler_avalon_scaler_source_data => VGA_Pixel_Scaler_avalon_scaler_source_data,
      VGA_Pixel_Scaler_avalon_scaler_source_endofpacket => VGA_Pixel_Scaler_avalon_scaler_source_endofpacket,
      VGA_Pixel_Scaler_avalon_scaler_source_startofpacket => VGA_Pixel_Scaler_avalon_scaler_source_startofpacket,
      VGA_Pixel_Scaler_avalon_scaler_source_valid => VGA_Pixel_Scaler_avalon_scaler_source_valid,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Alpha_Blending_avalon_foreground_sink, which is an e_instance
  the_Alpha_Blending_avalon_foreground_sink : Alpha_Blending_avalon_foreground_sink_arbitrator
    port map(
      Alpha_Blending_avalon_foreground_sink_data => Alpha_Blending_avalon_foreground_sink_data,
      Alpha_Blending_avalon_foreground_sink_endofpacket => Alpha_Blending_avalon_foreground_sink_endofpacket,
      Alpha_Blending_avalon_foreground_sink_ready_from_sa => Alpha_Blending_avalon_foreground_sink_ready_from_sa,
      Alpha_Blending_avalon_foreground_sink_reset => Alpha_Blending_avalon_foreground_sink_reset,
      Alpha_Blending_avalon_foreground_sink_startofpacket => Alpha_Blending_avalon_foreground_sink_startofpacket,
      Alpha_Blending_avalon_foreground_sink_valid => Alpha_Blending_avalon_foreground_sink_valid,
      Alpha_Blending_avalon_foreground_sink_ready => Alpha_Blending_avalon_foreground_sink_ready,
      VGA_Char_Buffer_avalon_char_source_data => VGA_Char_Buffer_avalon_char_source_data,
      VGA_Char_Buffer_avalon_char_source_endofpacket => VGA_Char_Buffer_avalon_char_source_endofpacket,
      VGA_Char_Buffer_avalon_char_source_startofpacket => VGA_Char_Buffer_avalon_char_source_startofpacket,
      VGA_Char_Buffer_avalon_char_source_valid => VGA_Char_Buffer_avalon_char_source_valid,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Alpha_Blending_avalon_blended_source, which is an e_instance
  the_Alpha_Blending_avalon_blended_source : Alpha_Blending_avalon_blended_source_arbitrator
    port map(
      Alpha_Blending_avalon_blended_source_ready => Alpha_Blending_avalon_blended_source_ready,
      Alpha_Blending_avalon_blended_source_data => Alpha_Blending_avalon_blended_source_data,
      Alpha_Blending_avalon_blended_source_endofpacket => Alpha_Blending_avalon_blended_source_endofpacket,
      Alpha_Blending_avalon_blended_source_startofpacket => Alpha_Blending_avalon_blended_source_startofpacket,
      Alpha_Blending_avalon_blended_source_valid => Alpha_Blending_avalon_blended_source_valid,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Alpha_Blending, which is an e_ptf_instance
  the_Alpha_Blending : Alpha_Blending
    port map(
      background_ready => Alpha_Blending_avalon_background_sink_ready,
      foreground_ready => Alpha_Blending_avalon_foreground_sink_ready,
      output_data => Alpha_Blending_avalon_blended_source_data,
      output_endofpacket => Alpha_Blending_avalon_blended_source_endofpacket,
      output_startofpacket => Alpha_Blending_avalon_blended_source_startofpacket,
      output_valid => Alpha_Blending_avalon_blended_source_valid,
      background_data => Alpha_Blending_avalon_background_sink_data,
      background_endofpacket => Alpha_Blending_avalon_background_sink_endofpacket,
      background_startofpacket => Alpha_Blending_avalon_background_sink_startofpacket,
      background_valid => Alpha_Blending_avalon_background_sink_valid,
      clk => internal_sys_clk,
      foreground_data => Alpha_Blending_avalon_foreground_sink_data,
      foreground_endofpacket => Alpha_Blending_avalon_foreground_sink_endofpacket,
      foreground_startofpacket => Alpha_Blending_avalon_foreground_sink_startofpacket,
      foreground_valid => Alpha_Blending_avalon_foreground_sink_valid,
      output_ready => Alpha_Blending_avalon_blended_source_ready,
      reset => Alpha_Blending_avalon_foreground_sink_reset
    );


  --the_Audio_avalon_audio_slave, which is an e_instance
  the_Audio_avalon_audio_slave : Audio_avalon_audio_slave_arbitrator
    port map(
      Audio_avalon_audio_slave_address => Audio_avalon_audio_slave_address,
      Audio_avalon_audio_slave_chipselect => Audio_avalon_audio_slave_chipselect,
      Audio_avalon_audio_slave_irq_from_sa => Audio_avalon_audio_slave_irq_from_sa,
      Audio_avalon_audio_slave_read => Audio_avalon_audio_slave_read,
      Audio_avalon_audio_slave_readdata_from_sa => Audio_avalon_audio_slave_readdata_from_sa,
      Audio_avalon_audio_slave_reset => Audio_avalon_audio_slave_reset,
      Audio_avalon_audio_slave_write => Audio_avalon_audio_slave_write,
      Audio_avalon_audio_slave_writedata => Audio_avalon_audio_slave_writedata,
      CPU_data_master_granted_Audio_avalon_audio_slave => CPU_data_master_granted_Audio_avalon_audio_slave,
      CPU_data_master_qualified_request_Audio_avalon_audio_slave => CPU_data_master_qualified_request_Audio_avalon_audio_slave,
      CPU_data_master_read_data_valid_Audio_avalon_audio_slave => CPU_data_master_read_data_valid_Audio_avalon_audio_slave,
      CPU_data_master_requests_Audio_avalon_audio_slave => CPU_data_master_requests_Audio_avalon_audio_slave,
      d1_Audio_avalon_audio_slave_end_xfer => d1_Audio_avalon_audio_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave => registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave,
      Audio_avalon_audio_slave_irq => Audio_avalon_audio_slave_irq,
      Audio_avalon_audio_slave_readdata => Audio_avalon_audio_slave_readdata,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Audio, which is an e_ptf_instance
  the_Audio : Audio
    port map(
      AUD_ADCLRCK => AUD_ADCLRCK_to_and_from_the_Audio,
      AUD_BCLK => AUD_BCLK_to_and_from_the_Audio,
      AUD_DACDAT => internal_AUD_DACDAT_from_the_Audio,
      AUD_DACLRCK => AUD_DACLRCK_to_and_from_the_Audio,
      irq => Audio_avalon_audio_slave_irq,
      readdata => Audio_avalon_audio_slave_readdata,
      AUD_ADCDAT => AUD_ADCDAT_to_the_Audio,
      address => Audio_avalon_audio_slave_address,
      chipselect => Audio_avalon_audio_slave_chipselect,
      clk => internal_sys_clk,
      read => Audio_avalon_audio_slave_read,
      reset => Audio_avalon_audio_slave_reset,
      write => Audio_avalon_audio_slave_write,
      writedata => Audio_avalon_audio_slave_writedata
    );


  --the_CPU_jtag_debug_module, which is an e_instance
  the_CPU_jtag_debug_module : CPU_jtag_debug_module_arbitrator
    port map(
      CPU_data_master_granted_CPU_jtag_debug_module => CPU_data_master_granted_CPU_jtag_debug_module,
      CPU_data_master_qualified_request_CPU_jtag_debug_module => CPU_data_master_qualified_request_CPU_jtag_debug_module,
      CPU_data_master_read_data_valid_CPU_jtag_debug_module => CPU_data_master_read_data_valid_CPU_jtag_debug_module,
      CPU_data_master_requests_CPU_jtag_debug_module => CPU_data_master_requests_CPU_jtag_debug_module,
      CPU_instruction_master_granted_CPU_jtag_debug_module => CPU_instruction_master_granted_CPU_jtag_debug_module,
      CPU_instruction_master_qualified_request_CPU_jtag_debug_module => CPU_instruction_master_qualified_request_CPU_jtag_debug_module,
      CPU_instruction_master_read_data_valid_CPU_jtag_debug_module => CPU_instruction_master_read_data_valid_CPU_jtag_debug_module,
      CPU_instruction_master_requests_CPU_jtag_debug_module => CPU_instruction_master_requests_CPU_jtag_debug_module,
      CPU_jtag_debug_module_address => CPU_jtag_debug_module_address,
      CPU_jtag_debug_module_begintransfer => CPU_jtag_debug_module_begintransfer,
      CPU_jtag_debug_module_byteenable => CPU_jtag_debug_module_byteenable,
      CPU_jtag_debug_module_chipselect => CPU_jtag_debug_module_chipselect,
      CPU_jtag_debug_module_debugaccess => CPU_jtag_debug_module_debugaccess,
      CPU_jtag_debug_module_readdata_from_sa => CPU_jtag_debug_module_readdata_from_sa,
      CPU_jtag_debug_module_resetrequest_from_sa => CPU_jtag_debug_module_resetrequest_from_sa,
      CPU_jtag_debug_module_write => CPU_jtag_debug_module_write,
      CPU_jtag_debug_module_writedata => CPU_jtag_debug_module_writedata,
      d1_CPU_jtag_debug_module_end_xfer => d1_CPU_jtag_debug_module_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_debugaccess => CPU_data_master_debugaccess,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      CPU_instruction_master_address_to_slave => CPU_instruction_master_address_to_slave,
      CPU_instruction_master_latency_counter => CPU_instruction_master_latency_counter,
      CPU_instruction_master_read => CPU_instruction_master_read,
      CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register => CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register,
      CPU_jtag_debug_module_readdata => CPU_jtag_debug_module_readdata,
      CPU_jtag_debug_module_resetrequest => CPU_jtag_debug_module_resetrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_CPU_custom_instruction_master, which is an e_instance
  the_CPU_custom_instruction_master : CPU_custom_instruction_master_arbitrator
    port map(
      CPU_custom_instruction_master_multi_done => CPU_custom_instruction_master_multi_done,
      CPU_custom_instruction_master_multi_result => CPU_custom_instruction_master_multi_result,
      CPU_custom_instruction_master_reset_n => CPU_custom_instruction_master_reset_n,
      CPU_custom_instruction_master_start_CPU_fpoint_s1 => CPU_custom_instruction_master_start_CPU_fpoint_s1,
      CPU_fpoint_s1_select => CPU_fpoint_s1_select,
      CPU_custom_instruction_master_multi_start => CPU_custom_instruction_master_multi_start,
      CPU_fpoint_s1_done_from_sa => CPU_fpoint_s1_done_from_sa,
      CPU_fpoint_s1_result_from_sa => CPU_fpoint_s1_result_from_sa,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_CPU_data_master, which is an e_instance
  the_CPU_data_master : CPU_data_master_arbitrator
    port map(
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_16 => CPU_data_master_dbs_write_16,
      CPU_data_master_dbs_write_8 => CPU_data_master_dbs_write_8,
      CPU_data_master_irq => CPU_data_master_irq,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_readdata => CPU_data_master_readdata,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      AV_Config_avalon_av_config_slave_readdata_from_sa => AV_Config_avalon_av_config_slave_readdata_from_sa,
      AV_Config_avalon_av_config_slave_waitrequest_from_sa => AV_Config_avalon_av_config_slave_waitrequest_from_sa,
      Audio_avalon_audio_slave_irq_from_sa => Audio_avalon_audio_slave_irq_from_sa,
      Audio_avalon_audio_slave_readdata_from_sa => Audio_avalon_audio_slave_readdata_from_sa,
      CPU_data_master_address => CPU_data_master_address,
      CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_byteenable_SDRAM_s1 => CPU_data_master_byteenable_SDRAM_s1,
      CPU_data_master_byteenable_SRAM_avalon_sram_slave => CPU_data_master_byteenable_SRAM_avalon_sram_slave,
      CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_byteenable_nios_system_clock_0_in => CPU_data_master_byteenable_nios_system_clock_0_in,
      CPU_data_master_granted_AV_Config_avalon_av_config_slave => CPU_data_master_granted_AV_Config_avalon_av_config_slave,
      CPU_data_master_granted_Audio_avalon_audio_slave => CPU_data_master_granted_Audio_avalon_audio_slave,
      CPU_data_master_granted_CPU_jtag_debug_module => CPU_data_master_granted_CPU_jtag_debug_module,
      CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_granted_Interval_Timer_s1 => CPU_data_master_granted_Interval_Timer_s1,
      CPU_data_master_granted_JTAG_UART_avalon_jtag_slave => CPU_data_master_granted_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_granted_PS2_Port_avalon_ps2_slave => CPU_data_master_granted_PS2_Port_avalon_ps2_slave,
      CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_granted_SDRAM_s1 => CPU_data_master_granted_SDRAM_s1,
      CPU_data_master_granted_SRAM_avalon_sram_slave => CPU_data_master_granted_SRAM_avalon_sram_slave,
      CPU_data_master_granted_Serial_Port_avalon_rs232_slave => CPU_data_master_granted_Serial_Port_avalon_rs232_slave,
      CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_granted_nios_system_clock_0_in => CPU_data_master_granted_nios_system_clock_0_in,
      CPU_data_master_granted_sysid_control_slave => CPU_data_master_granted_sysid_control_slave,
      CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave => CPU_data_master_qualified_request_AV_Config_avalon_av_config_slave,
      CPU_data_master_qualified_request_Audio_avalon_audio_slave => CPU_data_master_qualified_request_Audio_avalon_audio_slave,
      CPU_data_master_qualified_request_CPU_jtag_debug_module => CPU_data_master_qualified_request_CPU_jtag_debug_module,
      CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Interval_Timer_s1 => CPU_data_master_qualified_request_Interval_Timer_s1,
      CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave => CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave => CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave,
      CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_SDRAM_s1 => CPU_data_master_qualified_request_SDRAM_s1,
      CPU_data_master_qualified_request_SRAM_avalon_sram_slave => CPU_data_master_qualified_request_SRAM_avalon_sram_slave,
      CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave => CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave,
      CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_qualified_request_nios_system_clock_0_in => CPU_data_master_qualified_request_nios_system_clock_0_in,
      CPU_data_master_qualified_request_sysid_control_slave => CPU_data_master_qualified_request_sysid_control_slave,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave => CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave,
      CPU_data_master_read_data_valid_Audio_avalon_audio_slave => CPU_data_master_read_data_valid_Audio_avalon_audio_slave,
      CPU_data_master_read_data_valid_CPU_jtag_debug_module => CPU_data_master_read_data_valid_CPU_jtag_debug_module,
      CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Interval_Timer_s1 => CPU_data_master_read_data_valid_Interval_Timer_s1,
      CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave => CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave => CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave,
      CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_SDRAM_s1 => CPU_data_master_read_data_valid_SDRAM_s1,
      CPU_data_master_read_data_valid_SDRAM_s1_shift_register => CPU_data_master_read_data_valid_SDRAM_s1_shift_register,
      CPU_data_master_read_data_valid_SRAM_avalon_sram_slave => CPU_data_master_read_data_valid_SRAM_avalon_sram_slave,
      CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register => CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register,
      CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave => CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave,
      CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_read_data_valid_nios_system_clock_0_in => CPU_data_master_read_data_valid_nios_system_clock_0_in,
      CPU_data_master_read_data_valid_sysid_control_slave => CPU_data_master_read_data_valid_sysid_control_slave,
      CPU_data_master_requests_AV_Config_avalon_av_config_slave => CPU_data_master_requests_AV_Config_avalon_av_config_slave,
      CPU_data_master_requests_Audio_avalon_audio_slave => CPU_data_master_requests_Audio_avalon_audio_slave,
      CPU_data_master_requests_CPU_jtag_debug_module => CPU_data_master_requests_CPU_jtag_debug_module,
      CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_requests_Interval_Timer_s1 => CPU_data_master_requests_Interval_Timer_s1,
      CPU_data_master_requests_JTAG_UART_avalon_jtag_slave => CPU_data_master_requests_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_requests_PS2_Port_avalon_ps2_slave => CPU_data_master_requests_PS2_Port_avalon_ps2_slave,
      CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_requests_SDRAM_s1 => CPU_data_master_requests_SDRAM_s1,
      CPU_data_master_requests_SRAM_avalon_sram_slave => CPU_data_master_requests_SRAM_avalon_sram_slave,
      CPU_data_master_requests_Serial_Port_avalon_rs232_slave => CPU_data_master_requests_Serial_Port_avalon_rs232_slave,
      CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_requests_nios_system_clock_0_in => CPU_data_master_requests_nios_system_clock_0_in,
      CPU_data_master_requests_sysid_control_slave => CPU_data_master_requests_sysid_control_slave,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      CPU_jtag_debug_module_readdata_from_sa => CPU_jtag_debug_module_readdata_from_sa,
      Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa => Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa,
      Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa => Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa,
      Expansion_JP1_avalon_parallel_port_slave_irq_from_sa => Expansion_JP1_avalon_parallel_port_slave_irq_from_sa,
      Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa => Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa,
      Expansion_JP2_avalon_parallel_port_slave_irq_from_sa => Expansion_JP2_avalon_parallel_port_slave_irq_from_sa,
      Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa => Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa,
      Green_LEDs_avalon_parallel_port_slave_readdata_from_sa => Green_LEDs_avalon_parallel_port_slave_readdata_from_sa,
      HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa => HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa,
      HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa => HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa,
      Interval_Timer_s1_irq_from_sa => Interval_Timer_s1_irq_from_sa,
      Interval_Timer_s1_readdata_from_sa => Interval_Timer_s1_readdata_from_sa,
      JTAG_UART_avalon_jtag_slave_irq_from_sa => JTAG_UART_avalon_jtag_slave_irq_from_sa,
      JTAG_UART_avalon_jtag_slave_readdata_from_sa => JTAG_UART_avalon_jtag_slave_readdata_from_sa,
      JTAG_UART_avalon_jtag_slave_waitrequest_from_sa => JTAG_UART_avalon_jtag_slave_waitrequest_from_sa,
      PS2_Port_avalon_ps2_slave_irq_from_sa => PS2_Port_avalon_ps2_slave_irq_from_sa,
      PS2_Port_avalon_ps2_slave_readdata_from_sa => PS2_Port_avalon_ps2_slave_readdata_from_sa,
      PS2_Port_avalon_ps2_slave_waitrequest_from_sa => PS2_Port_avalon_ps2_slave_waitrequest_from_sa,
      Pushbuttons_avalon_parallel_port_slave_irq_from_sa => Pushbuttons_avalon_parallel_port_slave_irq_from_sa,
      Pushbuttons_avalon_parallel_port_slave_readdata_from_sa => Pushbuttons_avalon_parallel_port_slave_readdata_from_sa,
      Red_LEDs_avalon_parallel_port_slave_readdata_from_sa => Red_LEDs_avalon_parallel_port_slave_readdata_from_sa,
      SDRAM_s1_readdata_from_sa => SDRAM_s1_readdata_from_sa,
      SDRAM_s1_waitrequest_from_sa => SDRAM_s1_waitrequest_from_sa,
      SRAM_avalon_sram_slave_readdata_from_sa => SRAM_avalon_sram_slave_readdata_from_sa,
      Serial_Port_avalon_rs232_slave_irq_from_sa => Serial_Port_avalon_rs232_slave_irq_from_sa,
      Serial_Port_avalon_rs232_slave_readdata_from_sa => Serial_Port_avalon_rs232_slave_readdata_from_sa,
      Slider_Switches_avalon_parallel_port_slave_readdata_from_sa => Slider_Switches_avalon_parallel_port_slave_readdata_from_sa,
      VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa => VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa,
      VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa => VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa,
      VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa => VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa,
      VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa => VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa,
      clk => internal_sys_clk,
      d1_AV_Config_avalon_av_config_slave_end_xfer => d1_AV_Config_avalon_av_config_slave_end_xfer,
      d1_Audio_avalon_audio_slave_end_xfer => d1_Audio_avalon_audio_slave_end_xfer,
      d1_CPU_jtag_debug_module_end_xfer => d1_CPU_jtag_debug_module_end_xfer,
      d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer => d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer,
      d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer => d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer,
      d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer => d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer,
      d1_Green_LEDs_avalon_parallel_port_slave_end_xfer => d1_Green_LEDs_avalon_parallel_port_slave_end_xfer,
      d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer => d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer,
      d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer => d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer,
      d1_Interval_Timer_s1_end_xfer => d1_Interval_Timer_s1_end_xfer,
      d1_JTAG_UART_avalon_jtag_slave_end_xfer => d1_JTAG_UART_avalon_jtag_slave_end_xfer,
      d1_PS2_Port_avalon_ps2_slave_end_xfer => d1_PS2_Port_avalon_ps2_slave_end_xfer,
      d1_Pushbuttons_avalon_parallel_port_slave_end_xfer => d1_Pushbuttons_avalon_parallel_port_slave_end_xfer,
      d1_Red_LEDs_avalon_parallel_port_slave_end_xfer => d1_Red_LEDs_avalon_parallel_port_slave_end_xfer,
      d1_SDRAM_s1_end_xfer => d1_SDRAM_s1_end_xfer,
      d1_SRAM_avalon_sram_slave_end_xfer => d1_SRAM_avalon_sram_slave_end_xfer,
      d1_Serial_Port_avalon_rs232_slave_end_xfer => d1_Serial_Port_avalon_rs232_slave_end_xfer,
      d1_Slider_Switches_avalon_parallel_port_slave_end_xfer => d1_Slider_Switches_avalon_parallel_port_slave_end_xfer,
      d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer => d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer,
      d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer => d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer,
      d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer => d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer,
      d1_nios_system_clock_0_in_end_xfer => d1_nios_system_clock_0_in_end_xfer,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      nios_system_clock_0_in_readdata_from_sa => nios_system_clock_0_in_readdata_from_sa,
      nios_system_clock_0_in_waitrequest_from_sa => nios_system_clock_0_in_waitrequest_from_sa,
      registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave => registered_CPU_data_master_read_data_valid_AV_Config_avalon_av_config_slave,
      registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave => registered_CPU_data_master_read_data_valid_Audio_avalon_audio_slave,
      registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave => registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave,
      registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave => registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave,
      registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave,
      registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave => registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave,
      registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave => registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave,
      registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave => registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave,
      reset_n => sys_clk_reset_n,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa
    );


  --the_CPU_instruction_master, which is an e_instance
  the_CPU_instruction_master : CPU_instruction_master_arbitrator
    port map(
      CPU_instruction_master_address_to_slave => CPU_instruction_master_address_to_slave,
      CPU_instruction_master_dbs_address => CPU_instruction_master_dbs_address,
      CPU_instruction_master_latency_counter => CPU_instruction_master_latency_counter,
      CPU_instruction_master_readdata => CPU_instruction_master_readdata,
      CPU_instruction_master_readdatavalid => CPU_instruction_master_readdatavalid,
      CPU_instruction_master_waitrequest => CPU_instruction_master_waitrequest,
      CPU_instruction_master_address => CPU_instruction_master_address,
      CPU_instruction_master_granted_CPU_jtag_debug_module => CPU_instruction_master_granted_CPU_jtag_debug_module,
      CPU_instruction_master_granted_SDRAM_s1 => CPU_instruction_master_granted_SDRAM_s1,
      CPU_instruction_master_qualified_request_CPU_jtag_debug_module => CPU_instruction_master_qualified_request_CPU_jtag_debug_module,
      CPU_instruction_master_qualified_request_SDRAM_s1 => CPU_instruction_master_qualified_request_SDRAM_s1,
      CPU_instruction_master_read => CPU_instruction_master_read,
      CPU_instruction_master_read_data_valid_CPU_jtag_debug_module => CPU_instruction_master_read_data_valid_CPU_jtag_debug_module,
      CPU_instruction_master_read_data_valid_SDRAM_s1 => CPU_instruction_master_read_data_valid_SDRAM_s1,
      CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register => CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register,
      CPU_instruction_master_requests_CPU_jtag_debug_module => CPU_instruction_master_requests_CPU_jtag_debug_module,
      CPU_instruction_master_requests_SDRAM_s1 => CPU_instruction_master_requests_SDRAM_s1,
      CPU_jtag_debug_module_readdata_from_sa => CPU_jtag_debug_module_readdata_from_sa,
      SDRAM_s1_readdata_from_sa => SDRAM_s1_readdata_from_sa,
      SDRAM_s1_waitrequest_from_sa => SDRAM_s1_waitrequest_from_sa,
      clk => internal_sys_clk,
      d1_CPU_jtag_debug_module_end_xfer => d1_CPU_jtag_debug_module_end_xfer,
      d1_SDRAM_s1_end_xfer => d1_SDRAM_s1_end_xfer,
      reset_n => sys_clk_reset_n
    );


  --the_CPU, which is an e_ptf_instance
  the_CPU : CPU
    port map(
      M_ci_multi_a => CPU_custom_instruction_master_multi_a,
      M_ci_multi_b => CPU_custom_instruction_master_multi_b,
      M_ci_multi_c => CPU_custom_instruction_master_multi_c,
      M_ci_multi_clk_en => CPU_custom_instruction_master_multi_clk_en,
      M_ci_multi_dataa => CPU_custom_instruction_master_multi_dataa,
      M_ci_multi_datab => CPU_custom_instruction_master_multi_datab,
      M_ci_multi_estatus => CPU_custom_instruction_master_multi_estatus,
      M_ci_multi_ipending => CPU_custom_instruction_master_multi_ipending,
      M_ci_multi_n => CPU_custom_instruction_master_multi_n,
      M_ci_multi_readra => CPU_custom_instruction_master_multi_readra,
      M_ci_multi_readrb => CPU_custom_instruction_master_multi_readrb,
      M_ci_multi_start => CPU_custom_instruction_master_multi_start,
      M_ci_multi_status => CPU_custom_instruction_master_multi_status,
      M_ci_multi_writerc => CPU_custom_instruction_master_multi_writerc,
      d_address => CPU_data_master_address,
      d_byteenable => CPU_data_master_byteenable,
      d_read => CPU_data_master_read,
      d_write => CPU_data_master_write,
      d_writedata => CPU_data_master_writedata,
      i_address => CPU_instruction_master_address,
      i_read => CPU_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => CPU_data_master_debugaccess,
      jtag_debug_module_readdata => CPU_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => CPU_jtag_debug_module_resetrequest,
      M_ci_multi_done => CPU_custom_instruction_master_multi_done,
      M_ci_multi_result => CPU_custom_instruction_master_multi_result,
      clk => internal_sys_clk,
      d_irq => CPU_data_master_irq,
      d_readdata => CPU_data_master_readdata,
      d_waitrequest => CPU_data_master_waitrequest,
      i_readdata => CPU_instruction_master_readdata,
      i_readdatavalid => CPU_instruction_master_readdatavalid,
      i_waitrequest => CPU_instruction_master_waitrequest,
      jtag_debug_module_address => CPU_jtag_debug_module_address,
      jtag_debug_module_begintransfer => CPU_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => CPU_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => CPU_jtag_debug_module_debugaccess,
      jtag_debug_module_select => CPU_jtag_debug_module_chipselect,
      jtag_debug_module_write => CPU_jtag_debug_module_write,
      jtag_debug_module_writedata => CPU_jtag_debug_module_writedata,
      reset_n => CPU_custom_instruction_master_reset_n
    );


  --the_CPU_fpoint_s1, which is an e_instance
  the_CPU_fpoint_s1 : CPU_fpoint_s1_arbitrator
    port map(
      CPU_fpoint_s1_clk_en => CPU_fpoint_s1_clk_en,
      CPU_fpoint_s1_dataa => CPU_fpoint_s1_dataa,
      CPU_fpoint_s1_datab => CPU_fpoint_s1_datab,
      CPU_fpoint_s1_done_from_sa => CPU_fpoint_s1_done_from_sa,
      CPU_fpoint_s1_n => CPU_fpoint_s1_n,
      CPU_fpoint_s1_reset => CPU_fpoint_s1_reset,
      CPU_fpoint_s1_result_from_sa => CPU_fpoint_s1_result_from_sa,
      CPU_fpoint_s1_start => CPU_fpoint_s1_start,
      CPU_custom_instruction_master_multi_clk_en => CPU_custom_instruction_master_multi_clk_en,
      CPU_custom_instruction_master_multi_dataa => CPU_custom_instruction_master_multi_dataa,
      CPU_custom_instruction_master_multi_datab => CPU_custom_instruction_master_multi_datab,
      CPU_custom_instruction_master_multi_n => CPU_custom_instruction_master_multi_n,
      CPU_custom_instruction_master_start_CPU_fpoint_s1 => CPU_custom_instruction_master_start_CPU_fpoint_s1,
      CPU_fpoint_s1_done => CPU_fpoint_s1_done,
      CPU_fpoint_s1_result => CPU_fpoint_s1_result,
      CPU_fpoint_s1_select => CPU_fpoint_s1_select,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_CPU_fpoint, which is an e_ptf_instance
  the_CPU_fpoint : CPU_fpoint
    port map(
      done => CPU_fpoint_s1_done,
      result => CPU_fpoint_s1_result,
      clk => internal_sys_clk,
      clk_en => CPU_fpoint_s1_clk_en,
      dataa => CPU_fpoint_s1_dataa,
      datab => CPU_fpoint_s1_datab,
      n => CPU_fpoint_s1_n,
      reset => CPU_fpoint_s1_reset,
      start => CPU_fpoint_s1_start
    );


  --the_Char_LCD_16x2_avalon_lcd_slave, which is an e_instance
  the_Char_LCD_16x2_avalon_lcd_slave : Char_LCD_16x2_avalon_lcd_slave_arbitrator
    port map(
      CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_byteenable_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_granted_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_qualified_request_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_read_data_valid_Char_LCD_16x2_avalon_lcd_slave,
      CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave => CPU_data_master_requests_Char_LCD_16x2_avalon_lcd_slave,
      Char_LCD_16x2_avalon_lcd_slave_address => Char_LCD_16x2_avalon_lcd_slave_address,
      Char_LCD_16x2_avalon_lcd_slave_chipselect => Char_LCD_16x2_avalon_lcd_slave_chipselect,
      Char_LCD_16x2_avalon_lcd_slave_read => Char_LCD_16x2_avalon_lcd_slave_read,
      Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa => Char_LCD_16x2_avalon_lcd_slave_readdata_from_sa,
      Char_LCD_16x2_avalon_lcd_slave_reset => Char_LCD_16x2_avalon_lcd_slave_reset,
      Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa => Char_LCD_16x2_avalon_lcd_slave_waitrequest_from_sa,
      Char_LCD_16x2_avalon_lcd_slave_write => Char_LCD_16x2_avalon_lcd_slave_write,
      Char_LCD_16x2_avalon_lcd_slave_writedata => Char_LCD_16x2_avalon_lcd_slave_writedata,
      d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer => d1_Char_LCD_16x2_avalon_lcd_slave_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_8 => CPU_data_master_dbs_write_8,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      Char_LCD_16x2_avalon_lcd_slave_readdata => Char_LCD_16x2_avalon_lcd_slave_readdata,
      Char_LCD_16x2_avalon_lcd_slave_waitrequest => Char_LCD_16x2_avalon_lcd_slave_waitrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Char_LCD_16x2, which is an e_ptf_instance
  the_Char_LCD_16x2 : Char_LCD_16x2
    port map(
      LCD_BLON => internal_LCD_BLON_from_the_Char_LCD_16x2,
      LCD_DATA => LCD_DATA_to_and_from_the_Char_LCD_16x2,
      LCD_EN => internal_LCD_EN_from_the_Char_LCD_16x2,
      LCD_ON => internal_LCD_ON_from_the_Char_LCD_16x2,
      LCD_RS => internal_LCD_RS_from_the_Char_LCD_16x2,
      LCD_RW => internal_LCD_RW_from_the_Char_LCD_16x2,
      readdata => Char_LCD_16x2_avalon_lcd_slave_readdata,
      waitrequest => Char_LCD_16x2_avalon_lcd_slave_waitrequest,
      address => Char_LCD_16x2_avalon_lcd_slave_address,
      chipselect => Char_LCD_16x2_avalon_lcd_slave_chipselect,
      clk => internal_sys_clk,
      read => Char_LCD_16x2_avalon_lcd_slave_read,
      reset => Char_LCD_16x2_avalon_lcd_slave_reset,
      write => Char_LCD_16x2_avalon_lcd_slave_write,
      writedata => Char_LCD_16x2_avalon_lcd_slave_writedata
    );


  --the_Expansion_JP1_avalon_parallel_port_slave, which is an e_instance
  the_Expansion_JP1_avalon_parallel_port_slave : Expansion_JP1_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_granted_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_qualified_request_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave => CPU_data_master_requests_Expansion_JP1_avalon_parallel_port_slave,
      Expansion_JP1_avalon_parallel_port_slave_address => Expansion_JP1_avalon_parallel_port_slave_address,
      Expansion_JP1_avalon_parallel_port_slave_byteenable => Expansion_JP1_avalon_parallel_port_slave_byteenable,
      Expansion_JP1_avalon_parallel_port_slave_chipselect => Expansion_JP1_avalon_parallel_port_slave_chipselect,
      Expansion_JP1_avalon_parallel_port_slave_irq_from_sa => Expansion_JP1_avalon_parallel_port_slave_irq_from_sa,
      Expansion_JP1_avalon_parallel_port_slave_read => Expansion_JP1_avalon_parallel_port_slave_read,
      Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa => Expansion_JP1_avalon_parallel_port_slave_readdata_from_sa,
      Expansion_JP1_avalon_parallel_port_slave_reset => Expansion_JP1_avalon_parallel_port_slave_reset,
      Expansion_JP1_avalon_parallel_port_slave_write => Expansion_JP1_avalon_parallel_port_slave_write,
      Expansion_JP1_avalon_parallel_port_slave_writedata => Expansion_JP1_avalon_parallel_port_slave_writedata,
      d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer => d1_Expansion_JP1_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Expansion_JP1_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Expansion_JP1_avalon_parallel_port_slave_irq => Expansion_JP1_avalon_parallel_port_slave_irq,
      Expansion_JP1_avalon_parallel_port_slave_readdata => Expansion_JP1_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Expansion_JP1, which is an e_ptf_instance
  the_Expansion_JP1 : Expansion_JP1
    port map(
      GPIO_0 => GPIO_0_to_and_from_the_Expansion_JP1,
      irq => Expansion_JP1_avalon_parallel_port_slave_irq,
      readdata => Expansion_JP1_avalon_parallel_port_slave_readdata,
      address => Expansion_JP1_avalon_parallel_port_slave_address,
      byteenable => Expansion_JP1_avalon_parallel_port_slave_byteenable,
      chipselect => Expansion_JP1_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Expansion_JP1_avalon_parallel_port_slave_read,
      reset => Expansion_JP1_avalon_parallel_port_slave_reset,
      write => Expansion_JP1_avalon_parallel_port_slave_write,
      writedata => Expansion_JP1_avalon_parallel_port_slave_writedata
    );


  --the_Expansion_JP2_avalon_parallel_port_slave, which is an e_instance
  the_Expansion_JP2_avalon_parallel_port_slave : Expansion_JP2_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_granted_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_qualified_request_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave => CPU_data_master_requests_Expansion_JP2_avalon_parallel_port_slave,
      Expansion_JP2_avalon_parallel_port_slave_address => Expansion_JP2_avalon_parallel_port_slave_address,
      Expansion_JP2_avalon_parallel_port_slave_byteenable => Expansion_JP2_avalon_parallel_port_slave_byteenable,
      Expansion_JP2_avalon_parallel_port_slave_chipselect => Expansion_JP2_avalon_parallel_port_slave_chipselect,
      Expansion_JP2_avalon_parallel_port_slave_irq_from_sa => Expansion_JP2_avalon_parallel_port_slave_irq_from_sa,
      Expansion_JP2_avalon_parallel_port_slave_read => Expansion_JP2_avalon_parallel_port_slave_read,
      Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa => Expansion_JP2_avalon_parallel_port_slave_readdata_from_sa,
      Expansion_JP2_avalon_parallel_port_slave_reset => Expansion_JP2_avalon_parallel_port_slave_reset,
      Expansion_JP2_avalon_parallel_port_slave_write => Expansion_JP2_avalon_parallel_port_slave_write,
      Expansion_JP2_avalon_parallel_port_slave_writedata => Expansion_JP2_avalon_parallel_port_slave_writedata,
      d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer => d1_Expansion_JP2_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Expansion_JP2_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Expansion_JP2_avalon_parallel_port_slave_irq => Expansion_JP2_avalon_parallel_port_slave_irq,
      Expansion_JP2_avalon_parallel_port_slave_readdata => Expansion_JP2_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Expansion_JP2, which is an e_ptf_instance
  the_Expansion_JP2 : Expansion_JP2
    port map(
      GPIO_1 => GPIO_1_to_and_from_the_Expansion_JP2,
      irq => Expansion_JP2_avalon_parallel_port_slave_irq,
      readdata => Expansion_JP2_avalon_parallel_port_slave_readdata,
      address => Expansion_JP2_avalon_parallel_port_slave_address,
      byteenable => Expansion_JP2_avalon_parallel_port_slave_byteenable,
      chipselect => Expansion_JP2_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Expansion_JP2_avalon_parallel_port_slave_read,
      reset => Expansion_JP2_avalon_parallel_port_slave_reset,
      write => Expansion_JP2_avalon_parallel_port_slave_write,
      writedata => Expansion_JP2_avalon_parallel_port_slave_writedata
    );


  --the_External_Clocks_avalon_clocks_slave, which is an e_instance
  the_External_Clocks_avalon_clocks_slave : External_Clocks_avalon_clocks_slave_arbitrator
    port map(
      External_Clocks_avalon_clocks_slave_address => External_Clocks_avalon_clocks_slave_address,
      External_Clocks_avalon_clocks_slave_readdata_from_sa => External_Clocks_avalon_clocks_slave_readdata_from_sa,
      d1_External_Clocks_avalon_clocks_slave_end_xfer => d1_External_Clocks_avalon_clocks_slave_end_xfer,
      nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave,
      External_Clocks_avalon_clocks_slave_readdata => External_Clocks_avalon_clocks_slave_readdata,
      clk => clk,
      nios_system_clock_0_out_address_to_slave => nios_system_clock_0_out_address_to_slave,
      nios_system_clock_0_out_read => nios_system_clock_0_out_read,
      nios_system_clock_0_out_write => nios_system_clock_0_out_write,
      reset_n => clk_reset_n
    );


  --audio_clk out_clk assignment, which is an e_assign
  audio_clk <= out_clk_External_Clocks_AUD_CLK;
  --sdram_clk out_clk assignment, which is an e_assign
  sdram_clk <= out_clk_External_Clocks_SDRAM_CLK;
  --vga_clk out_clk assignment, which is an e_assign
  internal_vga_clk <= out_clk_External_Clocks_VGA_CLK;
  --sys_clk out_clk assignment, which is an e_assign
  internal_sys_clk <= out_clk_External_Clocks_sys_clk;
  --the_External_Clocks, which is an e_ptf_instance
  the_External_Clocks : External_Clocks
    port map(
      AUD_CLK => out_clk_External_Clocks_AUD_CLK,
      SDRAM_CLK => out_clk_External_Clocks_SDRAM_CLK,
      VGA_CLK => out_clk_External_Clocks_VGA_CLK,
      readdata => External_Clocks_avalon_clocks_slave_readdata,
      sys_clk => out_clk_External_Clocks_sys_clk,
      CLOCK_27 => clk_27,
      CLOCK_50 => clk,
      address => External_Clocks_avalon_clocks_slave_address
    );


  --the_Green_LEDs_avalon_parallel_port_slave, which is an e_instance
  the_Green_LEDs_avalon_parallel_port_slave : Green_LEDs_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_granted_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_qualified_request_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave => CPU_data_master_requests_Green_LEDs_avalon_parallel_port_slave,
      Green_LEDs_avalon_parallel_port_slave_address => Green_LEDs_avalon_parallel_port_slave_address,
      Green_LEDs_avalon_parallel_port_slave_byteenable => Green_LEDs_avalon_parallel_port_slave_byteenable,
      Green_LEDs_avalon_parallel_port_slave_chipselect => Green_LEDs_avalon_parallel_port_slave_chipselect,
      Green_LEDs_avalon_parallel_port_slave_read => Green_LEDs_avalon_parallel_port_slave_read,
      Green_LEDs_avalon_parallel_port_slave_readdata_from_sa => Green_LEDs_avalon_parallel_port_slave_readdata_from_sa,
      Green_LEDs_avalon_parallel_port_slave_reset => Green_LEDs_avalon_parallel_port_slave_reset,
      Green_LEDs_avalon_parallel_port_slave_write => Green_LEDs_avalon_parallel_port_slave_write,
      Green_LEDs_avalon_parallel_port_slave_writedata => Green_LEDs_avalon_parallel_port_slave_writedata,
      d1_Green_LEDs_avalon_parallel_port_slave_end_xfer => d1_Green_LEDs_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Green_LEDs_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Green_LEDs_avalon_parallel_port_slave_readdata => Green_LEDs_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Green_LEDs, which is an e_ptf_instance
  the_Green_LEDs : Green_LEDs
    port map(
      LEDG => internal_LEDG_from_the_Green_LEDs,
      readdata => Green_LEDs_avalon_parallel_port_slave_readdata,
      address => Green_LEDs_avalon_parallel_port_slave_address,
      byteenable => Green_LEDs_avalon_parallel_port_slave_byteenable,
      chipselect => Green_LEDs_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Green_LEDs_avalon_parallel_port_slave_read,
      reset => Green_LEDs_avalon_parallel_port_slave_reset,
      write => Green_LEDs_avalon_parallel_port_slave_write,
      writedata => Green_LEDs_avalon_parallel_port_slave_writedata
    );


  --the_HEX3_HEX0_avalon_parallel_port_slave, which is an e_instance
  the_HEX3_HEX0_avalon_parallel_port_slave : HEX3_HEX0_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_granted_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_qualified_request_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave => CPU_data_master_requests_HEX3_HEX0_avalon_parallel_port_slave,
      HEX3_HEX0_avalon_parallel_port_slave_address => HEX3_HEX0_avalon_parallel_port_slave_address,
      HEX3_HEX0_avalon_parallel_port_slave_byteenable => HEX3_HEX0_avalon_parallel_port_slave_byteenable,
      HEX3_HEX0_avalon_parallel_port_slave_chipselect => HEX3_HEX0_avalon_parallel_port_slave_chipselect,
      HEX3_HEX0_avalon_parallel_port_slave_read => HEX3_HEX0_avalon_parallel_port_slave_read,
      HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa => HEX3_HEX0_avalon_parallel_port_slave_readdata_from_sa,
      HEX3_HEX0_avalon_parallel_port_slave_reset => HEX3_HEX0_avalon_parallel_port_slave_reset,
      HEX3_HEX0_avalon_parallel_port_slave_write => HEX3_HEX0_avalon_parallel_port_slave_write,
      HEX3_HEX0_avalon_parallel_port_slave_writedata => HEX3_HEX0_avalon_parallel_port_slave_writedata,
      d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer => d1_HEX3_HEX0_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_HEX3_HEX0_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      HEX3_HEX0_avalon_parallel_port_slave_readdata => HEX3_HEX0_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_HEX3_HEX0, which is an e_ptf_instance
  the_HEX3_HEX0 : HEX3_HEX0
    port map(
      HEX0 => internal_HEX0_from_the_HEX3_HEX0,
      HEX1 => internal_HEX1_from_the_HEX3_HEX0,
      HEX2 => internal_HEX2_from_the_HEX3_HEX0,
      HEX3 => internal_HEX3_from_the_HEX3_HEX0,
      readdata => HEX3_HEX0_avalon_parallel_port_slave_readdata,
      address => HEX3_HEX0_avalon_parallel_port_slave_address,
      byteenable => HEX3_HEX0_avalon_parallel_port_slave_byteenable,
      chipselect => HEX3_HEX0_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => HEX3_HEX0_avalon_parallel_port_slave_read,
      reset => HEX3_HEX0_avalon_parallel_port_slave_reset,
      write => HEX3_HEX0_avalon_parallel_port_slave_write,
      writedata => HEX3_HEX0_avalon_parallel_port_slave_writedata
    );


  --the_HEX7_HEX4_avalon_parallel_port_slave, which is an e_instance
  the_HEX7_HEX4_avalon_parallel_port_slave : HEX7_HEX4_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_granted_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_qualified_request_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave => CPU_data_master_requests_HEX7_HEX4_avalon_parallel_port_slave,
      HEX7_HEX4_avalon_parallel_port_slave_address => HEX7_HEX4_avalon_parallel_port_slave_address,
      HEX7_HEX4_avalon_parallel_port_slave_byteenable => HEX7_HEX4_avalon_parallel_port_slave_byteenable,
      HEX7_HEX4_avalon_parallel_port_slave_chipselect => HEX7_HEX4_avalon_parallel_port_slave_chipselect,
      HEX7_HEX4_avalon_parallel_port_slave_read => HEX7_HEX4_avalon_parallel_port_slave_read,
      HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa => HEX7_HEX4_avalon_parallel_port_slave_readdata_from_sa,
      HEX7_HEX4_avalon_parallel_port_slave_reset => HEX7_HEX4_avalon_parallel_port_slave_reset,
      HEX7_HEX4_avalon_parallel_port_slave_write => HEX7_HEX4_avalon_parallel_port_slave_write,
      HEX7_HEX4_avalon_parallel_port_slave_writedata => HEX7_HEX4_avalon_parallel_port_slave_writedata,
      d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer => d1_HEX7_HEX4_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_HEX7_HEX4_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      HEX7_HEX4_avalon_parallel_port_slave_readdata => HEX7_HEX4_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_HEX7_HEX4, which is an e_ptf_instance
  the_HEX7_HEX4 : HEX7_HEX4
    port map(
      HEX4 => internal_HEX4_from_the_HEX7_HEX4,
      HEX5 => internal_HEX5_from_the_HEX7_HEX4,
      HEX6 => internal_HEX6_from_the_HEX7_HEX4,
      HEX7 => internal_HEX7_from_the_HEX7_HEX4,
      readdata => HEX7_HEX4_avalon_parallel_port_slave_readdata,
      address => HEX7_HEX4_avalon_parallel_port_slave_address,
      byteenable => HEX7_HEX4_avalon_parallel_port_slave_byteenable,
      chipselect => HEX7_HEX4_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => HEX7_HEX4_avalon_parallel_port_slave_read,
      reset => HEX7_HEX4_avalon_parallel_port_slave_reset,
      write => HEX7_HEX4_avalon_parallel_port_slave_write,
      writedata => HEX7_HEX4_avalon_parallel_port_slave_writedata
    );


  --the_Interval_Timer_s1, which is an e_instance
  the_Interval_Timer_s1 : Interval_Timer_s1_arbitrator
    port map(
      CPU_data_master_granted_Interval_Timer_s1 => CPU_data_master_granted_Interval_Timer_s1,
      CPU_data_master_qualified_request_Interval_Timer_s1 => CPU_data_master_qualified_request_Interval_Timer_s1,
      CPU_data_master_read_data_valid_Interval_Timer_s1 => CPU_data_master_read_data_valid_Interval_Timer_s1,
      CPU_data_master_requests_Interval_Timer_s1 => CPU_data_master_requests_Interval_Timer_s1,
      Interval_Timer_s1_address => Interval_Timer_s1_address,
      Interval_Timer_s1_chipselect => Interval_Timer_s1_chipselect,
      Interval_Timer_s1_irq_from_sa => Interval_Timer_s1_irq_from_sa,
      Interval_Timer_s1_readdata_from_sa => Interval_Timer_s1_readdata_from_sa,
      Interval_Timer_s1_reset_n => Interval_Timer_s1_reset_n,
      Interval_Timer_s1_write_n => Interval_Timer_s1_write_n,
      Interval_Timer_s1_writedata => Interval_Timer_s1_writedata,
      d1_Interval_Timer_s1_end_xfer => d1_Interval_Timer_s1_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Interval_Timer_s1_irq => Interval_Timer_s1_irq,
      Interval_Timer_s1_readdata => Interval_Timer_s1_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Interval_Timer, which is an e_ptf_instance
  the_Interval_Timer : Interval_Timer
    port map(
      irq => Interval_Timer_s1_irq,
      readdata => Interval_Timer_s1_readdata,
      address => Interval_Timer_s1_address,
      chipselect => Interval_Timer_s1_chipselect,
      clk => internal_sys_clk,
      reset_n => Interval_Timer_s1_reset_n,
      write_n => Interval_Timer_s1_write_n,
      writedata => Interval_Timer_s1_writedata
    );


  --the_JTAG_UART_avalon_jtag_slave, which is an e_instance
  the_JTAG_UART_avalon_jtag_slave : JTAG_UART_avalon_jtag_slave_arbitrator
    port map(
      CPU_data_master_granted_JTAG_UART_avalon_jtag_slave => CPU_data_master_granted_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave => CPU_data_master_qualified_request_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave => CPU_data_master_read_data_valid_JTAG_UART_avalon_jtag_slave,
      CPU_data_master_requests_JTAG_UART_avalon_jtag_slave => CPU_data_master_requests_JTAG_UART_avalon_jtag_slave,
      JTAG_UART_avalon_jtag_slave_address => JTAG_UART_avalon_jtag_slave_address,
      JTAG_UART_avalon_jtag_slave_chipselect => JTAG_UART_avalon_jtag_slave_chipselect,
      JTAG_UART_avalon_jtag_slave_dataavailable_from_sa => JTAG_UART_avalon_jtag_slave_dataavailable_from_sa,
      JTAG_UART_avalon_jtag_slave_irq_from_sa => JTAG_UART_avalon_jtag_slave_irq_from_sa,
      JTAG_UART_avalon_jtag_slave_read_n => JTAG_UART_avalon_jtag_slave_read_n,
      JTAG_UART_avalon_jtag_slave_readdata_from_sa => JTAG_UART_avalon_jtag_slave_readdata_from_sa,
      JTAG_UART_avalon_jtag_slave_readyfordata_from_sa => JTAG_UART_avalon_jtag_slave_readyfordata_from_sa,
      JTAG_UART_avalon_jtag_slave_reset_n => JTAG_UART_avalon_jtag_slave_reset_n,
      JTAG_UART_avalon_jtag_slave_waitrequest_from_sa => JTAG_UART_avalon_jtag_slave_waitrequest_from_sa,
      JTAG_UART_avalon_jtag_slave_write_n => JTAG_UART_avalon_jtag_slave_write_n,
      JTAG_UART_avalon_jtag_slave_writedata => JTAG_UART_avalon_jtag_slave_writedata,
      d1_JTAG_UART_avalon_jtag_slave_end_xfer => d1_JTAG_UART_avalon_jtag_slave_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      JTAG_UART_avalon_jtag_slave_dataavailable => JTAG_UART_avalon_jtag_slave_dataavailable,
      JTAG_UART_avalon_jtag_slave_irq => JTAG_UART_avalon_jtag_slave_irq,
      JTAG_UART_avalon_jtag_slave_readdata => JTAG_UART_avalon_jtag_slave_readdata,
      JTAG_UART_avalon_jtag_slave_readyfordata => JTAG_UART_avalon_jtag_slave_readyfordata,
      JTAG_UART_avalon_jtag_slave_waitrequest => JTAG_UART_avalon_jtag_slave_waitrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_JTAG_UART, which is an e_ptf_instance
  the_JTAG_UART : JTAG_UART
    port map(
      av_irq => JTAG_UART_avalon_jtag_slave_irq,
      av_readdata => JTAG_UART_avalon_jtag_slave_readdata,
      av_waitrequest => JTAG_UART_avalon_jtag_slave_waitrequest,
      dataavailable => JTAG_UART_avalon_jtag_slave_dataavailable,
      readyfordata => JTAG_UART_avalon_jtag_slave_readyfordata,
      av_address => JTAG_UART_avalon_jtag_slave_address,
      av_chipselect => JTAG_UART_avalon_jtag_slave_chipselect,
      av_read_n => JTAG_UART_avalon_jtag_slave_read_n,
      av_write_n => JTAG_UART_avalon_jtag_slave_write_n,
      av_writedata => JTAG_UART_avalon_jtag_slave_writedata,
      clk => internal_sys_clk,
      rst_n => JTAG_UART_avalon_jtag_slave_reset_n
    );


  --the_PS2_Port_avalon_ps2_slave, which is an e_instance
  the_PS2_Port_avalon_ps2_slave : PS2_Port_avalon_ps2_slave_arbitrator
    port map(
      CPU_data_master_granted_PS2_Port_avalon_ps2_slave => CPU_data_master_granted_PS2_Port_avalon_ps2_slave,
      CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave => CPU_data_master_qualified_request_PS2_Port_avalon_ps2_slave,
      CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave => CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave,
      CPU_data_master_requests_PS2_Port_avalon_ps2_slave => CPU_data_master_requests_PS2_Port_avalon_ps2_slave,
      PS2_Port_avalon_ps2_slave_address => PS2_Port_avalon_ps2_slave_address,
      PS2_Port_avalon_ps2_slave_byteenable => PS2_Port_avalon_ps2_slave_byteenable,
      PS2_Port_avalon_ps2_slave_chipselect => PS2_Port_avalon_ps2_slave_chipselect,
      PS2_Port_avalon_ps2_slave_irq_from_sa => PS2_Port_avalon_ps2_slave_irq_from_sa,
      PS2_Port_avalon_ps2_slave_read => PS2_Port_avalon_ps2_slave_read,
      PS2_Port_avalon_ps2_slave_readdata_from_sa => PS2_Port_avalon_ps2_slave_readdata_from_sa,
      PS2_Port_avalon_ps2_slave_reset => PS2_Port_avalon_ps2_slave_reset,
      PS2_Port_avalon_ps2_slave_waitrequest_from_sa => PS2_Port_avalon_ps2_slave_waitrequest_from_sa,
      PS2_Port_avalon_ps2_slave_write => PS2_Port_avalon_ps2_slave_write,
      PS2_Port_avalon_ps2_slave_writedata => PS2_Port_avalon_ps2_slave_writedata,
      d1_PS2_Port_avalon_ps2_slave_end_xfer => d1_PS2_Port_avalon_ps2_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave => registered_CPU_data_master_read_data_valid_PS2_Port_avalon_ps2_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      PS2_Port_avalon_ps2_slave_irq => PS2_Port_avalon_ps2_slave_irq,
      PS2_Port_avalon_ps2_slave_readdata => PS2_Port_avalon_ps2_slave_readdata,
      PS2_Port_avalon_ps2_slave_waitrequest => PS2_Port_avalon_ps2_slave_waitrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_PS2_Port, which is an e_ptf_instance
  the_PS2_Port : PS2_Port
    port map(
      PS2_CLK => PS2_CLK_to_and_from_the_PS2_Port,
      PS2_DAT => PS2_DAT_to_and_from_the_PS2_Port,
      irq => PS2_Port_avalon_ps2_slave_irq,
      readdata => PS2_Port_avalon_ps2_slave_readdata,
      waitrequest => PS2_Port_avalon_ps2_slave_waitrequest,
      address => PS2_Port_avalon_ps2_slave_address,
      byteenable => PS2_Port_avalon_ps2_slave_byteenable,
      chipselect => PS2_Port_avalon_ps2_slave_chipselect,
      clk => internal_sys_clk,
      read => PS2_Port_avalon_ps2_slave_read,
      reset => PS2_Port_avalon_ps2_slave_reset,
      write => PS2_Port_avalon_ps2_slave_write,
      writedata => PS2_Port_avalon_ps2_slave_writedata
    );


  --the_Pushbuttons_avalon_parallel_port_slave, which is an e_instance
  the_Pushbuttons_avalon_parallel_port_slave : Pushbuttons_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_granted_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_qualified_request_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave => CPU_data_master_requests_Pushbuttons_avalon_parallel_port_slave,
      Pushbuttons_avalon_parallel_port_slave_address => Pushbuttons_avalon_parallel_port_slave_address,
      Pushbuttons_avalon_parallel_port_slave_byteenable => Pushbuttons_avalon_parallel_port_slave_byteenable,
      Pushbuttons_avalon_parallel_port_slave_chipselect => Pushbuttons_avalon_parallel_port_slave_chipselect,
      Pushbuttons_avalon_parallel_port_slave_irq_from_sa => Pushbuttons_avalon_parallel_port_slave_irq_from_sa,
      Pushbuttons_avalon_parallel_port_slave_read => Pushbuttons_avalon_parallel_port_slave_read,
      Pushbuttons_avalon_parallel_port_slave_readdata_from_sa => Pushbuttons_avalon_parallel_port_slave_readdata_from_sa,
      Pushbuttons_avalon_parallel_port_slave_reset => Pushbuttons_avalon_parallel_port_slave_reset,
      Pushbuttons_avalon_parallel_port_slave_write => Pushbuttons_avalon_parallel_port_slave_write,
      Pushbuttons_avalon_parallel_port_slave_writedata => Pushbuttons_avalon_parallel_port_slave_writedata,
      d1_Pushbuttons_avalon_parallel_port_slave_end_xfer => d1_Pushbuttons_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Pushbuttons_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Pushbuttons_avalon_parallel_port_slave_irq => Pushbuttons_avalon_parallel_port_slave_irq,
      Pushbuttons_avalon_parallel_port_slave_readdata => Pushbuttons_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Pushbuttons, which is an e_ptf_instance
  the_Pushbuttons : Pushbuttons
    port map(
      irq => Pushbuttons_avalon_parallel_port_slave_irq,
      readdata => Pushbuttons_avalon_parallel_port_slave_readdata,
      KEY => KEY_to_the_Pushbuttons,
      address => Pushbuttons_avalon_parallel_port_slave_address,
      byteenable => Pushbuttons_avalon_parallel_port_slave_byteenable,
      chipselect => Pushbuttons_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Pushbuttons_avalon_parallel_port_slave_read,
      reset => Pushbuttons_avalon_parallel_port_slave_reset,
      write => Pushbuttons_avalon_parallel_port_slave_write,
      writedata => Pushbuttons_avalon_parallel_port_slave_writedata
    );


  --the_Red_LEDs_avalon_parallel_port_slave, which is an e_instance
  the_Red_LEDs_avalon_parallel_port_slave : Red_LEDs_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_granted_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_qualified_request_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave => CPU_data_master_requests_Red_LEDs_avalon_parallel_port_slave,
      Red_LEDs_avalon_parallel_port_slave_address => Red_LEDs_avalon_parallel_port_slave_address,
      Red_LEDs_avalon_parallel_port_slave_byteenable => Red_LEDs_avalon_parallel_port_slave_byteenable,
      Red_LEDs_avalon_parallel_port_slave_chipselect => Red_LEDs_avalon_parallel_port_slave_chipselect,
      Red_LEDs_avalon_parallel_port_slave_read => Red_LEDs_avalon_parallel_port_slave_read,
      Red_LEDs_avalon_parallel_port_slave_readdata_from_sa => Red_LEDs_avalon_parallel_port_slave_readdata_from_sa,
      Red_LEDs_avalon_parallel_port_slave_reset => Red_LEDs_avalon_parallel_port_slave_reset,
      Red_LEDs_avalon_parallel_port_slave_write => Red_LEDs_avalon_parallel_port_slave_write,
      Red_LEDs_avalon_parallel_port_slave_writedata => Red_LEDs_avalon_parallel_port_slave_writedata,
      d1_Red_LEDs_avalon_parallel_port_slave_end_xfer => d1_Red_LEDs_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Red_LEDs_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Red_LEDs_avalon_parallel_port_slave_readdata => Red_LEDs_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Red_LEDs, which is an e_ptf_instance
  the_Red_LEDs : Red_LEDs
    port map(
      LEDR => internal_LEDR_from_the_Red_LEDs,
      readdata => Red_LEDs_avalon_parallel_port_slave_readdata,
      address => Red_LEDs_avalon_parallel_port_slave_address,
      byteenable => Red_LEDs_avalon_parallel_port_slave_byteenable,
      chipselect => Red_LEDs_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Red_LEDs_avalon_parallel_port_slave_read,
      reset => Red_LEDs_avalon_parallel_port_slave_reset,
      write => Red_LEDs_avalon_parallel_port_slave_write,
      writedata => Red_LEDs_avalon_parallel_port_slave_writedata
    );


  --the_SDRAM_s1, which is an e_instance
  the_SDRAM_s1 : SDRAM_s1_arbitrator
    port map(
      CPU_data_master_byteenable_SDRAM_s1 => CPU_data_master_byteenable_SDRAM_s1,
      CPU_data_master_granted_SDRAM_s1 => CPU_data_master_granted_SDRAM_s1,
      CPU_data_master_qualified_request_SDRAM_s1 => CPU_data_master_qualified_request_SDRAM_s1,
      CPU_data_master_read_data_valid_SDRAM_s1 => CPU_data_master_read_data_valid_SDRAM_s1,
      CPU_data_master_read_data_valid_SDRAM_s1_shift_register => CPU_data_master_read_data_valid_SDRAM_s1_shift_register,
      CPU_data_master_requests_SDRAM_s1 => CPU_data_master_requests_SDRAM_s1,
      CPU_instruction_master_granted_SDRAM_s1 => CPU_instruction_master_granted_SDRAM_s1,
      CPU_instruction_master_qualified_request_SDRAM_s1 => CPU_instruction_master_qualified_request_SDRAM_s1,
      CPU_instruction_master_read_data_valid_SDRAM_s1 => CPU_instruction_master_read_data_valid_SDRAM_s1,
      CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register => CPU_instruction_master_read_data_valid_SDRAM_s1_shift_register,
      CPU_instruction_master_requests_SDRAM_s1 => CPU_instruction_master_requests_SDRAM_s1,
      SDRAM_s1_address => SDRAM_s1_address,
      SDRAM_s1_byteenable_n => SDRAM_s1_byteenable_n,
      SDRAM_s1_chipselect => SDRAM_s1_chipselect,
      SDRAM_s1_read_n => SDRAM_s1_read_n,
      SDRAM_s1_readdata_from_sa => SDRAM_s1_readdata_from_sa,
      SDRAM_s1_reset_n => SDRAM_s1_reset_n,
      SDRAM_s1_waitrequest_from_sa => SDRAM_s1_waitrequest_from_sa,
      SDRAM_s1_write_n => SDRAM_s1_write_n,
      SDRAM_s1_writedata => SDRAM_s1_writedata,
      d1_SDRAM_s1_end_xfer => d1_SDRAM_s1_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_16 => CPU_data_master_dbs_write_16,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_instruction_master_address_to_slave => CPU_instruction_master_address_to_slave,
      CPU_instruction_master_dbs_address => CPU_instruction_master_dbs_address,
      CPU_instruction_master_latency_counter => CPU_instruction_master_latency_counter,
      CPU_instruction_master_read => CPU_instruction_master_read,
      SDRAM_s1_readdata => SDRAM_s1_readdata,
      SDRAM_s1_readdatavalid => SDRAM_s1_readdatavalid,
      SDRAM_s1_waitrequest => SDRAM_s1_waitrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_SDRAM, which is an e_ptf_instance
  the_SDRAM : SDRAM
    port map(
      za_data => SDRAM_s1_readdata,
      za_valid => SDRAM_s1_readdatavalid,
      za_waitrequest => SDRAM_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_SDRAM,
      zs_ba => internal_zs_ba_from_the_SDRAM,
      zs_cas_n => internal_zs_cas_n_from_the_SDRAM,
      zs_cke => internal_zs_cke_from_the_SDRAM,
      zs_cs_n => internal_zs_cs_n_from_the_SDRAM,
      zs_dq => zs_dq_to_and_from_the_SDRAM,
      zs_dqm => internal_zs_dqm_from_the_SDRAM,
      zs_ras_n => internal_zs_ras_n_from_the_SDRAM,
      zs_we_n => internal_zs_we_n_from_the_SDRAM,
      az_addr => SDRAM_s1_address,
      az_be_n => SDRAM_s1_byteenable_n,
      az_cs => SDRAM_s1_chipselect,
      az_data => SDRAM_s1_writedata,
      az_rd_n => SDRAM_s1_read_n,
      az_wr_n => SDRAM_s1_write_n,
      clk => internal_sys_clk,
      reset_n => SDRAM_s1_reset_n
    );


  --the_SRAM_avalon_sram_slave, which is an e_instance
  the_SRAM_avalon_sram_slave : SRAM_avalon_sram_slave_arbitrator
    port map(
      CPU_data_master_byteenable_SRAM_avalon_sram_slave => CPU_data_master_byteenable_SRAM_avalon_sram_slave,
      CPU_data_master_granted_SRAM_avalon_sram_slave => CPU_data_master_granted_SRAM_avalon_sram_slave,
      CPU_data_master_qualified_request_SRAM_avalon_sram_slave => CPU_data_master_qualified_request_SRAM_avalon_sram_slave,
      CPU_data_master_read_data_valid_SRAM_avalon_sram_slave => CPU_data_master_read_data_valid_SRAM_avalon_sram_slave,
      CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register => CPU_data_master_read_data_valid_SRAM_avalon_sram_slave_shift_register,
      CPU_data_master_requests_SRAM_avalon_sram_slave => CPU_data_master_requests_SRAM_avalon_sram_slave,
      SRAM_avalon_sram_slave_address => SRAM_avalon_sram_slave_address,
      SRAM_avalon_sram_slave_byteenable => SRAM_avalon_sram_slave_byteenable,
      SRAM_avalon_sram_slave_read => SRAM_avalon_sram_slave_read,
      SRAM_avalon_sram_slave_readdata_from_sa => SRAM_avalon_sram_slave_readdata_from_sa,
      SRAM_avalon_sram_slave_reset => SRAM_avalon_sram_slave_reset,
      SRAM_avalon_sram_slave_write => SRAM_avalon_sram_slave_write,
      SRAM_avalon_sram_slave_writedata => SRAM_avalon_sram_slave_writedata,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register => VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave,
      d1_SRAM_avalon_sram_slave_end_xfer => d1_SRAM_avalon_sram_slave_end_xfer,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_16 => CPU_data_master_dbs_write_16,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      SRAM_avalon_sram_slave_readdata => SRAM_avalon_sram_slave_readdata,
      SRAM_avalon_sram_slave_readdatavalid => SRAM_avalon_sram_slave_readdatavalid,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock => VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter => VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read => VGA_Pixel_Buffer_avalon_pixel_dma_master_read,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_SRAM, which is an e_ptf_instance
  the_SRAM : SRAM
    port map(
      SRAM_ADDR => internal_SRAM_ADDR_from_the_SRAM,
      SRAM_CE_N => internal_SRAM_CE_N_from_the_SRAM,
      SRAM_DQ => SRAM_DQ_to_and_from_the_SRAM,
      SRAM_LB_N => internal_SRAM_LB_N_from_the_SRAM,
      SRAM_OE_N => internal_SRAM_OE_N_from_the_SRAM,
      SRAM_UB_N => internal_SRAM_UB_N_from_the_SRAM,
      SRAM_WE_N => internal_SRAM_WE_N_from_the_SRAM,
      readdata => SRAM_avalon_sram_slave_readdata,
      readdatavalid => SRAM_avalon_sram_slave_readdatavalid,
      address => SRAM_avalon_sram_slave_address,
      byteenable => SRAM_avalon_sram_slave_byteenable,
      clk => internal_sys_clk,
      read => SRAM_avalon_sram_slave_read,
      reset => SRAM_avalon_sram_slave_reset,
      write => SRAM_avalon_sram_slave_write,
      writedata => SRAM_avalon_sram_slave_writedata
    );


  --the_Serial_Port_avalon_rs232_slave, which is an e_instance
  the_Serial_Port_avalon_rs232_slave : Serial_Port_avalon_rs232_slave_arbitrator
    port map(
      CPU_data_master_granted_Serial_Port_avalon_rs232_slave => CPU_data_master_granted_Serial_Port_avalon_rs232_slave,
      CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave => CPU_data_master_qualified_request_Serial_Port_avalon_rs232_slave,
      CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave => CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave,
      CPU_data_master_requests_Serial_Port_avalon_rs232_slave => CPU_data_master_requests_Serial_Port_avalon_rs232_slave,
      Serial_Port_avalon_rs232_slave_address => Serial_Port_avalon_rs232_slave_address,
      Serial_Port_avalon_rs232_slave_byteenable => Serial_Port_avalon_rs232_slave_byteenable,
      Serial_Port_avalon_rs232_slave_chipselect => Serial_Port_avalon_rs232_slave_chipselect,
      Serial_Port_avalon_rs232_slave_irq_from_sa => Serial_Port_avalon_rs232_slave_irq_from_sa,
      Serial_Port_avalon_rs232_slave_read => Serial_Port_avalon_rs232_slave_read,
      Serial_Port_avalon_rs232_slave_readdata_from_sa => Serial_Port_avalon_rs232_slave_readdata_from_sa,
      Serial_Port_avalon_rs232_slave_reset => Serial_Port_avalon_rs232_slave_reset,
      Serial_Port_avalon_rs232_slave_write => Serial_Port_avalon_rs232_slave_write,
      Serial_Port_avalon_rs232_slave_writedata => Serial_Port_avalon_rs232_slave_writedata,
      d1_Serial_Port_avalon_rs232_slave_end_xfer => d1_Serial_Port_avalon_rs232_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave => registered_CPU_data_master_read_data_valid_Serial_Port_avalon_rs232_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Serial_Port_avalon_rs232_slave_irq => Serial_Port_avalon_rs232_slave_irq,
      Serial_Port_avalon_rs232_slave_readdata => Serial_Port_avalon_rs232_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Serial_Port, which is an e_ptf_instance
  the_Serial_Port : Serial_Port
    port map(
      UART_TXD => internal_UART_TXD_from_the_Serial_Port,
      irq => Serial_Port_avalon_rs232_slave_irq,
      readdata => Serial_Port_avalon_rs232_slave_readdata,
      UART_RXD => UART_RXD_to_the_Serial_Port,
      address => Serial_Port_avalon_rs232_slave_address,
      byteenable => Serial_Port_avalon_rs232_slave_byteenable,
      chipselect => Serial_Port_avalon_rs232_slave_chipselect,
      clk => internal_sys_clk,
      read => Serial_Port_avalon_rs232_slave_read,
      reset => Serial_Port_avalon_rs232_slave_reset,
      write => Serial_Port_avalon_rs232_slave_write,
      writedata => Serial_Port_avalon_rs232_slave_writedata
    );


  --the_Slider_Switches_avalon_parallel_port_slave, which is an e_instance
  the_Slider_Switches_avalon_parallel_port_slave : Slider_Switches_avalon_parallel_port_slave_arbitrator
    port map(
      CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_granted_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_qualified_request_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave => CPU_data_master_requests_Slider_Switches_avalon_parallel_port_slave,
      Slider_Switches_avalon_parallel_port_slave_address => Slider_Switches_avalon_parallel_port_slave_address,
      Slider_Switches_avalon_parallel_port_slave_byteenable => Slider_Switches_avalon_parallel_port_slave_byteenable,
      Slider_Switches_avalon_parallel_port_slave_chipselect => Slider_Switches_avalon_parallel_port_slave_chipselect,
      Slider_Switches_avalon_parallel_port_slave_read => Slider_Switches_avalon_parallel_port_slave_read,
      Slider_Switches_avalon_parallel_port_slave_readdata_from_sa => Slider_Switches_avalon_parallel_port_slave_readdata_from_sa,
      Slider_Switches_avalon_parallel_port_slave_reset => Slider_Switches_avalon_parallel_port_slave_reset,
      Slider_Switches_avalon_parallel_port_slave_write => Slider_Switches_avalon_parallel_port_slave_write,
      Slider_Switches_avalon_parallel_port_slave_writedata => Slider_Switches_avalon_parallel_port_slave_writedata,
      d1_Slider_Switches_avalon_parallel_port_slave_end_xfer => d1_Slider_Switches_avalon_parallel_port_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave => registered_CPU_data_master_read_data_valid_Slider_Switches_avalon_parallel_port_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      Slider_Switches_avalon_parallel_port_slave_readdata => Slider_Switches_avalon_parallel_port_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_Slider_Switches, which is an e_ptf_instance
  the_Slider_Switches : Slider_Switches
    port map(
      readdata => Slider_Switches_avalon_parallel_port_slave_readdata,
      SW => SW_to_the_Slider_Switches,
      address => Slider_Switches_avalon_parallel_port_slave_address,
      byteenable => Slider_Switches_avalon_parallel_port_slave_byteenable,
      chipselect => Slider_Switches_avalon_parallel_port_slave_chipselect,
      clk => internal_sys_clk,
      read => Slider_Switches_avalon_parallel_port_slave_read,
      reset => Slider_Switches_avalon_parallel_port_slave_reset,
      write => Slider_Switches_avalon_parallel_port_slave_write,
      writedata => Slider_Switches_avalon_parallel_port_slave_writedata
    );


  --the_VGA_Char_Buffer_avalon_char_buffer_slave, which is an e_instance
  the_VGA_Char_Buffer_avalon_char_buffer_slave : VGA_Char_Buffer_avalon_char_buffer_slave_arbitrator
    port map(
      CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_byteenable_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_granted_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave => CPU_data_master_requests_VGA_Char_Buffer_avalon_char_buffer_slave,
      VGA_Char_Buffer_avalon_char_buffer_slave_address => VGA_Char_Buffer_avalon_char_buffer_slave_address,
      VGA_Char_Buffer_avalon_char_buffer_slave_byteenable => VGA_Char_Buffer_avalon_char_buffer_slave_byteenable,
      VGA_Char_Buffer_avalon_char_buffer_slave_chipselect => VGA_Char_Buffer_avalon_char_buffer_slave_chipselect,
      VGA_Char_Buffer_avalon_char_buffer_slave_read => VGA_Char_Buffer_avalon_char_buffer_slave_read,
      VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa => VGA_Char_Buffer_avalon_char_buffer_slave_readdata_from_sa,
      VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa => VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest_from_sa,
      VGA_Char_Buffer_avalon_char_buffer_slave_write => VGA_Char_Buffer_avalon_char_buffer_slave_write,
      VGA_Char_Buffer_avalon_char_buffer_slave_writedata => VGA_Char_Buffer_avalon_char_buffer_slave_writedata,
      d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer => d1_VGA_Char_Buffer_avalon_char_buffer_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave => registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_buffer_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_8 => CPU_data_master_dbs_write_8,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      VGA_Char_Buffer_avalon_char_buffer_slave_readdata => VGA_Char_Buffer_avalon_char_buffer_slave_readdata,
      VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest => VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Char_Buffer_avalon_char_control_slave, which is an e_instance
  the_VGA_Char_Buffer_avalon_char_control_slave : VGA_Char_Buffer_avalon_char_control_slave_arbitrator
    port map(
      CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_granted_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_qualified_request_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave => CPU_data_master_requests_VGA_Char_Buffer_avalon_char_control_slave,
      VGA_Char_Buffer_avalon_char_control_slave_address => VGA_Char_Buffer_avalon_char_control_slave_address,
      VGA_Char_Buffer_avalon_char_control_slave_byteenable => VGA_Char_Buffer_avalon_char_control_slave_byteenable,
      VGA_Char_Buffer_avalon_char_control_slave_chipselect => VGA_Char_Buffer_avalon_char_control_slave_chipselect,
      VGA_Char_Buffer_avalon_char_control_slave_read => VGA_Char_Buffer_avalon_char_control_slave_read,
      VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa => VGA_Char_Buffer_avalon_char_control_slave_readdata_from_sa,
      VGA_Char_Buffer_avalon_char_control_slave_reset => VGA_Char_Buffer_avalon_char_control_slave_reset,
      VGA_Char_Buffer_avalon_char_control_slave_write => VGA_Char_Buffer_avalon_char_control_slave_write,
      VGA_Char_Buffer_avalon_char_control_slave_writedata => VGA_Char_Buffer_avalon_char_control_slave_writedata,
      d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer => d1_VGA_Char_Buffer_avalon_char_control_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave => registered_CPU_data_master_read_data_valid_VGA_Char_Buffer_avalon_char_control_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      VGA_Char_Buffer_avalon_char_control_slave_readdata => VGA_Char_Buffer_avalon_char_control_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Char_Buffer_avalon_char_source, which is an e_instance
  the_VGA_Char_Buffer_avalon_char_source : VGA_Char_Buffer_avalon_char_source_arbitrator
    port map(
      VGA_Char_Buffer_avalon_char_source_ready => VGA_Char_Buffer_avalon_char_source_ready,
      Alpha_Blending_avalon_foreground_sink_ready_from_sa => Alpha_Blending_avalon_foreground_sink_ready_from_sa,
      VGA_Char_Buffer_avalon_char_source_data => VGA_Char_Buffer_avalon_char_source_data,
      VGA_Char_Buffer_avalon_char_source_endofpacket => VGA_Char_Buffer_avalon_char_source_endofpacket,
      VGA_Char_Buffer_avalon_char_source_startofpacket => VGA_Char_Buffer_avalon_char_source_startofpacket,
      VGA_Char_Buffer_avalon_char_source_valid => VGA_Char_Buffer_avalon_char_source_valid,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Char_Buffer, which is an e_ptf_instance
  the_VGA_Char_Buffer : VGA_Char_Buffer
    port map(
      buf_readdata => VGA_Char_Buffer_avalon_char_buffer_slave_readdata,
      buf_waitrequest => VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest,
      ctrl_readdata => VGA_Char_Buffer_avalon_char_control_slave_readdata,
      stream_data => VGA_Char_Buffer_avalon_char_source_data,
      stream_endofpacket => VGA_Char_Buffer_avalon_char_source_endofpacket,
      stream_startofpacket => VGA_Char_Buffer_avalon_char_source_startofpacket,
      stream_valid => VGA_Char_Buffer_avalon_char_source_valid,
      buf_address => VGA_Char_Buffer_avalon_char_buffer_slave_address,
      buf_byteenable => VGA_Char_Buffer_avalon_char_buffer_slave_byteenable,
      buf_chipselect => VGA_Char_Buffer_avalon_char_buffer_slave_chipselect,
      buf_read => VGA_Char_Buffer_avalon_char_buffer_slave_read,
      buf_write => VGA_Char_Buffer_avalon_char_buffer_slave_write,
      buf_writedata => VGA_Char_Buffer_avalon_char_buffer_slave_writedata,
      clk => internal_sys_clk,
      ctrl_address => VGA_Char_Buffer_avalon_char_control_slave_address,
      ctrl_byteenable => VGA_Char_Buffer_avalon_char_control_slave_byteenable,
      ctrl_chipselect => VGA_Char_Buffer_avalon_char_control_slave_chipselect,
      ctrl_read => VGA_Char_Buffer_avalon_char_control_slave_read,
      ctrl_write => VGA_Char_Buffer_avalon_char_control_slave_write,
      ctrl_writedata => VGA_Char_Buffer_avalon_char_control_slave_writedata,
      reset => VGA_Char_Buffer_avalon_char_control_slave_reset,
      stream_ready => VGA_Char_Buffer_avalon_char_source_ready
    );


  --the_VGA_Controller_avalon_vga_sink, which is an e_instance
  the_VGA_Controller_avalon_vga_sink : VGA_Controller_avalon_vga_sink_arbitrator
    port map(
      VGA_Controller_avalon_vga_sink_data => VGA_Controller_avalon_vga_sink_data,
      VGA_Controller_avalon_vga_sink_endofpacket => VGA_Controller_avalon_vga_sink_endofpacket,
      VGA_Controller_avalon_vga_sink_ready_from_sa => VGA_Controller_avalon_vga_sink_ready_from_sa,
      VGA_Controller_avalon_vga_sink_reset => VGA_Controller_avalon_vga_sink_reset,
      VGA_Controller_avalon_vga_sink_startofpacket => VGA_Controller_avalon_vga_sink_startofpacket,
      VGA_Controller_avalon_vga_sink_valid => VGA_Controller_avalon_vga_sink_valid,
      VGA_Controller_avalon_vga_sink_ready => VGA_Controller_avalon_vga_sink_ready,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid,
      clk => internal_vga_clk,
      reset_n => vga_clk_reset_n
    );


  --the_VGA_Controller, which is an e_ptf_instance
  the_VGA_Controller : VGA_Controller
    port map(
      VGA_B => internal_VGA_B_from_the_VGA_Controller,
      VGA_BLANK => internal_VGA_BLANK_from_the_VGA_Controller,
      VGA_CLK => internal_VGA_CLK_from_the_VGA_Controller,
      VGA_G => internal_VGA_G_from_the_VGA_Controller,
      VGA_HS => internal_VGA_HS_from_the_VGA_Controller,
      VGA_R => internal_VGA_R_from_the_VGA_Controller,
      VGA_SYNC => internal_VGA_SYNC_from_the_VGA_Controller,
      VGA_VS => internal_VGA_VS_from_the_VGA_Controller,
      ready => VGA_Controller_avalon_vga_sink_ready,
      clk => internal_vga_clk,
      data => VGA_Controller_avalon_vga_sink_data,
      endofpacket => VGA_Controller_avalon_vga_sink_endofpacket,
      reset => VGA_Controller_avalon_vga_sink_reset,
      startofpacket => VGA_Controller_avalon_vga_sink_startofpacket,
      valid => VGA_Controller_avalon_vga_sink_valid
    );


  --the_VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink, which is an e_instance
  the_VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink : VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_arbitrator
    port map(
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready_from_sa,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid,
      Alpha_Blending_avalon_blended_source_data => Alpha_Blending_avalon_blended_source_data,
      Alpha_Blending_avalon_blended_source_endofpacket => Alpha_Blending_avalon_blended_source_endofpacket,
      Alpha_Blending_avalon_blended_source_startofpacket => Alpha_Blending_avalon_blended_source_startofpacket,
      Alpha_Blending_avalon_blended_source_valid => Alpha_Blending_avalon_blended_source_valid,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Dual_Clock_FIFO_avalon_dc_buffer_source, which is an e_instance
  the_VGA_Dual_Clock_FIFO_avalon_dc_buffer_source : VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_arbitrator
    port map(
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready,
      VGA_Controller_avalon_vga_sink_ready_from_sa => VGA_Controller_avalon_vga_sink_ready_from_sa,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket,
      VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid,
      clk => internal_vga_clk,
      reset_n => vga_clk_reset_n
    );


  --the_VGA_Dual_Clock_FIFO, which is an e_ptf_instance
  the_VGA_Dual_Clock_FIFO : VGA_Dual_Clock_FIFO
    port map(
      stream_in_ready => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_ready,
      stream_out_data => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_data,
      stream_out_endofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_endofpacket,
      stream_out_startofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_startofpacket,
      stream_out_valid => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_valid,
      clk_stream_in => internal_sys_clk,
      clk_stream_out => internal_vga_clk,
      stream_in_data => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_data,
      stream_in_endofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_endofpacket,
      stream_in_startofpacket => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_startofpacket,
      stream_in_valid => VGA_Dual_Clock_FIFO_avalon_dc_buffer_sink_valid,
      stream_out_ready => VGA_Dual_Clock_FIFO_avalon_dc_buffer_source_ready
    );


  --the_VGA_Pixel_Buffer_avalon_control_slave, which is an e_instance
  the_VGA_Pixel_Buffer_avalon_control_slave : VGA_Pixel_Buffer_avalon_control_slave_arbitrator
    port map(
      CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_granted_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_qualified_request_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave => CPU_data_master_requests_VGA_Pixel_Buffer_avalon_control_slave,
      VGA_Pixel_Buffer_avalon_control_slave_address => VGA_Pixel_Buffer_avalon_control_slave_address,
      VGA_Pixel_Buffer_avalon_control_slave_byteenable => VGA_Pixel_Buffer_avalon_control_slave_byteenable,
      VGA_Pixel_Buffer_avalon_control_slave_read => VGA_Pixel_Buffer_avalon_control_slave_read,
      VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa => VGA_Pixel_Buffer_avalon_control_slave_readdata_from_sa,
      VGA_Pixel_Buffer_avalon_control_slave_write => VGA_Pixel_Buffer_avalon_control_slave_write,
      VGA_Pixel_Buffer_avalon_control_slave_writedata => VGA_Pixel_Buffer_avalon_control_slave_writedata,
      d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer => d1_VGA_Pixel_Buffer_avalon_control_slave_end_xfer,
      registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave => registered_CPU_data_master_read_data_valid_VGA_Pixel_Buffer_avalon_control_slave,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      CPU_data_master_writedata => CPU_data_master_writedata,
      VGA_Pixel_Buffer_avalon_control_slave_readdata => VGA_Pixel_Buffer_avalon_control_slave_readdata,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_Buffer_avalon_pixel_dma_master, which is an e_instance
  the_VGA_Pixel_Buffer_avalon_pixel_dma_master : VGA_Pixel_Buffer_avalon_pixel_dma_master_arbitrator
    port map(
      VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_address_to_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter => VGA_Pixel_Buffer_avalon_pixel_dma_master_latency_counter,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata => VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid => VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_reset => VGA_Pixel_Buffer_avalon_pixel_dma_master_reset,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest => VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest,
      SRAM_avalon_sram_slave_readdata_from_sa => SRAM_avalon_sram_slave_readdata_from_sa,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_address => VGA_Pixel_Buffer_avalon_pixel_dma_master_address,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_granted_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_qualified_request_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read => VGA_Pixel_Buffer_avalon_pixel_dma_master_read,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register => VGA_Pixel_Buffer_avalon_pixel_dma_master_read_data_valid_SRAM_avalon_sram_slave_shift_register,
      VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave => VGA_Pixel_Buffer_avalon_pixel_dma_master_requests_SRAM_avalon_sram_slave,
      clk => internal_sys_clk,
      d1_SRAM_avalon_sram_slave_end_xfer => d1_SRAM_avalon_sram_slave_end_xfer,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_Buffer_avalon_pixel_source, which is an e_instance
  the_VGA_Pixel_Buffer_avalon_pixel_source : VGA_Pixel_Buffer_avalon_pixel_source_arbitrator
    port map(
      VGA_Pixel_Buffer_avalon_pixel_source_ready => VGA_Pixel_Buffer_avalon_pixel_source_ready,
      VGA_Pixel_Buffer_avalon_pixel_source_data => VGA_Pixel_Buffer_avalon_pixel_source_data,
      VGA_Pixel_Buffer_avalon_pixel_source_endofpacket => VGA_Pixel_Buffer_avalon_pixel_source_endofpacket,
      VGA_Pixel_Buffer_avalon_pixel_source_startofpacket => VGA_Pixel_Buffer_avalon_pixel_source_startofpacket,
      VGA_Pixel_Buffer_avalon_pixel_source_valid => VGA_Pixel_Buffer_avalon_pixel_source_valid,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_Buffer, which is an e_ptf_instance
  the_VGA_Pixel_Buffer : VGA_Pixel_Buffer
    port map(
      master_address => VGA_Pixel_Buffer_avalon_pixel_dma_master_address,
      master_arbiterlock => VGA_Pixel_Buffer_avalon_pixel_dma_master_arbiterlock,
      master_read => VGA_Pixel_Buffer_avalon_pixel_dma_master_read,
      slave_readdata => VGA_Pixel_Buffer_avalon_control_slave_readdata,
      stream_data => VGA_Pixel_Buffer_avalon_pixel_source_data,
      stream_endofpacket => VGA_Pixel_Buffer_avalon_pixel_source_endofpacket,
      stream_startofpacket => VGA_Pixel_Buffer_avalon_pixel_source_startofpacket,
      stream_valid => VGA_Pixel_Buffer_avalon_pixel_source_valid,
      clk => internal_sys_clk,
      master_readdata => VGA_Pixel_Buffer_avalon_pixel_dma_master_readdata,
      master_readdatavalid => VGA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid,
      master_waitrequest => VGA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest,
      reset => VGA_Pixel_Buffer_avalon_pixel_dma_master_reset,
      slave_address => VGA_Pixel_Buffer_avalon_control_slave_address,
      slave_byteenable => VGA_Pixel_Buffer_avalon_control_slave_byteenable,
      slave_read => VGA_Pixel_Buffer_avalon_control_slave_read,
      slave_write => VGA_Pixel_Buffer_avalon_control_slave_write,
      slave_writedata => VGA_Pixel_Buffer_avalon_control_slave_writedata,
      stream_ready => VGA_Pixel_Buffer_avalon_pixel_source_ready
    );


  --the_VGA_Pixel_RGB_Resampler_avalon_rgb_sink, which is an e_instance
  the_VGA_Pixel_RGB_Resampler_avalon_rgb_sink : VGA_Pixel_RGB_Resampler_avalon_rgb_sink_arbitrator
    port map(
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready_from_sa,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid,
      VGA_Pixel_Buffer_avalon_pixel_source_data => VGA_Pixel_Buffer_avalon_pixel_source_data,
      VGA_Pixel_Buffer_avalon_pixel_source_endofpacket => VGA_Pixel_Buffer_avalon_pixel_source_endofpacket,
      VGA_Pixel_Buffer_avalon_pixel_source_startofpacket => VGA_Pixel_Buffer_avalon_pixel_source_startofpacket,
      VGA_Pixel_Buffer_avalon_pixel_source_valid => VGA_Pixel_Buffer_avalon_pixel_source_valid,
      VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_RGB_Resampler_avalon_rgb_source, which is an e_instance
  the_VGA_Pixel_RGB_Resampler_avalon_rgb_source : VGA_Pixel_RGB_Resampler_avalon_rgb_source_arbitrator
    port map(
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready => VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_data => VGA_Pixel_RGB_Resampler_avalon_rgb_source_data,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid => VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid,
      VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa => VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_RGB_Resampler, which is an e_ptf_instance
  the_VGA_Pixel_RGB_Resampler : VGA_Pixel_RGB_Resampler
    port map(
      stream_in_ready => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_ready,
      stream_out_data => VGA_Pixel_RGB_Resampler_avalon_rgb_source_data,
      stream_out_endofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket,
      stream_out_startofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket,
      stream_out_valid => VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid,
      clk => internal_sys_clk,
      reset => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_reset,
      stream_in_data => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_data,
      stream_in_endofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_endofpacket,
      stream_in_startofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_startofpacket,
      stream_in_valid => VGA_Pixel_RGB_Resampler_avalon_rgb_sink_valid,
      stream_out_ready => VGA_Pixel_RGB_Resampler_avalon_rgb_source_ready
    );


  --the_VGA_Pixel_Scaler_avalon_scaler_sink, which is an e_instance
  the_VGA_Pixel_Scaler_avalon_scaler_sink : VGA_Pixel_Scaler_avalon_scaler_sink_arbitrator
    port map(
      VGA_Pixel_Scaler_avalon_scaler_sink_data => VGA_Pixel_Scaler_avalon_scaler_sink_data,
      VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket => VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket,
      VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa => VGA_Pixel_Scaler_avalon_scaler_sink_ready_from_sa,
      VGA_Pixel_Scaler_avalon_scaler_sink_reset => VGA_Pixel_Scaler_avalon_scaler_sink_reset,
      VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket => VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket,
      VGA_Pixel_Scaler_avalon_scaler_sink_valid => VGA_Pixel_Scaler_avalon_scaler_sink_valid,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_data => VGA_Pixel_RGB_Resampler_avalon_rgb_source_data,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_endofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket => VGA_Pixel_RGB_Resampler_avalon_rgb_source_startofpacket,
      VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid => VGA_Pixel_RGB_Resampler_avalon_rgb_source_valid,
      VGA_Pixel_Scaler_avalon_scaler_sink_ready => VGA_Pixel_Scaler_avalon_scaler_sink_ready,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_Scaler_avalon_scaler_source, which is an e_instance
  the_VGA_Pixel_Scaler_avalon_scaler_source : VGA_Pixel_Scaler_avalon_scaler_source_arbitrator
    port map(
      VGA_Pixel_Scaler_avalon_scaler_source_ready => VGA_Pixel_Scaler_avalon_scaler_source_ready,
      Alpha_Blending_avalon_background_sink_ready_from_sa => Alpha_Blending_avalon_background_sink_ready_from_sa,
      VGA_Pixel_Scaler_avalon_scaler_source_data => VGA_Pixel_Scaler_avalon_scaler_source_data,
      VGA_Pixel_Scaler_avalon_scaler_source_endofpacket => VGA_Pixel_Scaler_avalon_scaler_source_endofpacket,
      VGA_Pixel_Scaler_avalon_scaler_source_startofpacket => VGA_Pixel_Scaler_avalon_scaler_source_startofpacket,
      VGA_Pixel_Scaler_avalon_scaler_source_valid => VGA_Pixel_Scaler_avalon_scaler_source_valid,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n
    );


  --the_VGA_Pixel_Scaler, which is an e_ptf_instance
  the_VGA_Pixel_Scaler : VGA_Pixel_Scaler
    port map(
      stream_in_ready => VGA_Pixel_Scaler_avalon_scaler_sink_ready,
      stream_out_data => VGA_Pixel_Scaler_avalon_scaler_source_data,
      stream_out_endofpacket => VGA_Pixel_Scaler_avalon_scaler_source_endofpacket,
      stream_out_startofpacket => VGA_Pixel_Scaler_avalon_scaler_source_startofpacket,
      stream_out_valid => VGA_Pixel_Scaler_avalon_scaler_source_valid,
      clk => internal_sys_clk,
      reset => VGA_Pixel_Scaler_avalon_scaler_sink_reset,
      stream_in_data => VGA_Pixel_Scaler_avalon_scaler_sink_data,
      stream_in_endofpacket => VGA_Pixel_Scaler_avalon_scaler_sink_endofpacket,
      stream_in_startofpacket => VGA_Pixel_Scaler_avalon_scaler_sink_startofpacket,
      stream_in_valid => VGA_Pixel_Scaler_avalon_scaler_sink_valid,
      stream_out_ready => VGA_Pixel_Scaler_avalon_scaler_source_ready
    );


  --the_nios_system_clock_0_in, which is an e_instance
  the_nios_system_clock_0_in : nios_system_clock_0_in_arbitrator
    port map(
      CPU_data_master_byteenable_nios_system_clock_0_in => CPU_data_master_byteenable_nios_system_clock_0_in,
      CPU_data_master_granted_nios_system_clock_0_in => CPU_data_master_granted_nios_system_clock_0_in,
      CPU_data_master_qualified_request_nios_system_clock_0_in => CPU_data_master_qualified_request_nios_system_clock_0_in,
      CPU_data_master_read_data_valid_nios_system_clock_0_in => CPU_data_master_read_data_valid_nios_system_clock_0_in,
      CPU_data_master_requests_nios_system_clock_0_in => CPU_data_master_requests_nios_system_clock_0_in,
      d1_nios_system_clock_0_in_end_xfer => d1_nios_system_clock_0_in_end_xfer,
      nios_system_clock_0_in_address => nios_system_clock_0_in_address,
      nios_system_clock_0_in_endofpacket_from_sa => nios_system_clock_0_in_endofpacket_from_sa,
      nios_system_clock_0_in_nativeaddress => nios_system_clock_0_in_nativeaddress,
      nios_system_clock_0_in_read => nios_system_clock_0_in_read,
      nios_system_clock_0_in_readdata_from_sa => nios_system_clock_0_in_readdata_from_sa,
      nios_system_clock_0_in_reset_n => nios_system_clock_0_in_reset_n,
      nios_system_clock_0_in_waitrequest_from_sa => nios_system_clock_0_in_waitrequest_from_sa,
      nios_system_clock_0_in_write => nios_system_clock_0_in_write,
      nios_system_clock_0_in_writedata => nios_system_clock_0_in_writedata,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_byteenable => CPU_data_master_byteenable,
      CPU_data_master_dbs_address => CPU_data_master_dbs_address,
      CPU_data_master_dbs_write_8 => CPU_data_master_dbs_write_8,
      CPU_data_master_no_byte_enables_and_last_term => CPU_data_master_no_byte_enables_and_last_term,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_waitrequest => CPU_data_master_waitrequest,
      CPU_data_master_write => CPU_data_master_write,
      clk => internal_sys_clk,
      nios_system_clock_0_in_endofpacket => nios_system_clock_0_in_endofpacket,
      nios_system_clock_0_in_readdata => nios_system_clock_0_in_readdata,
      nios_system_clock_0_in_waitrequest => nios_system_clock_0_in_waitrequest,
      reset_n => sys_clk_reset_n
    );


  --the_nios_system_clock_0_out, which is an e_instance
  the_nios_system_clock_0_out : nios_system_clock_0_out_arbitrator
    port map(
      nios_system_clock_0_out_address_to_slave => nios_system_clock_0_out_address_to_slave,
      nios_system_clock_0_out_readdata => nios_system_clock_0_out_readdata,
      nios_system_clock_0_out_reset_n => nios_system_clock_0_out_reset_n,
      nios_system_clock_0_out_waitrequest => nios_system_clock_0_out_waitrequest,
      External_Clocks_avalon_clocks_slave_readdata_from_sa => External_Clocks_avalon_clocks_slave_readdata_from_sa,
      clk => clk,
      d1_External_Clocks_avalon_clocks_slave_end_xfer => d1_External_Clocks_avalon_clocks_slave_end_xfer,
      nios_system_clock_0_out_address => nios_system_clock_0_out_address,
      nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_granted_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_qualified_request_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_read => nios_system_clock_0_out_read,
      nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_read_data_valid_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave => nios_system_clock_0_out_requests_External_Clocks_avalon_clocks_slave,
      nios_system_clock_0_out_write => nios_system_clock_0_out_write,
      nios_system_clock_0_out_writedata => nios_system_clock_0_out_writedata,
      reset_n => clk_reset_n
    );


  --the_nios_system_clock_0, which is an e_ptf_instance
  the_nios_system_clock_0 : nios_system_clock_0
    port map(
      master_address => nios_system_clock_0_out_address,
      master_nativeaddress => nios_system_clock_0_out_nativeaddress,
      master_read => nios_system_clock_0_out_read,
      master_write => nios_system_clock_0_out_write,
      master_writedata => nios_system_clock_0_out_writedata,
      slave_endofpacket => nios_system_clock_0_in_endofpacket,
      slave_readdata => nios_system_clock_0_in_readdata,
      slave_waitrequest => nios_system_clock_0_in_waitrequest,
      master_clk => clk,
      master_endofpacket => nios_system_clock_0_out_endofpacket,
      master_readdata => nios_system_clock_0_out_readdata,
      master_reset_n => nios_system_clock_0_out_reset_n,
      master_waitrequest => nios_system_clock_0_out_waitrequest,
      slave_address => nios_system_clock_0_in_address,
      slave_clk => internal_sys_clk,
      slave_nativeaddress => nios_system_clock_0_in_nativeaddress,
      slave_read => nios_system_clock_0_in_read,
      slave_reset_n => nios_system_clock_0_in_reset_n,
      slave_write => nios_system_clock_0_in_write,
      slave_writedata => nios_system_clock_0_in_writedata
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      CPU_data_master_granted_sysid_control_slave => CPU_data_master_granted_sysid_control_slave,
      CPU_data_master_qualified_request_sysid_control_slave => CPU_data_master_qualified_request_sysid_control_slave,
      CPU_data_master_read_data_valid_sysid_control_slave => CPU_data_master_read_data_valid_sysid_control_slave,
      CPU_data_master_requests_sysid_control_slave => CPU_data_master_requests_sysid_control_slave,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      CPU_data_master_address_to_slave => CPU_data_master_address_to_slave,
      CPU_data_master_read => CPU_data_master_read,
      CPU_data_master_write => CPU_data_master_write,
      clk => internal_sys_clk,
      reset_n => sys_clk_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address
    );


  --reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_sys_clk_domain_synch : nios_system_reset_sys_clk_domain_synch_module
    port map(
      data_out => sys_clk_reset_n,
      clk => internal_sys_clk,
      data_in => module_input12,
      reset_n => reset_n_sources
    );

  module_input12 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(CPU_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000"))));
  --reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_clk_domain_synch : nios_system_reset_clk_domain_synch_module
    port map(
      data_out => clk_reset_n,
      clk => clk,
      data_in => module_input13,
      reset_n => reset_n_sources
    );

  module_input13 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_vga_clk_domain_synch : nios_system_reset_vga_clk_domain_synch_module
    port map(
      data_out => vga_clk_reset_n,
      clk => internal_vga_clk,
      data_in => module_input14,
      reset_n => reset_n_sources
    );

  module_input14 <= std_logic'('1');

  --nios_system_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios_system_clock_0_out_endofpacket <= std_logic'('0');
  --vhdl renameroo for output signals
  AUD_DACDAT_from_the_Audio <= internal_AUD_DACDAT_from_the_Audio;
  --vhdl renameroo for output signals
  HEX0_from_the_HEX3_HEX0 <= internal_HEX0_from_the_HEX3_HEX0;
  --vhdl renameroo for output signals
  HEX1_from_the_HEX3_HEX0 <= internal_HEX1_from_the_HEX3_HEX0;
  --vhdl renameroo for output signals
  HEX2_from_the_HEX3_HEX0 <= internal_HEX2_from_the_HEX3_HEX0;
  --vhdl renameroo for output signals
  HEX3_from_the_HEX3_HEX0 <= internal_HEX3_from_the_HEX3_HEX0;
  --vhdl renameroo for output signals
  HEX4_from_the_HEX7_HEX4 <= internal_HEX4_from_the_HEX7_HEX4;
  --vhdl renameroo for output signals
  HEX5_from_the_HEX7_HEX4 <= internal_HEX5_from_the_HEX7_HEX4;
  --vhdl renameroo for output signals
  HEX6_from_the_HEX7_HEX4 <= internal_HEX6_from_the_HEX7_HEX4;
  --vhdl renameroo for output signals
  HEX7_from_the_HEX7_HEX4 <= internal_HEX7_from_the_HEX7_HEX4;
  --vhdl renameroo for output signals
  I2C_SCLK_from_the_AV_Config <= internal_I2C_SCLK_from_the_AV_Config;
  --vhdl renameroo for output signals
  LCD_BLON_from_the_Char_LCD_16x2 <= internal_LCD_BLON_from_the_Char_LCD_16x2;
  --vhdl renameroo for output signals
  LCD_EN_from_the_Char_LCD_16x2 <= internal_LCD_EN_from_the_Char_LCD_16x2;
  --vhdl renameroo for output signals
  LCD_ON_from_the_Char_LCD_16x2 <= internal_LCD_ON_from_the_Char_LCD_16x2;
  --vhdl renameroo for output signals
  LCD_RS_from_the_Char_LCD_16x2 <= internal_LCD_RS_from_the_Char_LCD_16x2;
  --vhdl renameroo for output signals
  LCD_RW_from_the_Char_LCD_16x2 <= internal_LCD_RW_from_the_Char_LCD_16x2;
  --vhdl renameroo for output signals
  LEDG_from_the_Green_LEDs <= internal_LEDG_from_the_Green_LEDs;
  --vhdl renameroo for output signals
  LEDR_from_the_Red_LEDs <= internal_LEDR_from_the_Red_LEDs;
  --vhdl renameroo for output signals
  SRAM_ADDR_from_the_SRAM <= internal_SRAM_ADDR_from_the_SRAM;
  --vhdl renameroo for output signals
  SRAM_CE_N_from_the_SRAM <= internal_SRAM_CE_N_from_the_SRAM;
  --vhdl renameroo for output signals
  SRAM_LB_N_from_the_SRAM <= internal_SRAM_LB_N_from_the_SRAM;
  --vhdl renameroo for output signals
  SRAM_OE_N_from_the_SRAM <= internal_SRAM_OE_N_from_the_SRAM;
  --vhdl renameroo for output signals
  SRAM_UB_N_from_the_SRAM <= internal_SRAM_UB_N_from_the_SRAM;
  --vhdl renameroo for output signals
  SRAM_WE_N_from_the_SRAM <= internal_SRAM_WE_N_from_the_SRAM;
  --vhdl renameroo for output signals
  UART_TXD_from_the_Serial_Port <= internal_UART_TXD_from_the_Serial_Port;
  --vhdl renameroo for output signals
  VGA_BLANK_from_the_VGA_Controller <= internal_VGA_BLANK_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_B_from_the_VGA_Controller <= internal_VGA_B_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_CLK_from_the_VGA_Controller <= internal_VGA_CLK_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_G_from_the_VGA_Controller <= internal_VGA_G_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_HS_from_the_VGA_Controller <= internal_VGA_HS_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_R_from_the_VGA_Controller <= internal_VGA_R_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_SYNC_from_the_VGA_Controller <= internal_VGA_SYNC_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  VGA_VS_from_the_VGA_Controller <= internal_VGA_VS_from_the_VGA_Controller;
  --vhdl renameroo for output signals
  sys_clk <= internal_sys_clk;
  --vhdl renameroo for output signals
  vga_clk <= internal_vga_clk;
  --vhdl renameroo for output signals
  zs_addr_from_the_SDRAM <= internal_zs_addr_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_ba_from_the_SDRAM <= internal_zs_ba_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_SDRAM <= internal_zs_cas_n_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_cke_from_the_SDRAM <= internal_zs_cke_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_SDRAM <= internal_zs_cs_n_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_dqm_from_the_SDRAM <= internal_zs_dqm_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_SDRAM <= internal_zs_ras_n_from_the_SDRAM;
  --vhdl renameroo for output signals
  zs_we_n_from_the_SDRAM <= internal_zs_we_n_from_the_SDRAM;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component nios_system is 
           port (
                 -- 1) global signals:
                    signal audio_clk : OUT STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clk_27 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_clk : OUT STD_LOGIC;
                    signal sys_clk : OUT STD_LOGIC;
                    signal vga_clk : OUT STD_LOGIC;

                 -- the_AV_Config
                    signal I2C_SCLK_from_the_AV_Config : OUT STD_LOGIC;
                    signal I2C_SDAT_to_and_from_the_AV_Config : INOUT STD_LOGIC;

                 -- the_Audio
                    signal AUD_ADCDAT_to_the_Audio : IN STD_LOGIC;
                    signal AUD_ADCLRCK_to_and_from_the_Audio : INOUT STD_LOGIC;
                    signal AUD_BCLK_to_and_from_the_Audio : INOUT STD_LOGIC;
                    signal AUD_DACDAT_from_the_Audio : OUT STD_LOGIC;
                    signal AUD_DACLRCK_to_and_from_the_Audio : INOUT STD_LOGIC;

                 -- the_Char_LCD_16x2
                    signal LCD_BLON_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                    signal LCD_DATA_to_and_from_the_Char_LCD_16x2 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal LCD_EN_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                    signal LCD_ON_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                    signal LCD_RS_from_the_Char_LCD_16x2 : OUT STD_LOGIC;
                    signal LCD_RW_from_the_Char_LCD_16x2 : OUT STD_LOGIC;

                 -- the_Expansion_JP1
                    signal GPIO_0_to_and_from_the_Expansion_JP1 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- the_Expansion_JP2
                    signal GPIO_1_to_and_from_the_Expansion_JP2 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- the_Green_LEDs
                    signal LEDG_from_the_Green_LEDs : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);

                 -- the_HEX3_HEX0
                    signal HEX0_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX1_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX2_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX3_from_the_HEX3_HEX0 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);

                 -- the_HEX7_HEX4
                    signal HEX4_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX5_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX6_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal HEX7_from_the_HEX7_HEX4 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);

                 -- the_PS2_Port
                    signal PS2_CLK_to_and_from_the_PS2_Port : INOUT STD_LOGIC;
                    signal PS2_DAT_to_and_from_the_PS2_Port : INOUT STD_LOGIC;

                 -- the_Pushbuttons
                    signal KEY_to_the_Pushbuttons : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_Red_LEDs
                    signal LEDR_from_the_Red_LEDs : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);

                 -- the_SDRAM
                    signal zs_addr_from_the_SDRAM : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba_from_the_SDRAM : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_SDRAM : OUT STD_LOGIC;
                    signal zs_cke_from_the_SDRAM : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_SDRAM : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_SDRAM : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm_from_the_SDRAM : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n_from_the_SDRAM : OUT STD_LOGIC;
                    signal zs_we_n_from_the_SDRAM : OUT STD_LOGIC;

                 -- the_SRAM
                    signal SRAM_ADDR_from_the_SRAM : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal SRAM_CE_N_from_the_SRAM : OUT STD_LOGIC;
                    signal SRAM_DQ_to_and_from_the_SRAM : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_LB_N_from_the_SRAM : OUT STD_LOGIC;
                    signal SRAM_OE_N_from_the_SRAM : OUT STD_LOGIC;
                    signal SRAM_UB_N_from_the_SRAM : OUT STD_LOGIC;
                    signal SRAM_WE_N_from_the_SRAM : OUT STD_LOGIC;

                 -- the_Serial_Port
                    signal UART_RXD_to_the_Serial_Port : IN STD_LOGIC;
                    signal UART_TXD_from_the_Serial_Port : OUT STD_LOGIC;

                 -- the_Slider_Switches
                    signal SW_to_the_Slider_Switches : IN STD_LOGIC_VECTOR (17 DOWNTO 0);

                 -- the_VGA_Controller
                    signal VGA_BLANK_from_the_VGA_Controller : OUT STD_LOGIC;
                    signal VGA_B_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_CLK_from_the_VGA_Controller : OUT STD_LOGIC;
                    signal VGA_G_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_HS_from_the_VGA_Controller : OUT STD_LOGIC;
                    signal VGA_R_from_the_VGA_Controller : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_SYNC_from_the_VGA_Controller : OUT STD_LOGIC;
                    signal VGA_VS_from_the_VGA_Controller : OUT STD_LOGIC
                 );
end component nios_system;

                signal AUD_ADCDAT_to_the_Audio :  STD_LOGIC;
                signal AUD_ADCLRCK_to_and_from_the_Audio :  STD_LOGIC;
                signal AUD_BCLK_to_and_from_the_Audio :  STD_LOGIC;
                signal AUD_DACDAT_from_the_Audio :  STD_LOGIC;
                signal AUD_DACLRCK_to_and_from_the_Audio :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal CPU_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_status :  STD_LOGIC;
                signal CPU_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal GPIO_0_to_and_from_the_Expansion_JP1 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal GPIO_1_to_and_from_the_Expansion_JP2 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal HEX0_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX1_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX2_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX3_from_the_HEX3_HEX0 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX4_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX5_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX6_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal HEX7_from_the_HEX7_HEX4 :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal I2C_SCLK_from_the_AV_Config :  STD_LOGIC;
                signal I2C_SDAT_to_and_from_the_AV_Config :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal JTAG_UART_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal KEY_to_the_Pushbuttons :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal LCD_BLON_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal LCD_DATA_to_and_from_the_Char_LCD_16x2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal LCD_EN_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal LCD_ON_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal LCD_RS_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal LCD_RW_from_the_Char_LCD_16x2 :  STD_LOGIC;
                signal LEDG_from_the_Green_LEDs :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal LEDR_from_the_Red_LEDs :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal PS2_CLK_to_and_from_the_PS2_Port :  STD_LOGIC;
                signal PS2_DAT_to_and_from_the_PS2_Port :  STD_LOGIC;
                signal SRAM_ADDR_from_the_SRAM :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal SRAM_CE_N_from_the_SRAM :  STD_LOGIC;
                signal SRAM_DQ_to_and_from_the_SRAM :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SRAM_LB_N_from_the_SRAM :  STD_LOGIC;
                signal SRAM_OE_N_from_the_SRAM :  STD_LOGIC;
                signal SRAM_UB_N_from_the_SRAM :  STD_LOGIC;
                signal SRAM_WE_N_from_the_SRAM :  STD_LOGIC;
                signal SW_to_the_Slider_Switches :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal UART_RXD_to_the_Serial_Port :  STD_LOGIC;
                signal UART_TXD_from_the_Serial_Port :  STD_LOGIC;
                signal VGA_BLANK_from_the_VGA_Controller :  STD_LOGIC;
                signal VGA_B_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_CLK_from_the_VGA_Controller :  STD_LOGIC;
                signal VGA_G_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_HS_from_the_VGA_Controller :  STD_LOGIC;
                signal VGA_R_from_the_VGA_Controller :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_SYNC_from_the_VGA_Controller :  STD_LOGIC;
                signal VGA_VS_from_the_VGA_Controller :  STD_LOGIC;
                signal audio_clk :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_27 :  STD_LOGIC;
                signal nios_system_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios_system_clock_0_out_endofpacket :  STD_LOGIC;
                signal nios_system_clock_0_out_nativeaddress :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal sdram_clk :  STD_LOGIC;
                signal sys_clk :  STD_LOGIC;
                signal vga_clk :  STD_LOGIC;
                signal zs_addr_from_the_SDRAM :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal zs_ba_from_the_SDRAM :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_SDRAM :  STD_LOGIC;
                signal zs_cke_from_the_SDRAM :  STD_LOGIC;
                signal zs_cs_n_from_the_SDRAM :  STD_LOGIC;
                signal zs_dq_to_and_from_the_SDRAM :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal zs_dqm_from_the_SDRAM :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_ras_n_from_the_SDRAM :  STD_LOGIC;
                signal zs_we_n_from_the_SDRAM :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : nios_system
    port map(
      AUD_ADCLRCK_to_and_from_the_Audio => AUD_ADCLRCK_to_and_from_the_Audio,
      AUD_BCLK_to_and_from_the_Audio => AUD_BCLK_to_and_from_the_Audio,
      AUD_DACDAT_from_the_Audio => AUD_DACDAT_from_the_Audio,
      AUD_DACLRCK_to_and_from_the_Audio => AUD_DACLRCK_to_and_from_the_Audio,
      GPIO_0_to_and_from_the_Expansion_JP1 => GPIO_0_to_and_from_the_Expansion_JP1,
      GPIO_1_to_and_from_the_Expansion_JP2 => GPIO_1_to_and_from_the_Expansion_JP2,
      HEX0_from_the_HEX3_HEX0 => HEX0_from_the_HEX3_HEX0,
      HEX1_from_the_HEX3_HEX0 => HEX1_from_the_HEX3_HEX0,
      HEX2_from_the_HEX3_HEX0 => HEX2_from_the_HEX3_HEX0,
      HEX3_from_the_HEX3_HEX0 => HEX3_from_the_HEX3_HEX0,
      HEX4_from_the_HEX7_HEX4 => HEX4_from_the_HEX7_HEX4,
      HEX5_from_the_HEX7_HEX4 => HEX5_from_the_HEX7_HEX4,
      HEX6_from_the_HEX7_HEX4 => HEX6_from_the_HEX7_HEX4,
      HEX7_from_the_HEX7_HEX4 => HEX7_from_the_HEX7_HEX4,
      I2C_SCLK_from_the_AV_Config => I2C_SCLK_from_the_AV_Config,
      I2C_SDAT_to_and_from_the_AV_Config => I2C_SDAT_to_and_from_the_AV_Config,
      LCD_BLON_from_the_Char_LCD_16x2 => LCD_BLON_from_the_Char_LCD_16x2,
      LCD_DATA_to_and_from_the_Char_LCD_16x2 => LCD_DATA_to_and_from_the_Char_LCD_16x2,
      LCD_EN_from_the_Char_LCD_16x2 => LCD_EN_from_the_Char_LCD_16x2,
      LCD_ON_from_the_Char_LCD_16x2 => LCD_ON_from_the_Char_LCD_16x2,
      LCD_RS_from_the_Char_LCD_16x2 => LCD_RS_from_the_Char_LCD_16x2,
      LCD_RW_from_the_Char_LCD_16x2 => LCD_RW_from_the_Char_LCD_16x2,
      LEDG_from_the_Green_LEDs => LEDG_from_the_Green_LEDs,
      LEDR_from_the_Red_LEDs => LEDR_from_the_Red_LEDs,
      PS2_CLK_to_and_from_the_PS2_Port => PS2_CLK_to_and_from_the_PS2_Port,
      PS2_DAT_to_and_from_the_PS2_Port => PS2_DAT_to_and_from_the_PS2_Port,
      SRAM_ADDR_from_the_SRAM => SRAM_ADDR_from_the_SRAM,
      SRAM_CE_N_from_the_SRAM => SRAM_CE_N_from_the_SRAM,
      SRAM_DQ_to_and_from_the_SRAM => SRAM_DQ_to_and_from_the_SRAM,
      SRAM_LB_N_from_the_SRAM => SRAM_LB_N_from_the_SRAM,
      SRAM_OE_N_from_the_SRAM => SRAM_OE_N_from_the_SRAM,
      SRAM_UB_N_from_the_SRAM => SRAM_UB_N_from_the_SRAM,
      SRAM_WE_N_from_the_SRAM => SRAM_WE_N_from_the_SRAM,
      UART_TXD_from_the_Serial_Port => UART_TXD_from_the_Serial_Port,
      VGA_BLANK_from_the_VGA_Controller => VGA_BLANK_from_the_VGA_Controller,
      VGA_B_from_the_VGA_Controller => VGA_B_from_the_VGA_Controller,
      VGA_CLK_from_the_VGA_Controller => VGA_CLK_from_the_VGA_Controller,
      VGA_G_from_the_VGA_Controller => VGA_G_from_the_VGA_Controller,
      VGA_HS_from_the_VGA_Controller => VGA_HS_from_the_VGA_Controller,
      VGA_R_from_the_VGA_Controller => VGA_R_from_the_VGA_Controller,
      VGA_SYNC_from_the_VGA_Controller => VGA_SYNC_from_the_VGA_Controller,
      VGA_VS_from_the_VGA_Controller => VGA_VS_from_the_VGA_Controller,
      audio_clk => audio_clk,
      sdram_clk => sdram_clk,
      sys_clk => sys_clk,
      vga_clk => vga_clk,
      zs_addr_from_the_SDRAM => zs_addr_from_the_SDRAM,
      zs_ba_from_the_SDRAM => zs_ba_from_the_SDRAM,
      zs_cas_n_from_the_SDRAM => zs_cas_n_from_the_SDRAM,
      zs_cke_from_the_SDRAM => zs_cke_from_the_SDRAM,
      zs_cs_n_from_the_SDRAM => zs_cs_n_from_the_SDRAM,
      zs_dq_to_and_from_the_SDRAM => zs_dq_to_and_from_the_SDRAM,
      zs_dqm_from_the_SDRAM => zs_dqm_from_the_SDRAM,
      zs_ras_n_from_the_SDRAM => zs_ras_n_from_the_SDRAM,
      zs_we_n_from_the_SDRAM => zs_we_n_from_the_SDRAM,
      AUD_ADCDAT_to_the_Audio => AUD_ADCDAT_to_the_Audio,
      KEY_to_the_Pushbuttons => KEY_to_the_Pushbuttons,
      SW_to_the_Slider_Switches => SW_to_the_Slider_Switches,
      UART_RXD_to_the_Serial_Port => UART_RXD_to_the_Serial_Port,
      clk => clk,
      clk_27 => clk_27,
      reset_n => reset_n
    );


  process
  begin
    clk <= '0';
    loop
       wait for 10 ns;
       clk <= not clk;
    end loop;
  end process;
  process
  begin
    clk_27 <= '0';
    loop
       if (clk_27 = '1') then
          wait for 18 ns;
          clk_27 <= not clk_27;
       else
          wait for 19 ns;
          clk_27 <= not clk_27;
       end if;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
