library ieee;
USE IEEE.NUMERIC_STD.ALL; USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL; USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--------------------------------------------------------------
ENTITY lab5 IS
port (clk1 : in std_logic;
      seconds : out std_logic_vector(5 downto 0);
      minutes : out std_logic_vector(5 downto 0);
      hours : out std_logic_vector(4 downto 0)
		);
end lab5;
-------------------------------------------------------------
architecture behavior of lab5 is
	signal sec,min,hour : integer range 0 to 60 :=0;
	signal count : integer :=1;
	signal clk : std_logic :='0';
begin
seconds <= conv_std_logic_vector(sec,6);
minutes <= conv_std_logic_vector(min,6);
hours <= conv_std_logic_vector(hour,5);

 --clk generation.For 100 MHz clock this generates 1 Hz clock.
process(clk1)
begin
	if(clk1'event and clk1='1') then
		count <=count+1;
		if(count = 50000000) then
		clk <= not clk;
		count <=1;
		end if;
	end if;
end process;

--period of clk is 1 second. Counter Divider
process(clk)   
begin

if(clk'event and clk='1') then
sec <= sec+ 1;
if(sec = 59) then
sec<=0;
min <= min + 1;
if(min = 59) then
hour <= hour + 1;
min <= 0;
if(hour = 23) then
hour <= 0;
end if;
end if;
end if;
end if;

end process;

end behavior;