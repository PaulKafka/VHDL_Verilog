  --Example instantiation for system 'nios_system'
  nios_system_inst : nios_system
    port map(
      AUD_ADCLRCK_to_and_from_the_Audio => AUD_ADCLRCK_to_and_from_the_Audio,
      AUD_BCLK_to_and_from_the_Audio => AUD_BCLK_to_and_from_the_Audio,
      AUD_DACDAT_from_the_Audio => AUD_DACDAT_from_the_Audio,
      AUD_DACLRCK_to_and_from_the_Audio => AUD_DACLRCK_to_and_from_the_Audio,
      GPIO_0_to_and_from_the_Expansion_JP1 => GPIO_0_to_and_from_the_Expansion_JP1,
      GPIO_1_to_and_from_the_Expansion_JP2 => GPIO_1_to_and_from_the_Expansion_JP2,
      HEX0_from_the_HEX3_HEX0 => HEX0_from_the_HEX3_HEX0,
      HEX1_from_the_HEX3_HEX0 => HEX1_from_the_HEX3_HEX0,
      HEX2_from_the_HEX3_HEX0 => HEX2_from_the_HEX3_HEX0,
      HEX3_from_the_HEX3_HEX0 => HEX3_from_the_HEX3_HEX0,
      HEX4_from_the_HEX7_HEX4 => HEX4_from_the_HEX7_HEX4,
      HEX5_from_the_HEX7_HEX4 => HEX5_from_the_HEX7_HEX4,
      HEX6_from_the_HEX7_HEX4 => HEX6_from_the_HEX7_HEX4,
      HEX7_from_the_HEX7_HEX4 => HEX7_from_the_HEX7_HEX4,
      I2C_SCLK_from_the_AV_Config => I2C_SCLK_from_the_AV_Config,
      I2C_SDAT_to_and_from_the_AV_Config => I2C_SDAT_to_and_from_the_AV_Config,
      LCD_BLON_from_the_Char_LCD_16x2 => LCD_BLON_from_the_Char_LCD_16x2,
      LCD_DATA_to_and_from_the_Char_LCD_16x2 => LCD_DATA_to_and_from_the_Char_LCD_16x2,
      LCD_EN_from_the_Char_LCD_16x2 => LCD_EN_from_the_Char_LCD_16x2,
      LCD_ON_from_the_Char_LCD_16x2 => LCD_ON_from_the_Char_LCD_16x2,
      LCD_RS_from_the_Char_LCD_16x2 => LCD_RS_from_the_Char_LCD_16x2,
      LCD_RW_from_the_Char_LCD_16x2 => LCD_RW_from_the_Char_LCD_16x2,
      LEDG_from_the_Green_LEDs => LEDG_from_the_Green_LEDs,
      LEDR_from_the_Red_LEDs => LEDR_from_the_Red_LEDs,
      PS2_CLK_to_and_from_the_PS2_Port => PS2_CLK_to_and_from_the_PS2_Port,
      PS2_DAT_to_and_from_the_PS2_Port => PS2_DAT_to_and_from_the_PS2_Port,
      SRAM_ADDR_from_the_SRAM => SRAM_ADDR_from_the_SRAM,
      SRAM_CE_N_from_the_SRAM => SRAM_CE_N_from_the_SRAM,
      SRAM_DQ_to_and_from_the_SRAM => SRAM_DQ_to_and_from_the_SRAM,
      SRAM_LB_N_from_the_SRAM => SRAM_LB_N_from_the_SRAM,
      SRAM_OE_N_from_the_SRAM => SRAM_OE_N_from_the_SRAM,
      SRAM_UB_N_from_the_SRAM => SRAM_UB_N_from_the_SRAM,
      SRAM_WE_N_from_the_SRAM => SRAM_WE_N_from_the_SRAM,
      UART_TXD_from_the_Serial_Port => UART_TXD_from_the_Serial_Port,
      VGA_BLANK_from_the_VGA_Controller => VGA_BLANK_from_the_VGA_Controller,
      VGA_B_from_the_VGA_Controller => VGA_B_from_the_VGA_Controller,
      VGA_CLK_from_the_VGA_Controller => VGA_CLK_from_the_VGA_Controller,
      VGA_G_from_the_VGA_Controller => VGA_G_from_the_VGA_Controller,
      VGA_HS_from_the_VGA_Controller => VGA_HS_from_the_VGA_Controller,
      VGA_R_from_the_VGA_Controller => VGA_R_from_the_VGA_Controller,
      VGA_SYNC_from_the_VGA_Controller => VGA_SYNC_from_the_VGA_Controller,
      VGA_VS_from_the_VGA_Controller => VGA_VS_from_the_VGA_Controller,
      audio_clk => audio_clk,
      sdram_clk => sdram_clk,
      sys_clk => sys_clk,
      vga_clk => vga_clk,
      zs_addr_from_the_SDRAM => zs_addr_from_the_SDRAM,
      zs_ba_from_the_SDRAM => zs_ba_from_the_SDRAM,
      zs_cas_n_from_the_SDRAM => zs_cas_n_from_the_SDRAM,
      zs_cke_from_the_SDRAM => zs_cke_from_the_SDRAM,
      zs_cs_n_from_the_SDRAM => zs_cs_n_from_the_SDRAM,
      zs_dq_to_and_from_the_SDRAM => zs_dq_to_and_from_the_SDRAM,
      zs_dqm_from_the_SDRAM => zs_dqm_from_the_SDRAM,
      zs_ras_n_from_the_SDRAM => zs_ras_n_from_the_SDRAM,
      zs_we_n_from_the_SDRAM => zs_we_n_from_the_SDRAM,
      AUD_ADCDAT_to_the_Audio => AUD_ADCDAT_to_the_Audio,
      KEY_to_the_Pushbuttons => KEY_to_the_Pushbuttons,
      SW_to_the_Slider_Switches => SW_to_the_Slider_Switches,
      UART_RXD_to_the_Serial_Port => UART_RXD_to_the_Serial_Port,
      clk => clk,
      clk_27 => clk_27,
      reset_n => reset_n
    );


