��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ��>�(Ŗ�6�eQ�d*e��!i�v�4G[�\)C��S� y3�Xv��XcϷ�z���B�}��uE�Oz��q��̷s��n~܌W2����C�x��.ם:��˂S	�J�����ڐ�
�^ �	s�'�%���gM7�� �7���8�߻�So����@��>#�wiE�]�Da\E�ʙψ"�՘~z�X��)�f��D�y&�-��8R}qI���=-@Z.�������&�B�p4Z��q��M��c���j�R���AFW��\�T�Ɏbof�#<Y�^��c�=�|Xi�/7��� �#F�	Z�om�&��0�{��Ph۟p��_��s�-�|3�b����߻Ș�2���U�L�g�'Ň�&����!q�4bs!�V�#6��F���BGo�f�y�IU�o-(ޡ���W@�B��,��T%�*�a�i���jӄm�������H�C����ޟ���u2�g��'�Tf 4x��7�c
�^�N� �rR��/�7����n�U����'��b(�|��*U`�%�U�m�EQ����n���8���!*�O���0��3:�q��D:	�]a��N��^�Sk�9o᥅�l�SP��&������<��a~��+���CO߿EI��M�	*���tQ��SP��s:�[hl��_q�1��Qcp�?u�W!L��ႲW�Nïy&`�;KrS�6��5m���I#���^$o��0]�mE�FH.I]p���K3҇4���R\�7�^��	���
�E��7�w�,�$˱����eΨ���ow!9�����y8@�l��۷��7�:#.�A
�/G�e��+g"���BT�w�W���s�x�jgW'욦����/��@g�}�F2��w(Kzg�؃ba���*���������u����h�`]8x�#2jx�I�Ɨ�
�����: ����t���4NU?�S\�>g�q���3�=���Y��%X��D�F_�{�u����u���� ��v^���p���5Bp³�"�
u������W�N�����.�;`��+�ߴ�-;,2��jRQ���� Ȳ-I	&9��w�������W$���%^�mwEA��&=�˷���WEx�2��#`PJ��U߷7��gA(�)�D��X��M�9Ap9x-\�͇Y�&cbc�X+V�'+3���S+)�';���f�k�T����ir-�IA����ϑ�%�3.�{�SI@*>ϖS��!ԯ�k��=-���,�^Z_6�B�z+,-=�� ]!�L����g��!���<��~v�=cz;Z�Ո7��-5�;f툃� ��w�~,]p� Qn!�����F����=�C�yɀ�e_B�����2#�:�%��xMi� �sT�=�Z��CWy�cv.����xF��5�$�K�˘6ᖷp-W��T�8�����n����U����[���e74Q��:�:va����y����~9k虯�h�
�Cܳ%/dR�-�ͼ�����Ş����� �)���&W�*�u��#��[�i����7���C���&�X�lT�����Fх)�z�a���\��S�R�6���}]��m#��B��l��Ҿ.����o�FrZ9�٨�K��n^��Z�EFGx,ht�+65�&�b*ǂI�׆��"�X��O)��M�#VV��C?6��T��� .Ԍ�R����_C�e˲C1w͖#��g�u��n��x̖�{�[��t]�s�q�D^��h�soȃ`�V�췴��^P�����I5c9c�Gg�B3��4�q���ĩ
���;h�:�%\��琮�����E�v�����{���q~��,l���<��K��P���WL<��+~�e>N)R&ɷ%.Yˬf�`?L��IC@�֜�L�zM�Gu�4w�ҥn�?5_{�hG\��\d��qB�Ac_�>���zFAW�GpGL�a��L�Ÿl���y1�q$c �k�����}��
yo��e��=A���4�*G�r*w��m:�6<�X�T�I�s��L�#��-׎D�~4��2�Ye_ܸD��J�Z�3�"�L�(�%kr26��
�]W53L&Ѡ���6/�\=��/��7-�$�t+�}��M"��{��D���F�r���̱R�S��e� 8|'��CM������q��c:TKq�Dx�IV	(��
V\9����26��+��ب�db�U>T��ĮQxڒ��Z{<�㒩�o؝�N'�/�$\���7�F�w�R��3c�nw�,4%�A�Y;# y����H��j���T,�ЩW-~�G���s���ɑ��*�]�6w# ��>t�Ў�Sؐ�*�#���y�G�	~�ߌ8���b�@�ƥ�j�I��&��Gb��l�]���ZA\��|i�p:J�R��\��>��ˉ�y�Ϣ�P�<Z^I⢸e�tM�1���J��K����"}*���]��������f�d"��Z��1��r�E�aۄ��Y��T� ��g4K�Q�=D�&�\�uV�.�qɪ�xJ�#w��f0/g۞d1�i'-Qb��~���8r�H*��W�V��;*��Mt��_�@�H�e�F� ix�s4��ύj�۞��1��FU��C�,(q��+�	��J�UFtڞ�Ih	��ݻ7S-�-��Uv,�I4f!N�pc0+�@��X�K�n�S�lf >l�Y���̀ǈ3��eazʥ�c�˾��ɮ� �L�&f,���53D�'�����ׯ�N��8ߊj3J[23ɲ!�]F#�f�x��`ȥ���B��jg$8���F��b���N���c@��n�o��c6Maq[)��ݗ�,T��z��͋�<��Y����=ť��ɹzbw��I�3���x��}�D�Dz�w͊w�-���˼��mG��#����A6�i���`���1��)6��c迪�s���9k��1I�H�G�i(����oh\/b<5s�4��/e�pŷFQ� ꁱ+�ȖA��CƁ5̶���}�V���k�|�艛��eH�4NXl	$SL��9c�8�侶��4��w⟰�WUW��ol�9eS��H�"Q��g�1j(�U�$?�oW \�MO6�:o��|�=x'㜑�X�C�{rU"����B��iJ�|�*�cŝ�(�31ٶu��E �X4q�*�Ymٵ�a�(d}l̺����u�#"ny�"
W a��>ͦ_�./�nUhO6ʙ��[k����q�x��z�Ώ�,��(B��0r���k.��-�.��ΪI�"Ֆ�\Mjpy�˹\�\�ޭT�Ք� 3�NE�]��y�
�+e��ue�P����L�rkR��_��%�A���Vr7y��{�XWd���1����a��X���F���O�9�?4�+�֐b��C�eȈ��'���g��3#'K�u�Ic�����L.먖	�6��0[�J��bzb��q�1�T2�&�~tI�s�:���P���F����!���y�;����O�)��vvse��u:�g��T�V��TX���dza��2o��h
����5ʅՇI�b���&������P�38`E`V�_-,l�M��٫��n4Th���d���*�����S�'�%zeO��'��J���Z߶3�ZHi�+6�G�j')�%{�{b�7[�]ёdo�v���!�1}�S'^���L���"փ�5�TIhb}&���7���'N�Z��?�	���+�8�QE3�rz��-$��Bl���/q;d�V�$�d�?� Vtw�j���<6VT	��H��iQ�60Qlj,�FV�Xxrnc��#)1I�0?"�����1�@d��A>�֧ ?��o�'�8hr�q�l�8ո���2����}!h�S����xT���=M��������q�%���a3q�bA���#g��}n�
ዷ�p��w2l�o8�}8iZ� 5���<x�5��:*A���ξ(�bi��Ӛ�� ��e=�E���G�qh���2�=�1*ǥ�Q�ռ	ΖV�e��;{�ĸ�P
g��q�[����J�-x>xs���ۘ�:$�}���'0��/cL��H�xO\y�ý�K6,�9�����@�%�U��h���;���U���t��n��>I�£�����1ϵ�GH��7�v�k�©o��,R"�M���v�Z��\�� �u���#��h^�p�6R<j�	s�}�W��CA~/4�.���M��1k.|x#����j��6��>��.�>|-�=رN?|;����K�;��H�BC��U����怒�H�H�3.J6oػ���3y�j=����VIIF�@ѕ��oܐs�!��]Yґ��9����s�9;��jc�.���|\��
,u���Y��:I�s9��*ykf�oG�HoO_H��å+�A4���6	*�[5!o����4:6����(<�5ڨ���Ao��T��cs�HE�I-a�	a���^H��a<ot��������t0�V�P�{>�w�5�[���<>1r3M�{g[��
	�2�/΀�!�Dr�f��M4Q`}]���u���M�>Tw˭��s���$�<����V*�OGd8.���`[]y+K.��|i^�oT�mɝRD^�ci�$D�2E�B]�����l�	�
�we�O�AS.sIb�@Q���9��#����z�qR�9_T$�OaVT�^&Q�w�@݆��՟�?�)b���g^ ��	ԗx��8-�K8��`(	j�*��J�P�)��D�j�֒I����𥮵 �cqD�W��k��x�#G�4A�o�ym=UT[���E�'�Ƈ�$�7���f��Z2�P�'�v䘺5�/	��^�=~���8J�p���.#�� ��B������T��pF�u������cG���uZ
Ls1�/%�`����(����Dl����Y��r�nY������� �k���N�@K��Y\/�q
�8�M�~������!-��7��|�cDW�x�@��(�*���y��1�U�FY�(剛�����ٕ�z3�@-��ho�>h�R)�L��s���R(���KS�A����t�J8:��,u\��x����T��N��N�\��UU���]H��u�1"�F1��J���?M��!pd��F�D#�R�5ˡ2;�jA����B��j������{?`-ּ�a-qN�lF���c�m�-m���{�՗e�K´��3����
��xF���Y~h��䳽xQ��ѳ���l�9"xc�񰎋m&��O����Fk��?�U};^ׇ����(���؉
�������2�Q��Wu�g���}2���B�+'�r(3�UG#Ğ�Ǻ���
ckC��g		���^�hk4�/l�"_�oI��ҋ�b���굣��^�4�6�D]O����x8������ϐ�F�>�4)�C_��S�����K�3z�P�����r��a���?�؀:�ʨ	 |n���#y��3�N�z"�����:���l�]����:G���Ą*hDc�隸4�̍�c�B��%���}-���/�|���/Mxi���XI���=.f�@���
1Z�ҙ�FA�ƪ�r4m<#�_9�S�o�eF@0�~����p����޽uﳫ����u��aD+L�@�9&My���V(~���h���7+�t�ާ��s.�8�+c1��E��� Qg����W >3��%�*��0 ����0���}�o/
�1��d��B�ޚ#���څ���S}"U�@�U������ U���`�y�����!Z���_���5em��,������u�%��Vԫq�ɩ��Y."V
JC}C��͂�a
-H�RҔn�e%`=up0���� ��ܫ��RQ�9w\����� |�;���L�_ZW�qX�ehw%E�L�04�Ř-��rF��� ��ڭ"���ߥ&J=7��`�;e�8H�&H<�\�	���9�$���+�9�_^���V��0aw�K���mk��z�����s��?�Q��MI�71����@q[�ph³��s��ZU;O��_�B�!h�r���π~�l6�T �� ��x����Z�IT�C'�_0�c���$9�\T4E�?�6�j9�r�s��H�K=/p-U��*�*��o ���.��N��c}�
�� ��X�k�K����Z����5y��:�옴3j�Fi7��[0M8���'`����I/H �������LI"����RI��ȓ#�0;k{�n� ���|�R��~�M�q0PcW@��k�6��$��Uې����;�vr�r�+��bl�i�5����&�����!�{K��V4���:}���+��0S��^kW$vإ�]��	��C���ؒ-wg�w�L��J���wFR�XUA1h��{R���{x�_�˵m��L��db� պ�,Δ�d��z?E9S�ø*�3)�s�/7��	��{��Y��U��f�Yw��aD"�<��p0O�WT���E&�x����e�Eaܲ��|F˫G�ů��('�+�vj<����)'u9x�z�x=��k.�)>�cx�"�WrˋBS������h2�����5n�x���q�����*׍D�`w��M�n#�x2����g�ا4��;"�]5����F"g%)U������7]�@3�¥;���h��H����5+�\l�q�B#����S��Ko��+����LA��d���8��N��%�\�ڑ� �&��
X��<�M�@��� �C;&��GlW��1a|Ni��^�cV5�bgu5������iߊe&�4Mޒ�:�=b�F�Ǝ3���,�K#n��ڼu�#�Ӻ�M/�|G�������ꣷ��,��ӟ�`�X�r�[R	8��iR�Y���&�r��X�ʲ�NV��k3�X
�4w��Q�j�}gb���sޘ.mh�*�k��7����T�(6���6�PWG0Ufė,=���?�zJʢ�gǤ�K�!/]�A���L������5T�XL���/�S���N�"�z6�#R4I��� ���x�@��ȳJG���ԙ��L�t����f�'�>eg枎�Nw��A>�ؿ��D� �ӏ�"�O%45�n�C�6Rճc���5��9{���M��2J�"g�
ɚ�%jt�&|�zzJ|�ߓ���<ɐ��������V�U��,N$T9��V��OK$q�5��eq�A���x�_�B˚h=/��%C��!#9�����2����!��,��)�� �0�u<�Á��Z�8ֱѨ���생�`���Ьꇆ*z։5 ��*���2��'�÷�:�0B����(�$$��؏�OJ3��U:/bûl�+��_O�y�y�F��{�I8�^����05�㦢|Ҫ�.�򖓝��mr��Q�84ƙ�ꉦ�4����s�Eur���K�~]t0����'���9O�=�y���յI�9N��m4���Zxs0q��7cOG�~յ&�φ�!��ƨ�\�ì�Q���(��H��K���̟��a���'5�$� ��"<�uΥ5;Pm�����&w��,�Į�K��}��D�S4HG��-�j�2}�V�5۾�ʠ��toc�Q^.���!.���������G�HdX���A]	�=���Gb���&ky�޹�L��<�T�4�9��k�I0̞o�;	�#���*��޺@��;�m��\� m'"򧵇�/�%�N,�4���R�cN�H��`C=��5�%&OQ��V��@f#m�a�2�Z�2�� �B�ղ5h��k!ѓ͖����TL	�]�gh^/M��F��D�|�{@'��U�U<Jp�6		.������D
�����@��:F��avSk.�j&*D2+*e+I��C��5�!:F�c1���Ҳ=�:r��&��R���4����֏"m�	��r����q��-�W ��g�0oI��"��ot�l,�x��0-���V{� bgژ�-�&&��������AR����ί;��~c���z%K? � �lo��_�N�V��<%yF�:�:TF-����cx�z�3���t?RXA��බ�:|��e5C*�Wbr��RxP��˒���O�3}�)A�Yq����<-$
e)�]��+��vUg��LPs�| *�������
��F��+,�`���C���@�,
�� @uD��q_��Ě���̩�D�ًo'+e�8p&����JmF��y�%��-	ܖ��G���\��l=�f� ����L�f�]$��r\�ʬ:�3C�l}��\�� ��z�G�!Y$�aEs��̳��
'�Vf,�^�+�����u�?�(�'����b�ʊcG���>�A�ءs��?h�S�6]��}E?;"�*I�����������ϒO�xӜdٔo��Թ"��@�3���ܷ^ɂ��k� ��`�yv�SJt$#n���$�@����>*~��;.vìݹ�Oh���s�mLk4]���n�VҘ7n�P/�Hm
'��+;yV�:4(Am��G�Hߊ]�]�8 Ezo�C7JK�=��,O�PJ[�j�7rQc<ǟ�~�Dȏ��sC3!��o�,>� ��Y�Ň�CR�峏H�G*�ǁB��W�ܐ���܃$4�޸U0��1����]��l,�6݆."R��ܒ;.�+8���X N>/0�;��'��05�B5�h����'B-�����x����\Z;
��OU��i���P�A��O�;34���V��e�����H�^4�q�Jum�ه�;.�m�x'A�^�q}��;���M�3R�=W:�{�2�,|!� ��I�� ���	s�c՜v�!�L�-N�JO�=���!�P�JMd�Ob�g��9�i5
Ju]}��HU������AB�E�a��R�!�~56���dkh=y^ߢ��T&5�XT7�w�/�����E��0KXW��_�'�j6��ϭ6��*�';�S��������g(M>F���̗��'��0��1T�&�Ɔ8I���Z�	�����	�_��il��w��tm�i��э��mD���s�F�S�i4}�vfI���p톇]��>�q����[l��HzFlD�1��5!���/ʇѣ�O��b��W.��<��؀0۱�'1X_f��<o��MS.�z�зZ�����&�x@����)�Zj��^���w�8�����3�~-���������1�J�S���W��Q�X^��	�Kvm�o�`cbk���bs��8�AA�xϊnO��p�A�!���'�W����{4Mَ�&�n��'�s�9��2��a�n}�d���O��o�}B�!ad�(�9����-�.��)��Ɛ'��[=��oO(��Y�8hL� $����~��N?�H�#|/�H�%^��Z�v�Ӆ��,�"��a�`�� Ҝ��"�*�j��$\:���:�e���<�|�w��\��D˕*�:�	���Q�/Q־)��	��IH-P���	e��T��^�w'B�+���~��A�}���%��S����ٖ٩�L���O�?���~<�6��@�K¬�$pÇ@*�ns�M�r<$h}
�mi� �h1h�iMG(�6���w٦�'~WMʳ<�.�WypRB2VD����
1j �����z�8���W�K���bOr���!�'����6x���Hm#�O�*�_��I����z9��Z�F�J��EMJ�]ڣ�_�1N����A-�ӄw��|=00w"�	u��C8k}LȸE�v���,pLx�Hſ�(���	j��P3M
(M���3��<�@�0N����B��Q,��._�~��iW����\)�!a��/��/��d�+�.ΰ_���P)P��N"�����h<؜�|8���/�2WB�p���.��|�D��Z���|��@�pD�ԫ�67-�E������ A���8���q�Wȱ(&H�T�����MV�	�$��1j����B+?,y�胖g>�� cj�9n�$���tэ�Sߏ���}:X��V�����$�,q��D0�)��G�O�WCóui1�
;��C�^�!�����ˇj�|������ZI�ۋ�A Q9͞��o��(~��x�ʰA��:���r:."t���	���YZ�C4F�w!�>/��c�����c�E��j�������:�l�����Yxi���)�Vf��r����[�0��5���k
1��^�<k��W�D���T#�q�'u���9JH���u�r268&�:~|��Y7~}y�����W&�i���_�.*x�`yV�sM{u%q`W{�q�t�Wi*�
I��wd������s��u�fo�
eO*0�e�I�ޅx��)MFv��������s�(�&���#�J���jn���̑}B���tG4�}=�񨖰�T*���ʰR�D���Or+�4p����� �G�'3ɾ��E�-�.׈�Hv�7P���*$h�o�u���c��������4��W��H�jNѝs�֩���{)}���[%��>�/� Rls�:d=��P���Ha�5�"�1܎*t�΅{y��&��X,g�MVM��s�C�A�4�fO~N�S.lӕ3Y����A����c��̢D��C��Bc��_g&�,5!��Ě��V��aL>y��7(���`�swt�pd���x捺�<�i�G�1x������&��NU����*
���V��S�p�>H7��	�O�<5 ��R��&*�2{
HJI��?�ԵW`�}��9�� .� �Ե��������'n��;c�`UYU�Hћ�D��(ntr�y*�W���3Bf켢{��q�@l���ژQyZ|���h{�7+`�VJ|H�W���?��%��G � �<�Mw{~��V
E�õr+�����{˧�A�e)�� ǣ��u]�h ��c1@k����/�L ?i���]�yX�~<�FL�	?4��R�-�������R���4�u�҅ ��$E'M����	V�4U_�#�?�\ym7uo	n�bx�Fp�]�û;Z��b߻�63'Jj���@T�U�ya������^lg��8"�kv8�|.�C*-4_��b�/G�=����$�>x�&:��\։�OAEl��b�A.h���R}����Bo��G�����HuR-d���m��X�wj2%�u �Fb����6�xͧ��[��!�,�(SyN�y"��!��&#���?�?�jL� ��g0��.7j�C�h�0��S	�m����W�C�3͛n��쯷D�ϒ�1�{�ò�m:��������i������g� �Za�I����/7g�Y�t�����Ybe"F9N�^�.�����h�aq!�-���p�&��q����u$.�EG�"=3I��!vG5U3�נ�;x��=�P�Ŭ�ЩAz
�X	ܠ3�����T�
"�Q�!�spcɻ�'D^�R;Pֲ��ED�Sw>�+2t3�[��u$-�Tm]��9#�!㟖�*��@T��T���v�ν�J����=s�ݰ���9����&��5<�>+�+J�ZH�3bF+���*&��O
��^���������&�Cg�v�Zc��X��?�58�FP��w�v�+� ����ՉX��jB0�V�{�E�����x�-ӿ��c�6zý��Y���}_����� tH�@�[j�AA����������6v���ۥ��Ilr��k�Q��>C���F_dv���[˶ɧ�nþ�,����ay�!���ׂr:�+=��rr���E�˒5y�MF`��0�tĖ�7����n?������%j��E%g�yc@�0m����բk�\pPr������Ŭ�ly�G)���%����V�ן���W��bB�z�#K�鳦�8�K<����i�� 3��)� �?2<���Cٷ���$���c�?�t
���,ck��D$Ɲ��bWj1�Qp��xW�/JF�@.�0S��@���ow��?�f��Ak�Rʒ[BZ�����5Wk��K��.�n�yD��W���<�(he��Q�aIЀy�}|�t�b�Ћ��)�b��pʻ̲|�H��Gk�<�@�m�O˨�O~�|bꕜ��Wgd�F��~~�jC��֒���(��)� ��QOv�-o�Л2K�*��uC�b�2#��
�>�o6*٨���{*��(�hsjʢ��+���1c?C�������~X0r��x� ��MTc���C%�5𢒒ٓt׽a(I�+��Y͘7��w�I&���P�ꭠ�o�.w�f��NE����C��Q��џiGM���z;:�yZ ��tcZ��;�?J/��&'h�cA�fJѺ��ޟV���.�noQ"�����qx�k�+�Q���3�� yu���f�?�z��]!�vv	�1[���Vù��v���z�6ʲ�*��!�\-ΧG�]9��ڸ�P��dH��ֿ�����j��&��N��Ͽ�mb�N>�A$t�����C��m����~�R'f�8��bN: I�r���� ��&��:i�\]������?�/��7�]����G�z��TЖ���墔Z�r�F�Z�Ӯ�T�l�?�*��?��1�|a����̽�#\�C��Z�p�2-���9�vT2A`�5�1�� !����,D�?�K#^EPJ�o�B�J�EG%�`�\����͢�q���)Ó��C��w�V"v1Qr �{�J���3�T]�;Y��J5�'��:�k�΋P�ڸ����A3���o�+�_i1��$[P�gh|��i�����������Ŏ��]�>���brH$yW���.��Z�Y���*�b�����!Sf U�����O�LB�Eh��N���>��ߋ��ZPNˋ�diƴ�z@9� :��wOS�����8iեW�a���-'�[�I ���s=/w2����J�]�ܗf�D�t� u�1?Qw�;�a���Dt�ŭ�Xgͷ4���)w�"�/2kW\�yP��{��!����'+=l���7��,�.�}�u>���)�ǵ��� ������T|5oLZ�2s������Yn�BH�W�-T��#�es"6������5�I����|;-jA��.C�6'*�;��ۃP�iz�i�I�K�[�w�_V���{�i��:��,�߽m�.l�6��oZ�t���)�b+�Ggr/������8�+*c��CĖ3�����ĸ�X�&LM�pN�ڹ�5��<0�A�aQpz@�k*���!��(&W�ƌ�a�sXT���}��/T)�8rRQ�[$�J���:��R�.܄3H �j9���O<5�W�h'��)���8����.��B�[D��N�^�Ѿ���0	KY,��/)�!�/��p<I �ݭ���|��Nt=�v��S,M�����m��Y���W���ou*֜������ ̷y��	z�^���%W�\R;q�ƃc=�����r��W'�����`�#�{����}���i]йx%�;�� �u� [��%r�!{U����']�r���(��~�~�?�4]�J���@"���$T�\��7决��i��_̿�� �>���D�S�h1���cAo	��B�� ����GV�ܼu�XnI�R�q��U|;L�g;ӄ^B�z	�_T(l,��k��W���-l\�)�"˯�^V�NbE ƈ?�Bh$��!/����rI#��ʇ=����*M\���(��&�.\t|*r��}�����U����6K�~�7X��Ȧ�Tt x�f��,�& �X��;F��J���A�)s���K�e�S��{ۅ
@h +��_��$
�iל^ �3B�<'� �*�_Λ�~���%�m�H�Y���f��i5�oDtkky�}�۱���A�R����}���n���=�
�`uH �T׍�+�L�3�Q]��>�����C"$��]�޸K��uz��;���W��ݼ�d�FVc��f�IǮ*_E��/��z�}*�L�Ͷã4}X�$o�%'}�z<�t��m��L'"�}���P�o��g�_��A�FNW��3M1�l>`���v$o���j��j�8Y�� ���jٶk5o��c�,I�FR�d��ϲ
8�|�s�,f9ބ�^��m�nL]��YL���W�w`ߪn�P^�敁Mm�0䍚��T?�ݝ������uA�����k���>>��WH�߃��bQ�Q�`=�݊k�<���]m�i�����Ӕ����,a҈
�3�*�"�?u�=�Q��'7�����IC+��V����͗�>�i�4�R)'�/=��5`��ѥ�G�,�7�ƺ�?�$J��swl�o�.9��Jh���3˘.x�N���Ͽ�����Ye�V�<ٮL��s��Y���VB>e;���z3l�b��������5�/
f��蝶�*��A�&�&0p�쫞�dđBWxV�&��U�` ����Bm��
p���6��y�&�-B�J,���s�G��z�����&
c�G>1���*7E���<�L�Jk}���l�u��
�.ȣ�>qtkh��8��u�������}�1�DD|�����-�)����R�6j����o~�~C�b�UJH�"�b`{��eB����Tгo���oU�9u�M��c���b_z�iP���%F���ۼ�~H��~����*� hb�3�6�^k���1A^�����JKo�sj �>/��`9�*�Dig��LĮ��w����.�����i;w����q?�,�ay��K����km��T�3��I�>�<���V�3숊p-�RIwF�A����@,�e�@����PKC�B廻$y��%k��;��a��M�Ѝ���EY.-E�QM��`��m-�\�U~�R�86�5o�1�Â��O�a�p�}H_B�����7rI����}�)��MV�.Ҭ�桁x����>��gZ���(�N������{D���Ǔ}���� 3ƁN����}�v�r��
���"�D	&�th�<L�(,� ����j�1�c���J% ����dXF���s&����n��!�������mj��D��U<(�]�ga�gLb_�����/�za4
|(\Ҳ�ns�Z�k��m6J�jC�r^�/�EB�F2���c@0h��m�/k}����{�K�{C�{κ!�n}��`�9@s��O��w�L�9���-Dy"��J����8��?�q�
����o��|Vא�n��o�}k�1�̞�x]s����r���}(P�Վ�Z�vh��������ࠎA�Ή	��Oa���tNS�p��.�gۨ�,/��v3mR�c�($4"Rl,�&4�{��X:,���*c�o.L���([�I��5��`�k�`ل����>Hh&���K���%��uٗ�in�"4�q�r�1٫&��h$�����l���ӜX�: �T�X�_kъ���I�']߃θ�P�e�����T��6�f���}]7!;K�XBR�O�Ri�8���,�3��h���1V�tVR��h�ٸe�%8�$ѧ�q/���,<CNz��HL�1zC�����תY�7L��t�t��RwD�A��QW�����F��ȐI��5!wI�[�j��R0�QY�8>5���)�5�b/���zPi���:z�:�TC���B��q{�'��|�g��i4���7�+f����!�7�J~u���KH���}����mc��<w��D�F��{JTP(Q�B�`���.q���X�5��y��W�C�l}he��Fu���=`�J=t��t�]Sn�ے�wm3Pe�1��0��8�SU��t�+��07�d��F~��9�<�~`x^ŧ�Bp��ң*�i>7�N�h��0�]��G�m�����R���p�6St1��͛�6NXYu�e�������2�B���ʍd�?D�Kj������V�	�)�p�w���?]ٜ:5TQ�6�Jv{�n�����7��8�yH�o2H���̺T �T�i��?��Q�!:1���7כ#�����q!�>���j�g4�+��=Љ�I"8�g��	oh'L�S�XS�'p�����L���>B��߀U�dP.nK'lӠ���(	,p�,��{�"�۩	�Dn
�I6@-�^�Kn�}�x�릷^�?]a{�Z�^�苜���^Q�Qi�LdԭŭQ�<�s����x��/�3�f�<.���[e>��˽"��{H��@��/d��@}P��"UoG���E�Pk��ͽ�������o��ɩ�1�@��JL���k����ޟB'�=�9�y8�9'	�Q�SQ�&���q���#ф0��O�
OFa�r8R��LB o�~�Ґ~�u%lQhWn('��#��aP���&Y��.&ا��N��#DcWlQ��e�K��o�.F?]\[�q.��O��E���]1)φm˺�|0��%�[�*��RU�����q�i��e��	��s�˽Kq�_o	����� tlL���;%�O]�Ѧ�#\�{��>��>y}B]�T/���д�R��{^�Pt�P�TO�@�n�-�����vl��h 7�	�_z$Y3��InҖ5�FlU�i�$uHuk�6&�����!�� �Ŀ�Fd���t2�,$��3i����%Gw�eC��~f>o�Vاpʨ�p�,�>�O��Y-�(��ڟ0yK��PtOv�,^w��۫� �y�S�~�yQ�r����\[1���Il�Aݦ_�B�%AZL��%�)Wq�jAEm\	�1;]�a�vj1����d<x	m|l�q RSQ�����>��O���� <X� �l��E�"׵�Ġ�e21���Ne��JB�)� �$�����e�b�)��1@�{H}bC+�݄V:�y������$�<�M��_�*t��4(��(<%�)�r�l#�n����lfx+��U�s��RY��@l�鉵YQπ��lu,F�DY�����W��.�V]�/U�/I��(b�j6�hs�B�!$�(�9e�(�pX���{(��r6��+t��#�r�Hjt�7�$�?����t��t�07d�U�̈́�]�R[i���6z�GZ	O�x����9����Q�t�J_�F�F�y��	}��X�U��|���_Ց}o�����g
;J��fv�!E�ڕ��AjzҒI���3O9O$���W�:�6�Ir�S,d_&$e��k�>�U��0��k}�<z
R/��l�N{��:Y���I3���Μ�H�I��py�a*ߤ��B/D
�F���OD�|��Z�nV�'���ژ%қi$���ډ4�:�2��j��璈C�@V�����K���Zj�cb��)ȴB������(��z�Eq�ݱ��];p	I�*��*�Y�炂�@���W��Mnq�^�z���rJB�M2f
��h��4:�Ԯ�*�N��5M'�F�~)�`YQ�v�S�����(�H�v���M�p�m���?����\􆇫�{����{htU��9<�F��m7@k������{�%N�aziB���SW` 'VV�A���bW^�������������\�L85���e���J�AF/��u۳AX��ڒ�h}g}���4��Y���i����]�X8�>���7Bͼ2xo��@~-��RQ������8d��.j�����'�")����˒�~��+��V|�4��!w_�HX��]�:,@lg����\��! |�'��LώS�[�2�=C~F�H
zY�7�1q��$���A�) f���r��eQ�Kɹ�j�FK]�f:#�>�@�_ܙ��;���+ȼ׋n�p�s��q>O��t���E�U�0]����Nժ+��{?�?i&������������e�d\����0���+��W���_���D#�E@�*Lk$X%z?|�{C�9V��9 \��Uذ���m�M֞;�	KhJ���z#�^�Uը�U��[�rVi@�8o��+���좕|���"������2�L�F�b� ��y�% ��r�)�,u�����z&C8�܋���|T�G����>W,�Y� ������BMF�F,�30LO��}�?�Ǖ���R/Z��X�*�3?"�/ �E8���6��x��3��'Q`1<~�y�0��R�v���(���g�=6�W}o����a�i������[���G���c�/���\�r!t�7�-���q���HH�f@'���#�?؞o�$�pn�_�x*���>���4%�h��p�����UP��S���N�:ѡ��4c2��Y��.Y���	Z�ڀxjO��yn��kYw[r@:#+��e;�?Ҟ��30�3�q���1Y�(+�uʂ�VU{�y7("3m�G��z�a�b�ҽ�4<�
|kc�{�<�N-(!�Q:��J��;gS՝��s>��[H@�0OM����ȃ=0jeN��	����@��6�Ne߿�,zBS�Ks@t���k|V�x�%�}��Cѓ>�edD}�Z�WK�ua8%���ă8!*�%pF��TV��Dv��1�sBb�]w�����j�76��}Q����0��U4 �e�+f��|�
�fkj�o�� U�ز�`��ϙ#�&�i��-	��_r7�6�D�J���w�5L���k�AzG�N�E��UjQq&4Q�;oX9�<���
�MQ�/6��9<r�qG��触]JK_1��hj.3j.$�P懇������we��E����B�+���a�������/)4�5q��q��14�)��\q݋�zO	V���Z:���a��S����)线X6WϬO�V�}>��@Z@�Q �gBB���!H #:ZI��[#׈��-��� ��6�� �����8�I�t8�$�s�^�%yAtɦ_Ga68��fz����E{��x];�3e�>-�,��O�b8�}�)P���ْ]*�S�9Zam$� �f���X♔�<&���(Ii�`�#jq��`v<�a �$�C�hv�Q:6��{��ѰI��$`��ݪ���v3s�����,�ig��HZ�D��0�.d�N*�=��ρH���`�&���{�z�A�4����X/p3�����k���䌏_(��J�Ʋ�
,;z����X�k
��r,�H�'n�(�J���08�,�&Qli^�����K*�o��-��-~�㉥��moi�W�U0�M�kp�d��=4��Ȟ���^o�]�ԡ�|,�< �~���.��v����l�������=��c�l�Xߔ�7ٰ��Ӆ:D��Z)p�d/�?"����m�����?]����I:��o~�.��V퓮,k˫�J�KId5�M��X\?ɬ� fb����-��u�0�A,��#�{h+�[�F�8��U� z�<g��e��ǋ>�Kwr}�(�u�Ma��tb9
�@��c�������N���̂�����N�x�z:i~�9�N�O�
S_��>� ܍vAw�3�Գ���ܾ��KM���@���`|~�{���qo�h���C��sDh4cW�y8T$��g�#�\M����`xjߕ\D���0�Ioc�;Fs���'�`�7��gR�>'ykm�h���_y�i����I� �;4�T�"6�f��0!y����V�

1�;iąV.,�n������)���j�5�c�x��p��iŗ�<$��)3�.�֬|ġe�Eك	�&_��a������?����p�R���̖n�&�EOZ�}�R3�+wѴ�\�ϟL�p
�?鯼a5���{x/P%�ʨPR�p��O�m.���g���1[��(bH6P8�x�f�+��v��E�U/zV+�(�g`
B�C=8]1~w�0�8������ʇ@�o��4�V�������Z�hX�A�?���1QA��)5kʕA�N��*LW�
s�+���Qz@���M@��U���l"b)�
����'s˘'�n��AX�Vkf�1�횞��0�C�O� V�S�{���U�.� .�~yH�]E�,v�v���6f	$�H������wR�H��\�>V��J��q��ērW ��ʊ�w�n��3��� Qd'�g�Y+߬�,OF�
O��7[ ^YRj����IH�9�#u6$��FX/�<c�;��~�3ė�x�P��~�8ռc��^��r�;"��Pɲ�eU�D��r8�e�,���Ə�%<+�1����Wy����zW�ze�Ǥ�1�dV�����l��Sx��K`���@<�{�'���φ����^z���T]�5�H�0����K��X�J#`3����3�u\)��TH��E�A�Hn�.��v��+�����ŋ~�[ڀl�6=�,�}ڔ��.7��;~�Dچl���h�M�-�l&\;�x�g�H���Eu_PP��JqE˃L�$���K�� +f�.�'[���J�)7�u��?�R����%+^�%+{t�+��F�iN I<�����"@�|u'�I���P:�p!?���*��9v�د��Q�&ԫZ<q!+.*�t� I�M���3ʤ濇�'��+�.'>ڶ-��c8���B�gP�~�.X�S��I[t´f�	��w��}���T"�f��\�B��vZ������2��4��ݩ�yZ�(5xy�x5�z�Q{��B��",
������`�� �m$�D���BQ�}�W>���b���������6sW���D�8��/�E��I��->�$`�p�"YO^1��0�P�>��w*���ޔ�O��f� �*1h8 ߢR��V �Y�k�Q�Ls�Ѻ����\��b>��U�Z#�u5Y���q�������w���`� ț΋8Z��t#�p��R�,y�
lm**�(��j>�?*�3G��o�����=-'S8��Y�o|tt $���9����& �|���g�u�Ij�A��$#b�;���]g�_�g���'�u���Ls��_y@X.�I�e�`gc(��}��J���;�v��I��cć���a���JQ���&oݴ��IH����
za�M��J��k҂jB�gzU��\���g��/w�6����<�f���Uȥ���3�p�*�;�ⶵW����l}�{��WZ��"]q6��t��6x
��Tu�\J��x�
�j�!����	�S����<�nbN��w~4i���PM�L��TS��?��+�������-��$�I�]j\�'bg�h5\��b�Wn�I,�<��4Q��EU�Mx�
�3p�Ģ{i#{]��}��_���-6�U�;��.ԗM���*�����P]=��ZJ<�~y�\c3�̚�v#��6�%^�� R�	���8?���Ɂ�*�r�����`�_z*�V�x��\��BT_��{fғ�EӋZ��ti��S�q�H�C�a-cF���6S�&�C��~���r1B���T�$�	'��P?/5-ZO�|&��`���� ��#��x*h�O�<�PZ=�F�? �"0؆D��8�������f��?~�(���T�@��k���'bA�$`�Kg��2�I����5zK:�~k����`�-�R0��e3�SU�T�x�+x ,�H{����N����_U��d�ִK�;U�1��ws��* �&�[�\QDh�z��4��zY/Q4��7��k�X����9.j�����n�3w�\���{�qLYbS�H�Ý[�v^��� ��B�w�M1���>�ʳ���<�W�:=��{��I'��?�}ˁY��=R��H1|l3�(�^�L���Xl�-���N�]-�н����4%�ӟ���cj��:
M��*� �"�2���)��«Ys��J�XT&���� s�/u�U���R��1�~Ar��uB�:������(��Ld�r:���xd�C�d�y8
���r&�~U(�4��2o	��>y� ��){ke{!�ɑk���jk��(���h�II�EWABMc7R��>\	D<�K�b���5nFe'=e���?�dE<2(4���C곦����$�ֵ���}U�uDp���_Z�$�)�L]����^u8�4R$fe�g�W*����=��=����W��"j0J`�薎����R>0�T��^��m��B	�X:r�=eOa���U@9�/c]�U�����f��K`�@v�$&\�j1��� �*���D��T0Mb1��5{�)�n��]D1 ��fJ *{��4�  w#Q���X/c�Y�'�G�*�f�h(Yn��ڤ�N�?N���h�I���,�Zv&����q�>�9:���]N6m�f4U�؟b��Eɷ��6!�Wt��~��6�����׆���v^��5]��x�2��?N�֏�{�:�(�}�<��_�h_�QXFz��}����4�6Ϋ=����e�mY�x.�$/'�R�͍f1��y�},V`�z� ����p�H�
�#�����hΨ#�.���,�Ŕd�«1�M(���߂���'%��C��Z��a����Ȯ�����g�rbn�@��<��toq�sU]dxe��Q��v����@���b��X�4���is<@��+`"	���5�M��{�Y�~�Ǟ
�u�`�_ݽ��j�~��\��,R�f�:�� �:}����;O�E��ԥdG�6���O
��ڀ�n^����D�1���R����}
p
f��`TlyJ71v7�'%q����Eȕ)^�Ⳛ_���$��0��6�� ���^SP��iw��5ۅU�hO��]�E��
S��0hv[�d؃V�d����:NѻJያH���H@����&�3�D^��令f���~y�!�P�j�bwbN��
���X�j=��}�V�Z>MVY8�v����1��q�c���ٚB�ŧ�p��"��-_�+ؐq��ٝ�!^\>��z�U��Bx��Y�y�7���+&�	�X��m&|���[���]�A^��!|*H���_���������[4�N2!2�[�>8ʨ��
��J�Qɯ�;u)�x�ls��6�0z�Ad����7�I�N�vsܶk��~�b�R�H2
�0a&{��K�Ľ��7&2��&v��F[���i��������1];�>A�{��k9"����]a�ޡ��m���8f����'��_��g��@�sloy#��p�'�������C�\��IyX�+�Ȧ�\nq�I���N��!��[P᝝�X	��$C���:�����t������5��{��h���&M��X⽝ ��zyU�<$-%� ��`��;-7�/�;6T�ʚo���9�dk�� f���T?ҪǽQ}��wB����G�dl 3a2>��~R�ڌ��5��bc5(S�%�9Y l�!R��-N:<^ Ԇ���o���oD��&��ci�qg���<�l�r�fEB1D�4�a�T޿��]n�3,��{�;�i���%�ibߛּ�Zm�u�֫ ���q�zZ�+;I�F����@(��IP���4,���W6��Bm�p?Rf�R��!Х�'�0&����%���7�e)kX�z��0�DfPE��8`X�*Ձ���@�.�0��>��f�DaAe8� F��	�(l��$�"D8�g��V"B�N(��ŘZDkr��{�ן�,_�f�� @��Y[ċ wP��5��=��� �w3�֊n��ʸ;�!� �I2es�r�icE#L��r)�m^:=M������w�!�r��ٿ�KҌF�O�Y��Hʒ���DP�H���HqH�}]2��5R}�r,�*H�e����9�8���ښRڏƚ�j�fy��;j����M��e�Z�T/���$��Y���*v50n��}�'����Ң�HA�!}�b+���8�2\ѧgy�����3Ǐ�hk�|}��K�Oq��=�s�]c)�~�lO@����l�e~F��W�8��*d�+�����^�y����"����@��1-���-����4���;΄ǽ_C���A3ӷ�du�ָLa���ߦ$$S׈��mUҿ �I�1$R��n{���ܥKJĤo��o��4�"0�1.?z�)�S���m�Ƭ���7���:TbS��$ҭ��+�0-��k��k$\��p�6ۄ��.L&|k4�N(6�Ժ��ӟ9푟Uoj!���e���prn�IG���2#6uIF�_F��y� 5�,+B}C�^R��a�[O�u�2QV���(lN&�Bz�P�]��M=ZuVX[��ۤv�"h\�kJH���	^Ҩ��͙b:��4V7����ڀ�qw��t�>���B�-k�D`�a`�p��aX�}��EB�}r���a$�J=�|g<A�
���΅�5�c��"��\"A?��&�HN2���pHiyF�X>W�CT!����E�.0��oLJ�m�WW0E�IHA�?�T�ǅ��cYt��W9(�9�������8�WT��ESO�B/��a��h�l�κ��)y���}�ؑ����k/[C������y@�����;Q�l��SO*��7?�t�9N�S��1
n�G��CT�C��9n���;O���~��ߟ�|��T�qH%GĻ�E{�
8�k{}1�|�B�\�T��#ɛ���yO/��� GF*U�cU2��0Z��z�en�n�@����jg{���o��+�-�6�����e�2�X]�&�m�ŷd�m��� ?�0ơ�þ��~J�p����Hag��^k�� -��������IL��S�k��E}@i8�a��2��
#GVr���*:��Y��DE������ȡ{��ϥ��"��Z5"�P�^�u�^�XӀ[��P� ���mA�.cW)�1cAtƟN0|�d�25j�Rvn�y�L-z>@����4��K��:�MXu/$٭��5�i��V��G�6-ڊ�WCmvL���
N����TA�z�����F�cqf��K,(У�Oת��O���T��u+�@X����ϝna �C�<�P9Np�>!\�X��h��B�*;��E��Y�����\J{�j������ħ��`M=�a��:�ߛ� �*PDوN�V�]��t�pCMGk�E���N��"ͷ-q�ct��hzI�*�uDkε�J��ٹ�x�zhO��"��?�������;�aՍ�P���ֹ���O�����K�ly���{�r D.X��G�����/˯�Ǫ��S������c;���pqn�> �&Kcf��3<]*���Q�K��{Q>��"ů�I���z�?[F�j����]�<���,�$*c+U����@4�q�1��0?���N�d0?��8(/����4ڜ����9HA�L�W~�oa{�cPR<N��=���;��L��Nq�6�L^!�bd겗	��̞t3��\�3�k��5hg?w�#v4ݍRR z&�����D����M+io �/`�Զ2��~d���D�'X�� 5�i�ǥ9��R�@��o҂2�r��zI�M�jB�ar�^��|�>+mT��#g���]ɔ�0�����!H��0�dR�J�o�L�c����V�۶���=�Qř��$6+�JQ����7�#a:mԏ�o�+��a�*�N&�'�T���gA)��dhg ��E���דB[��X|�7��i6���Ӓ#�A�K}��۬	^�z
Z�wwMa����
����:A��\-�(蜇��s�͹.�g������T)��6��+�(
�`�>�`��t����v��0cF>���������_=�-뗉񄴊ʊ0�A��S�����@��T@��'�-��f��uaNh���r���N�'ws��+~��T�W�a%�yj���3�]�f���tM��Lǩ��&�h��\�� W�֯D� �aB@�Z����h�6&�|���b �	2ŹH��c!��X��xH�{�.i ��Á\X6u�B���9%_��9OxQ��[�1[:e�I�����@ %�jp �?���|p����t�x�7�b>��X9p�(�}��DT��r��=8j�Q+4s�_���b@95�D��^�_�t��A�;�Bb`�ڠ���n��}4��������2/�\�>Hd������I�sn�ڽ#��D�Ds��E�/fXa@�$�]�g�8G�e ���a��u4Z�K���uG|��8u\7��zgs'd�� \ͅdu�����JA�������>R)I���'OT@��]㻓7-��I�j0ƍU��3��Y?k<i��2<(�%G9F�s��7�nh<:���ZMI�E��,Q(�F[���>28q*�|H��\q6h$�2����I�pEm���`�*{��*%ʪ��#�����}��]'�KNV hڟߖ�n�;3��Op���1��Mm#ǜjLrrǻ�Ǥw���N�\W��- ��F#f+3�}�7��lA�i2>3�V�V���/���l��$���$I�m�<=��{��e�Ǉ^�i ]�4�P��W�w��.;0c[V�Dt�΀�{� 5���ؔ �1��u5{�LMl�E>�y����d�7��̑��p��:�<�暱�N���Clc�O�<�}4���K[��O�gS;��d��#�;{æ�2�;������O�LP1ɳ�Y�����1���Z�Nt��$Z����Kw��~��a�g�G�R%]�m�*��P���D$$rY��;&F~��e��2+���-��ɘ=F��sϛ�O���NxK�>q��>��h!o̒��Su�V��#�!�4���Pו0���I�2�)a�y�9*�W�j�K3�*îiA'�֦{�i�1S�J,��\�{+3*s���C$��+�ٖ�Z������fUf��~��K��������A���/^��F_�u��a��u�\ �٬y�Čm�J�dD[g�?�,�C�<����������d^����KC��6�?���E/x���?�u�[敁�Ͼ��������֨ڠ�����1諚K������5�c@�ۉ$9�jT���zH\��>b^�n��X�$p"$�R��
٧Rh�o-��y$~���#�1��0×�h�9�H�@Мp�I���-��\#K���T,�k��%�1��	(�G��:�s�tl/�P1}'��p"ܡ"�|�0?�j&����s����{�q~�ݘ���ӯC�ԍ���R�/��<.�*�-�
W���j�����0�ކ{�t "N����#�1{�����9V�����;v,�}�}? �5�1ߣ&�j4���mL�-=K�^�aI���ƺ&���OQ_��{s�F�3��Eܿ�)� *��X
Wd.|0r#Χ!�m�Uٲ������n��~���x�ywV��k���,cl�S���i��h��]1���;ĠN�3v˚���T�Nb���q�)px����`Wb��L(Fw���*J��As���q��jy�oy(s����hCI��B��ZU�\�of�^լѣ{=$�+�	l�-�$�2�1N��ڔ�z
U�6�[i�݅���|&�l���"�G�����AT�[��t���&a�� n��C��D��0/�H�V�� s�`�'���/r>�%~;�b���62j˫�o��-����*�4�@Up��I2;+A��,�'7�&�;�=nV @�w�ɗ�:<��%���������Q�a�"�t�&����yAF��]�	#%g�]����ji�0�b��y�y��k:�N)�]����;������Z����2�����:b,��`v�����>�[����ÊW�!�A�_U6Xױ�<�����	2�ă��T�#���S���0�=5�y;������/�ދ.�~2h݂���{ ���3�)����,�z��������� GaQ�U	F&�|DH��ݍڈ��\�$���_�QK_���ڮ�d��p�@�hn:b�[*%���z��=:�]�'���2���92I!�Bѹ�ř�<߷ҌA���V���Sc� ��~o��]�Q��d�jئ�&Z���A�H���2�uK)����C�/Xf�ڄq����MӃ�t	�bK{�<vn�qvsp��]q=�����6_&�s�T&͛Y?нe�Y�ϑ464w�~-���DB�(������=`�/�AI����P61�f�M8������ �4D�l��S�W�F�"������{J�	Ec���^�� L�� �6MD�������|K��-��$���_d�c��F��*��`�Iڟ\d՞�d��h�5Y帻~�������5Q���!�0fCc���N�э?Äω7�aL�9?�RC�(��I!k��`��)�N�A��?/�F����0d���^��6Bm��S\�G1w�d蚟����łE�I�ȤM1�CG��v�� �
�Z�1KE��ࡒ��[�z��ܚ&8\���^�R{(��I�s�n�Q� ��yL�>�������x�i���A��*�|��� �u<?[�U�p����yơ��W��HE�S�����|^��#��g���
wْB�,ؖ0��{W�s��:��%�����t��b�Ss*��E���;��8 R�G5���ʔ���>:Q��5�U�/����1O,/X#�,�/���peR�}�5^�u֝S�Usn�v�ҍ�fg� �E '����E���$B=��L�7O5����]+}��g���������4�3�NVFv��(���K�¹�"�yf e�zAk�Ԙ�g	�����U����h%�c��6�(�&���g�ϟ'��V����;���s�\�7),Wl�w�u�Z�	`=Q����h�I���k�����=�~�2f�T8�bqL�����<�������o�J�~���£Zs���!Qj��!u*3U�'��Ãx�DI����K]F+A��$�6W��T ���Q
3y�3���|����v>���F��yf���;Ou�y��bC(�j!d�84#ICo��G���F�e@?E�Y[Ƚ�������~"G5��h��x��9���ߝ D�|)N�o>�T��P�	���^�F�h$p�)�$v�]n��@ycB�!j{`u;��H�)�A1�3��C�f��T9�|��[1Pt�7%�Y�v� ԝ�(>	������;C�ը��l�E�S�4�?m��ؖjB��� �|����7���l�Q�6���G�4ᡥBf���9�H`F���� E�Q-J$h3�-s՝�"7���0���+�R�=��W�dڸv���5��J���Z�L��.:�'�pp,�v�׭������L�dYw�R�. ��G�{�-�S���K��}�C��}ӆ�ЗT�p ��D՟.(����(�+j=��s���EFh���
,J���U�Z�b��޺�0����"%w�s$c�p$�Q7���tyIȫ�U�͡ҷ2�Fsowg�!Y�A�����W��`y@�o�ˣ�H��]@��	�J��V7�D����w��C��j�468����5�a��S0��e[1虯��=I�89ٙԄ��&���遨�jc2e�*oM��(f� A
�x�� ��vDG�}��QF��Z�:����c�02q|�Nk����z�����mڢ��o)s�B��>?�^k��0R�x�>`��@V�78��ĀR�_|&	�%����K�����=d-�����Lf�rP��Q˶.�����G�Z�Xp:P��[�����P�5o�6��t��̤�#?���+�èe{�2�SYׄ���-T��3�N��n�L����|�>�:����P��'kZ�8�P�Z�wyl�)��ȉh-*h2t��,[8d��ʓ�tc�ŬT£�1�w�S-ũ��z=��.�s�ʾ�%����^�4�oQ��>��|6;����k4<��\�|a:�02�]�bb�7�\wJ,�o�u��l��Ǥ�)4Qoôm�z!��?����Q��a_�����|5�溼1�
�6���[ �D=/�$�{��jr���\�b�Z�,�P{x"�x���8�/I{Kc�m�=�?Hk��z/W�=�]ڋ�f�R�d�K%7��}�N�� �ޘq�W*��qS��\~D#h��"���rGJ��e�򵚲\��S�.9�ۓܩ#�<� 4���i�D��ݝ�pSj�66��ؠRZ﭅U��ܗ�z���+v���C��u�@�fK���u�.'�~��4��ED�Za���	+����2,ճȱԺ�<�|� VQ64�=�����4�&���ilʶ����G�ƢKB��(�8_��$#�����ՍD���-g����"Y;��t�� �nֳ���{�Y���������	c{��p�N�|�(L�|t���$�+}�Qv��Ȋ����ʼ�l�,;>��~|�t#R�x�`ˉs��!�;:E������ʜSr����O��Y`vtTI�4E|y�_�/���w����6r�?1��I1��VR���|؄#�[��"l�/�
��oF�����r" �G������{}'�`Nˋ�{v���^��LKB���)�T���E������|V�T1�����[x����Fo�<Ə|(h�/J����f�e�H�v,��Rt6AĖ�6�1*�E��{�u"F@@c����~�Y1)�C���7�@�C;�,�Z9Rģ����� !�/B��LPf���X��P����O��F��"�ܢ	TI�����w�8�5(ѦW��;�aw�%m�i�]<���89 �)���S֯�f���65�J�ݗܶ�*i#��;7�M*���ax��}t�)�Be�L0T	�]	��:av�*`�pY�ްx�»�Kڂj���*%�`���Q<#�ܨc�D�&�7��8������_M\��
.>TQw���[��i`/�"lK�O���w��3�dʦZNa\�^�^�~�-��&���?^���t-Ɨ�!��yÿ�"����,�S���T�O6Շ�0�2X}�(X<1���GY?�H��p��0�O��OW���K��>&�Fq2�ܔ)!���{>�����)8ʜ
F�@"_�<{3���:���psW� �{��75=�e���#�&)�i�A��L��"��\�n��>�en^��O.��)�"��`��Gd��30;7%�F�)Վ��-˙�Ҩ�Z���Td9�W�^����������#���ն�������C�He�rƠƇp�9tUƋ!���4��V.\��`GB�)ƞ��t�2����z��'���1�،W�0������İ��1.�^�뾾��F: x��
��{�sۓ��`�Sn��bn�[��׊7ۥ��3̧1k�Q|�����Kdp{[7�J�gO;�R�S��L����_ӄ=��������R����%�M��e����u�a��xFo��d�%uq�G���	��t�M�����$Y��%����G��5$^�ڛ�k�)�3R����U�*T1�����l���L� ��@�
kr9��օ��;��m"�o'QuN+&�R;Nc����%�q?�i�/����a�ZO�s�������$}s�l�<�%��:�`�g��̍W�j�Cۂ�8˶g}�JiY����������� �D�4 ݍxY��&=�������
i׾� �ɇ��_���m�ō���έ"�����J��8K�-$>x�����FQ^θm�fZ�ł�E�l��'� �'[٣����B�������� ���y��4[��v���]J����F�f]�&t�a?*�:��̺�a��n��Mv1���k�m��2d�
�=٭�{��"
fvZ�c���Gr�bh컫�<r�����!�R\0T �MŮ���[������%��
���r~�S窺���,Wܿ�m�q�҄��8�&f5�}�-Xpd�;�na�0�~�Q3���v��݋C����4Cvq�|��Z�O8Ud���D�Q�>�%3�U22��w�+�,�5i�h7�H��[��,�.#�}f2ړs�Pu9�!�*�5��GHm���%~ۗ�uD�:�,6�(�%=�=�I0���XO7p����;�0��fq`�ƣpH�tY�,��2H���ǃv&Y������PK"kI�p�T�4J����Q�˞��]�40�}
ӿ�؃L���s0���S� �������VxP�����{�H��E^��e@��J�{ ]~9�XY�x���-�d���ڲ*�qf�ĳ��+(V�:�,x���\�s=K��Z�	ذ��p��z��fi�)>%p�5���ę�jU���<m�6�݁��V%z-�n�5|��7�O45;����S�
�� Suss��DTv9I{��p��?A�!x���/�Ey�4��G�i9�N~�r��
���#���xib�"�z���v��Wᴬ$�Azq_2zФ�wԍKN����t���ʨQ�uu��r��+�����Q|�dI|�^����+�5�_Ż(��VLj�,��؍��І���i^�	��{݉d���Q*������8l��^�
13I�1�1�aC�7�^mM��\\P*���=��b�$����wNAӡ�P�-�xȓK�碔�.���S��v��D�g�WH�L�͒S��i���Vyy�:ߧ�h�͉��� �vf��@�v����[�;�J�FXJ�P��凗�U�QJr���H,[\�%�nf�lc�Ԕ5�y�24$��'�$�:'Xߛ,�7��]"�-�����d��"�C�pe 5�U��\C���S��M�=�#���� �Ʃ�	b���Kc��h�a�*)���ɶ<���Z8�s�!�_�[5��I3Ъ�D�賟'PN��7��1h�E�Ҵ�i�E��4�u�� �6:��$\��QŕM��O.,<H����t@�ߣmҧ��[��5�o�e������(١�����[<��j������y�+S5s�X�3�TJ̝���A�&tL�L��������t�hge��R�U�i�kT��yuY̲t��q;�ܟ����z��K�sC���?rp�qE�ԥ���l��s�zsd�\�Bx<��0�C^�W��U%�T���� �w�RP+��H�[�ǨqO��́�M� �-�PQ�ms��
���$E�J}� �.�V`����Շ�C!��R��}���������k���8��㮭�W��l��+=�;�~���P+F�FW�ۣ@��"���e�`5�Stz�d�T9��Y���_�7?8�[�eoz�%QQR����䰎Ox�xF� %��NzI�(�l�[A��Y=����ϲ��;+*�̺������-��	3d�ֈn?�1��i5���O�߷��vIt�98�/,6��)\��@-2�('$#�Ǳ�?�Q���cgܙ\���7m6��O�T�6�z�5�hz=�V��<�<��������X梙AS����}XG������^�ue#�&�d��Y�+�m��T(�!$�>֣G�~�I�W�8�5mL��!=����$��(v���;Z�\s�ꢒ�(��N�{�!"�x;�ۯ>`ߘx�!�#muG��u�*H�N����TB�0$��6=
i���Wc�E7��KC�_����`Z�Ls�CPY�e����}ՙz����*+8;R��ڃ(���@�����{R3�f��d�l!6��\��g˂�k�9�k�����/D�aF����q��M�B���h R����S2�����$p���!��W��{�
��� �t4Fb�Ė��[F��ǅu�<��\G���I�LÓ��u�UC?Iq�t��P���YD�Q� �����H*~X?���(��}v<m?�	����^66�oV�����Vvb�,0�W��w hbg��<���g�g��C����ؾ����;�"z�6����ݎ��K�OӫiyL�q�)���r]o�	�s�QK�r�Vk��4�u׬24��_U�ǐ���3�i�B�B�	*m���ZNfI�x ��,�Z�v�p�=-�V
��]�a�_+���Ȥ֒�8�:��8��Mw�֞M�f  ��^c�5��H}���l+���(u
R�
S^2"R�\���K'c�l��f�WZykf"�ݰ�t�~����B��o�%<�u�x1�'�]����$Q������%��f�$׽�9����[[��ve������'�f
�K�/��j�R��1����Hk�3����FV�d<kd�B��m:�#���i{?h@c#�SX�����[��������"V��1�C�Ԧú8�K�g��j��Ai;!<�b��C���^�	�����φ�$so�bvϟ����c����x��*��{�5�k�eU����0=X4T)��D��j̏��k��6V\J�\+X���f� �ʳ����u$�h쩌AB����w����v�����d:���y /�@C{V.��:�T����8�����ϳ��Ofё��xgt���J9; ^�ß��H����_���n��	�S��;�`	z��sD�\��OP�S�D�@d�WMȺ8�Z[ёW���}<;�Ti}�.�P��*��/������[~t�v��4-�v���D������<�z�H#t�����ڱ�i*P��H��̃��q��~��~��5ʳ �"��HX>��e���������������4a�V��h�A�wѹ�K{+-q��\��}���2_�t��O*��V��9:��ౌ*�'�,�t]K@[�O<�v�薹�yv=���=�3��4�t�I�Z'�/��ӕ�Xa����.Tn�/�����[Q䎮:9�׍�{Ġ(�}���z=�=�����Ew~&R��"پ8~ز���\sU�c�piAB��L!�
*S*�Ư�z���CcZ����첞�g?⸾�����2�)g�D��fr3���3��P�!R�����Xs0��渵��)P'�U�p���D�����$��Je`u%��J�ܶ���5�����h�FW-�'�,��z��x���W���"�36�)6H�
h�h��*ۘ�x=.U��t��\,ˏ�ل.a�\���zҋ�R�8[O�^���8	$����b뱢���"��p�QR�����'���.���(���A	��Ѕ���ܐZ�>c#��N�����G�%�O�--9�C<F��φ�ܴ��d���ށ6t����QdU�*�Z�T��	x����}Λ	�Faj��]���+��$�Js�]�Ԇb7Mߟ�6�~Y�����[U R>O�8c���n]I���	�xq�����;;�S���Q��%~���
��b[����Ԭl�i��?H��/�/<+��0����͎[�����Y^��I�2ݍ���7;�	2���B��P��9��3��`\��i�8�9f�bInc��
�M��H�����g���V@�μ�y`����0.���d��eKNtGd��~�`QQ�[��a�*C"SK��N�cPy�mmI�ώ4q3u�Z��HH�+��t(D��M$0N+>�ЊLi�������H�sW�E�~����%4d��*铗�H4;������RX�j�����%{��\KU��5��������볭�ħk������[��2m󐣴.d6^���4l���S�}�='�U� �45�1�;�Epl�6��)�=c0�����ۃI�X��{z_ /�HN�	�-�f(�~����%���g��s�L���"���n�v���v����r�7��d���}����q�"�L�- ���8n8E�$<@I$<�c�A(��N���S�>m�0ު���\���Wn���N�~�Dӂ�sČ�`�aͽ�J t��s���8���!:� on���v��z�%z���Ҧ���k���T�C�"���>�����Z���S����}�D����,X������������	�9W�v�KyF=��������<"��8n�C��~k&�sR�^Ñ��Z��Kp��%����c;k�0��N�:RA�e�U�/Q	s������&�n��Ñ��0����Y⿮�[�W4�7����1��r.������`�i���}� �^����++�LΖ���F�'C�j�V*���m�O�)�ʯ�QA�}���E��G��R�S���p7�t��K�7�]q\�p�����?�k�a|�-�
q�l�D2��.[�+�
��Dt(=Z OUL=��� ��6|:��\��ҢEU^;Y�H�mQ�i6�Qp�]	��5�ac`�95�⌥�s�H�l���#���'�k�v
�Q�;>B�����U,�Z�q�h�����6����?3��yi���e�� �p7��Q�z.XH����ݖSWңuH��*>-X^ʨLvMo�N�����p2#�?s^l��]L�Hބ��	�ٝ��se	�-9�M��
����r_C��z��7V&�`r���v�Rڏ�6�@tR��M��#Oȇ�5m�8cn\���zD�J�,��9u@�r������u|,�J2û�!���U�I�]|��̓b�h�H�y%��]�y����&K��>r�DԪ���uV���O�����}��aAa�׎���8�>R}"+!hzu���=,΋�_rRG!C)�Y��E�ʤ�R�nK:5��1��U�J�MG�Z$rA�=�7��.��Z%q�O�g\	�v�X�X�%��dR^a&���O�ҍ]Fk���������^]{����w���ik`=�&�o8w���Fz��'�e���u�~�m��n������'��Q���l�鷋�)�-��߿�&�Q�\�s1��G�R�X�������I��t����䳤�X��}=�/�G6��Ž���(d�Hf�g�wYT��!�h��o-Z�@u�3u��$L����aaW���yj�5b@���wr#�i���R�+�T�T@)Z������)������&�lH�~W��.�J��g���L�%�n�&V�l�BY��&��:RP�ʊI�X��%�t�#X���7�@ƫ�h��f�Ԛ����I�<�Jo�B�X��Q�B5�	S�JT+��sA�� �u-�Z�R��\N8�E�m���U(՛��l�5��.�#9��i#��oD�{X⥜bċ\���;�C�б�+H;o��������O(����ܙ�E
*S I&P�w�7r�;Qj��t2[l_y2q�Ц����ъע�
S� ��W�=�5 �\�n`ک�Vi�(�H_x:T#es�T�)�'_��%#%M�5�It<:}����ib�Df����L=��]O�
m�}Okm �>=��ɻ�}LMʺ d>m���ji��}%$nH/3��_T���3|c��YwSDM���{]�)��/b4����R0;,�z�Ғ���i�L��E��kFg:�T2qw�^�^��Ob�E7��
X-E��Pgu�EA���b\��i�,��ʂ����ԅ�9��OnZ�4
�H�~ԯ����%�8�l)�'��?#h�G~&�6P�-īƆ����<KrƔ��O�pT �6�3%��8|[����dBqs}��Q�)�g�ğ�9H�z{�x+��9WФ��4���8�ohLg���N�r�.�:�E	7^(�o�B���zSD�is�[�tnΩ�d�Ʀ{F I�o#o7Tr�T�FU�	Q�;��aMӑ�9ˀ�$�9�"�_	m��$�1Q�Rc��%K���e���,�fG���T`xY�K���[!�+�6_��x��m�Q%;;H�ά*)�������)���J�Z��P���Q�[��b�RQ:+����YJi��!t>,������A�:�h��O��|T~��l�*��sL��M1)��Z�<�Va��*�-9�)����؎+p�RPm9I��7�X����ĥ��S{/nw%ÍC���I c;������럋�͆Q����E��2��:�@Y��TԲ8/�9j%q�Jy�E[�F^	���"���Z�B������2���2�'ˉ�,_$d��kq��l<�y,��eݗ��'�G�5�P���Մ��@��_.� f%���E��◂��Lé�d�I���s��
n���5�%
�&��:d���L&ܯ.�l�fU��G���j!�\�w��/v�F��r1��ӗZL�����~|,Я�4�N����,�����e:{Oc���Ϡ\#X�U׶2��W�L��MG%���a���zo1��"��N2���֜���˩�k�)����vi����o�z���o~U��x!72�v�I�e����XG+i'bw�X]O�����b-�����#0�k��@wfϽ%?�+�
�	-���c�����uD5*R92��l�3�mJ\l-h҃(8d���ā_�� �d���g��[��;�m:8~��k�> ��p�0�̘eB ~�T�Gj"��Bd��jNcN����R����Z3R�a�S���lS1���M@7�h�\A�	t�6���k��Û�^׉;?��U1+��w�!;r����8S������9�B�$ЏzUJ�����L�G�<�@|	���\n;v-qk3f�όL���\��C����-�Ș����@�M[�}�e4g��#s" �NKjV�yx_�UpSj��$�zx�@��P�-��c1j:�pK�?�n���ﮉvyt0�'�%��`"t 	 ��eFR�7E��z���1N[��v҉��9#
WY�鰿�w,@ OdR_B�*���	� �\}�����G;�F�>K�*ަ�_-���N2��x�Q�y���kc����YA�':%*���R����z{�]u�+��|_?ɤ$U�lYanlZ�`�k?=��A��S���	t���F��N`�@Z{���K�=Mt��HoW�>6"g#��N�T���j�jJ/�����CϏ�uG%S����Y�A�)W���/k�e<Qf[�
�D��L�����W�In�1�b�6�@g,��w�y���\)�R��S�I%?D�B�i4�;��T�������%xL��T�����ڀ�c��;�c嫟<��]X�Oq��k�չ�p����&�I��� /9LU���.����.�t� ��d���y����$g뺇�ܳ�a9yX�Պ\��sb����q&a=�� �z��b����\x��ܹ ����<#r�����8����|�|k����	���_)0��ا�Sc�)��[T�Э�0���㕇��P<Q	�7�ę�"�*=��D�E�����n��N��:|�J�w��Jք��ي ����*�_b��!�N(��|��'��$�=o��E Uŋ���[��v6�c=��P����q�҅9��;�)���kA�Y�R�`R�z_0\�XkS����0�km3�!-�q��10��<�E\Zu�5�s3�+�B�W	&cꝗ���ք#�Xo�g�/���wLD���.����c��I�ncf@�#� ���K�w��++[���*�*L2�>�m��d�z3b]S(A�rYƀΉ���>�B��!��m��t���`����c�_Ù�m��5��҇�"ul��,j�ء0����/%�!��e�[��ԭ1��K֕=o�3*����,1vu��̵B�#�II�^��멫���mh���c2*Y{�sZ�~�I��f+�[����x3�Ϸl�~iVO��|@j�j�����_W�,9-����`�IA��W�9��bD��L/��?<r眶֛��D^�3K�Djq�؂�}3���]�n�[j��"�a���|�����72Fn�J]8BA�ƭPߺ����80'z���� 	���TM�R����I� �j���3f;�YaO�׎9���yl�c��q��2�2���VR�(]�!O��xu�]a=�v�n%q�Z�=�C�\�0~`Uv�Y�$��%2���sE�"Q
�4����ɫ2�a�a��EX���������k� o���@b�s���o�ǰ�z[$�U�(������dY�:�KQ4�)΂T�+d�OYj�i�'a�tw"��k��*fH�\F���o����K�a�|2s7M��-t�M�R���F�����^4��s����ҭ�fp��o�F+�E6���)�w%
����ۡ�������C�P������W.l̫��g',���y�����e�@� �e�S�x[���1�~:��\	��e�����D��� n�P,�dh��P.Dy�D�F3�/����R�w�.O��#��}E�Ҡ��D���Գ/��Q�l�E���i��T��ݍ:}XS[�����R5<"$�!�<��M����g/��o�a!yz%�y]��ŋZ�:pp��?�r:�����yz5�Jd�^Ē��k �Hp�YqA-��2��g ���6�F�j�ܗ��u�o6������g�7 [ny��R�)¡�V�s90I��Xi��@�Y�@��d��7mI
�(Gz�Vz�!��}�y�7���G���z{�����4t=�ܽ8p-�|[�j6���H�՜��o>"T_�//v�[�-k��o��*B߶Z6
pX��x�l�do�!��voL�7:}:V�b�ASD�#�F�1��c$����Z�{<�7:m��7^Oפ��1�Ju�]K4���b$��d�NcX@4��AY���2�_���z��+����e�Z��l��B� z��y�ϛ��ǌ��q�<J���(((�~-�ϩp��۞��K� 9�����C�MaW�ȑaX��lՉ��aG��~���`���w��U�i��E*��%?u�-�4��E��n��{��58�R���E	]CK'��̺�V=G���f�l}>�G�+���dM��K��7��[�𪑡��t�$K[죹1����[�y�,�:�ǜ�����B���	zx!���h�� s3�����	~����˺j�3�wU�)�sr�H�*�!�\aM�
�8��r��l���+͗�'��;��ņ��GW�httJ�~���6p�VI�z�׿�O�ril�=�o�[�"�l)��!�M�4�R�Z�����F�gD�}xkc;L,P�E"$y�h�C�{F�Ô�0�����Q�UBk��G����m��J���t[	�S�Pd�\��Gܿ��`��h�q�ؙ���c�� +�5�_�hz.Wg�Q��:��O�ht�WK��d��)��F$C��h���v�����#�"��Ru��}%̇;��:-�X��!ӗ�\HX&aL������RB��K���ys#���H\��1_m%���n#�(�D3��"a!7m���,A�`��gF�&�"p���s��o���  B�D,�
�Mӣ���qY�2o|��m�� �(�$�d�?�ݙD�N���lU��x+��,΢$`V>�^��N/��m5֌���P�|1��9�'=;	�?Dfj�f�[�� ���x%6��Sr����
�X#�Kb5���=Ʋڡ�B;��Z�M��#�x_��1�k�=#kN\�A��'Jq*u�!M�!����Mt�/<ة`�֕�y���6~�f�f�X��) ��[���3�3	v?���Y/���d��=䳨zF�f�U��z}�t��s�:}ӧ���>�>�@���S�2v%WiGH�m��}2�:�=)�R�I��A��g��
4�^�t��ěi�H!��T�Y�s���\�6�����k��+��U�o	Gr��Ιi>,�8��*��5�a��ĝ�k�ɟ��_{���)��͗����?P������.}{DO62͝,=�N�M��*Q1YK=�3��}?={���Y
�K�����Ȇ���<���Ґ�&�B;����@Q@eM��]���`dɅ8Ҳ�������B=����`�Ʌ�:ҹ��K4{J��a nz�W�Ĝ8��x׌�2�p\�Y�K�ES�T����� ��ׯ�+�@�b��W:��-YI�@�b/�]�GW��8
�3��,��[��t�߹�Dg�(����oDb^Y�l������I �NC�(��$�|��+��iXΪ��0�����g��q��ri�`���V�S��`]��4`�.���p6���p�M����&࢒����VU���{��?ua�����J!���|����4� ���~9،��}�l9 ��#��E��ܽ!QJV�&,�HZ�����9�Xn�:udbb��d�_�G��]� 8�Ӹ0bs�Oܶv�;�p���u�$�}��7aǈ"9u�af�G�\��9@Z����V5�8%l�+���N��A����;�z��+�CZ�q���5E���:Q�ᢶݭ.�81��r��>W����^gm�]�uC��C���%u�)"��궋�3��iW�FT8u�>����~�1��-?_|!d�@
�	Y�o���y�ع�,�����	��=]�o֨u�2/��,�g_6�B�*�a[�N�:���~]m�`�C`]
��Au?@$�+4��>Ĵ�u����0����T�K[�b'qSS���7I�5�2Eu-�hvw&�9�� KIշ����A��W2b���� ��c��"oZl˔I ��=CP� �s�g	�R��H:� �lF���n�-b#v*f*��J@W�%d���͖�#.���j�.�a5h���(��Z>,U�U��m���-�m��z�'hW]j7x�9��C�8E�*�
��:�C�@ڱ���hţI���LbB����w���(T�|�;��=�~��s╥\�e�i�c��23H��Ύ*�	�K1�'���j�6��C��rU��4K�#}��v����¿�ga�s\�r7����s��n�^�I M�� ����j��/Oe%��t�_�d�5�QHѨHr��h|y�,��B(6�w��[��5�bV˃��9����	�췅�}�-a̝���<����v��be;륁�dxM��p��jYn@і-=E��3�#b�h8*�.y{bĔY���6�x��~���-��#N�l����ɂ�N{�VWm��!Ǟ�Y�$��~�?�@!@e7�`���T��ᾘk3p�)f�{�$숖�"�J/�(HS>ԸE%��B�d�dr���w��ӾAdb�D�D5�f^PS(�x��9�F�gݯ����1��C�]e�ŪT�Q���0&i���>p�C�q>γ��Ԉ@e���?0��i�<ZY[�W��rk��rUw�������.�_/�ow ��w k�Q�?�!�U�:�t�^��␴����¹������Ou&9rXMg�cD���y<i8�yp�+Un��r�+�ي-�m-���n+u���iY�h?���=4 ��iӅ$W�<�l�Qi{����'!�؄����چw��w3�~/F�X�Ger΅��f��%՘i҉OӽǨv�}>�EA+�^���8��J��D�@��b�������U�Bm}pe-I��j>�'�!#G(�$�uF$V�ֺ�:�';G˂�|l�j��VJ��,�B���:ئ����Is<Xb}>ֆ(�������v�:�N��sS{�dK,�������㷆����
�S�P�!�eh�:hsk.K��"?է�@�b�8E�	ߟܚ_��1j
�h>`ɤ+7�vi�@L�Y�/�p.x�R����*�o��'K7v�����뼉jL*��,@���* �z�V��2&�6�i���w15����D�efw̞�B��7�~���sI��Դ7����!+�\�ࡄ�A1��k7��Ź��W��Qh��a��j*?)%0���:2�sA*��	xy�d��fzu/�������HTQ�5rB8�=@��Nx}��~���K����,��٤�B�����q��sQ�/ԑgC�F����jf0$ָ>���K�E=*5u�ĸ��
�U%%E���X�U��$H����)�~n5E��X�$�9�K�*����&�T��◮@��I�R�CN�6�#�A9��������/�u"�~*Sm���&!!�	V�k�m0�S�\l"]=�����+V��ݠ>�=4�@��qf���h�p�� ��0�5�R��5eiWzZ�^<KÆQI�(��q�Y�~�^���P�~���ܵ����Q��M\YM����t�|��ꘔ8_���onܨ�x[gFjKe����U�o�=����wxm��ce̟{v�*����R�h��p^D�Om��t߷?�NCO��)~��$d�i��/oi��6�="��;�:����3ڐM����phN�2��
�]g���L��bPw�'5*R1�H��EM6�o���� =��+�����)_Z��׹-}�X��:�(�|�\ߤĦ7�I�D����-�[��r	$��'�(�]��$�&�w�i<���ta"��:Ba/�Ds1�wd'�
Mg� �a}�A�Rw���S�S�̃a!V�\�Y9�8�1ڤP�����&ȭ��0m���OO��<�<te�����ѿ���=��)>��٪�ڱ�h�%�w3d�kA_T@�D��|2���f�g�%J�k��uq����`��=�ٯU�'q�z�qқX�jGk.��œ^�@!D��i����6<�r�����V�u�.�i9^���=A-&�bSַ��B��\�㜐{�Yg���0��ݫ� ���2�FL�S�1�$'L��������!mPq�g�ުz��"0�xz�hB2��DQ�dk���5M{K�x�%���G]�c�fG������A�(�A���d�Jz@��+��E��V���uc��r8\�T�
]�}��*������e���� x@��;X����9�a�*i�V��H�� �C�;�SP�b�"{�-�@0�wޙ��IM�����:��T���(���`*������Z*:ǭ���*��7���p��^�u`��l˒E2�Hj�_����i����rچ�@?|W�l����J &!@ ��Sˍ�#�2�/}�����C\"Mu���{����&|� �X3�#�����%��`�GBd�j�ʈcK��:�.,ĖJƪ�N�Ť�l����`?�\�p���~^��FҋA�Y���U*��8�a�.�B�%���he��i(&Ӳ�ɳ
̡�c�� W���D�T��Tm��Z58�3���x.�gH��]�����j����Uj���;9�ƍX�\��/O@&�%��@.���NAYY�`n|Y>��|����i�!�a��� rF ����9�A��GM���d�H�$�T��O�5�A�:sL@�0�nѶ+T`�j?NKb?�*^���I;5�������G{T	.n���_h��qlY�'�;��Rv�v��X�����u����FW�
ɪB��/rB���@�d�[�M%`�=�%ԯ��Vw؍u�e��S=\��x��K4ɖ������#������[�rF�y%�'�~�
h�����`UL_]����E���r0�>�^4n�������Ee�3�{���Y�x��Z���\�띅�&��09��{U�{f<�F�1]�*_�������6͏i7]���nX&�M���J�x�(��>1��×��X��D���|����T��O����gU`����O�\S�-���"��Iwdei�R]Q���jW=����}&Y�j�r����9��/�į8���3�Acژ��V `jz}�V{΅�b%����1��R8m��ƞ���
]36u٢3D%-S�=aXcsuE ,8��� �i�)��+��֡�����0�a�彝�hh�
�=�����p���aH2{��,~e|�8tO"6�,e5�i�x
3�؈5�v����L�t�V]"˶��v�x�B�	.0��
��:�<Hu'9 c2��v��y���b+o�T���QO���q�M1��*Op�K4���v��Zn�?Y먙�0�@���EJ�J������ݛ�ǡ�N!��w�<�;+)�|��dЋ4�b���)$>$�? D���v��|��7�I�)h`�̳K��d�|s�ا<�V�.������o�E��mx沌�rO`��6����x���G������5]\6�_guF4<�[�h��g���Mq��3KG~-ʼP��D��Q��x�J[O+Ҫt!�����o/����\&���1{2j����u �:z-�s�@���p_�*8a���6�E0_�L����I#9h!�G��x���tgoE:"
���tN�OB�!�+����2�GR�ɠk��DR�.�[7�5}L�N+Vm_��s�՚D��1gs���V�t=m'	��ʴ�z�T��/�(�h4HJ����H���TCO �7~�]+}�޿��!��&��P!����J18�j��-�5�5@
��`�+b�I_E.���X��:��m�0c�m�H�ϯ��	vq(����x�\� ����e	9(�'��닜�پ�����;�F���6����Zm�	������̼z��Lg&>#������uv���n}��#����o���{F�N��nw��m��;8na������Y�;��X��V�-�||lX��v�g<x!ĒѠ�l�f��7�m�Ƈm�_�2P\��`��[+���\ǁ���dOፅ��aȒ4�9�]��|���
�y���qW�+����B&W�K��gU�����/^�;�}H(���b�(~�����R�[ň�y��Y��d6���	INC��;�c�����q�JܶhR�k��"hM!�P����ehտ�V��:�x0�"�/��M���Wq�6��Ȗ?��^�
N?*{�0�W���g�?y��d��πVʖj;N��+�v\�Z����d��pB^��"��p�qǘ��s�޿�����y�fp�`d7��/2����NkeEl�R�~[�M{u��W�a���U�E���X:yz����o3�&�AK��(aje)"��h�y��O��0��m8iq]��V��[�a@3=o6��k{�e@Vg5���"4�l	��WL�m��ʄc�� (|[(l�K�p'V��Dkܨ�j6g�R]�X	�n��8y�'\��W�j��#BS	b����H�g��7���q�r6�9�QpE�1}�h-��c��X.4Ћ.VcK��k` � 6��Q:+�6�|�	�=(� CM�{7A��޸ؑ����W+gʯ�U�s���LP���m'@�e���M�ԟh��s�l�t]�6��:n����<�A�(�����}�������\�kq��&�g�G�`n�@��b��iYn�/�,|��2#��>��Ga]�#%�����/N�C��]|NG�=l����P.����Sv[�`穫�d�w��`��/�8bm/ˌ�s<�b���;�:�Uc��.9��y4�W�L[�h��\���.l��UkU�&Q��8��8U�H���ۊ@�K������ »A��y���M��~ �+�+�M%pC������iɾ�$��>�TR#�7UY�Y�:U�B��X��(a����z���/r�-@�K����Af�}V�����c~s~���g����	�nj˧���2pAW��BZ|�'�ig�g�Q�4����5h���YT����q(��щ �kQw`���(��>S����M��������B�μԵ�}������(9��W��ӓy�R:�H��#�;K(-�J_�n�L�]T`�!��yT��*{�����b�)t��f��n�[`v��
��!S�Բ�[�C��Z����VY="#v0������kM �zE��to����pa�����*� [���5"id�+ �M�.�$ qY�Rh������Ş��� !�ѬVa��ύū&En�#Gµ㮌�=����L�Q�Θ��>'�-?��e�o�r�.+��Pv=�%je����8�܃se
�/u;vU���S���X��}{!v.7=��A�?N��U�Ήr|d�c�ÿ��� q�S_h?��=��dA���%��_�ghT�LV[���lOkj�x�������>�gS�Ll>�9ݡ��J&xO/�T[MK��zύi�}-�F6�c��_� ��:�bT/�x��[ybB�wsE�HH ��
�;@NY�X�SM��7�'���*q��s _�r5"�,��6�?y��FB����u������u�~�>n5Z���Nc%��u�4�֫b\u�4��&��6�c�g�
��?s͊�U.3N��rnob|%~:� ��������!���b&Ó���t���c#�"��������ڽ���Q�LA� �p���p���> �#�E�oyc��&���˩�q�
Ku;U/8��vZ�d��ςUϚ5�XFH#9�Ort�</�������`%��J7�we����W��b4zp8:����u�R��P�(�y�0$E3(0�OA�%��}�J�c�	�[Jgg"'��&�8��3ρ���#�\��&��&lم��_y����@J�vL>�+�ox�)g�Sa�Z���uwe<�ۃ�F�D�Ǝ'�J�����Y�p�PL�Oܙ��Q~��ɬG�]�:%!�Nx_z�*�3'`��(VL�v���ru_'��cAxW�e��$�7}Z[��i��sH6|0��[sǏ�?��^i��G�%'j���*`��Т�ofa�j3>�hBZ�<�\�J]}Ϗl��=p?�hV�b�\9h��l�Ec<���� �:;�8<�]Aw�%�8������׮`�.�
z�
X���~3��,}�Ըߐ��)���K�id,��%E��E�^��N�������S��BC�FeWe��>���5/���A���?��\�k� 5��Pl��u)y��K�up�%��4j��/V�������9���#]E�J�����v��Q�dM)G��<� ��yd��-�F0�.#j&ϑwY>�C��m�񿷵�t��LNH�T���#r�Ta'Ӥ*���L���z��@���5+��B����E��{;[dh?�J)��<�9�	�VA�l�4z�2�Fq-���J%wjG��x�B�h�dU5��a�I7Ͽf���f��?e�W|�Tr�+�)��d�)YF�_-+�򶜘��FW���:���p��E}��76Svto��������o�����8����1�R����ӑ�X��IlR�^N��i`�P��[t=S�l%0���[V��ލ��>f��QX��ҀzD�����f$;	c��1#�,TW�� R7vFl�s	~���W�*z跌���>qd�Bs5�#�w���IZF<�� �p�Цy	H>��)�S	D /�:x�����>�CyX������=���NCi��iM���Lo��˟��F1�LW�<Q��H��}q�^�o��Yx�}W*���j{	yO��|0$�����t����+	��$M�1���I�:��1 �I�۱�x��ϕ�d�ï�f1��te���WH��(�P+�_��+U9�.Ym�� �� �}����%��6�|� ���#�����K�O��Ek3@r�7��/�$k��v&�f��� ���E���,�A���c�ii��yu���x��g;���B�`�#����
����M�dk�V��kϡ�	ŧ0�����q��>�����=[ɂeL��&q���Y�P���ŝ�vTKh������/�d�d�(\�9��f5��S���9H�`�^}��tx��O�ʯj�H�L0��+�.E����g7T�&�l@}_�'��C��w�_|�Rp�=����ۧ2I*>��D�n<ĕqj���9l��A���(������L�B�D�{�Z�5�~dGSi�1��}|�p䮆<W��+}�������}��	�S�Z��'�H�4�|�� ȬF����*�����)�Q����~�]`e�\�)$�>������[�>�R��L8���� >�l��M���c�UBR8�1�Z�.*D/~��Ux j7�Z�ꍗ[N*x,��)= \r�bVT��)�%0�� -�ݧ�|���k*�.V�M�9]�U�V�uBP��C��C����@О�2� �F#5\���$�5����B0�F�.��ö���_JA�"]�y�!�R\�]zmb���ǐ�΋ɱ��~��F"7]��/8��;�>aP��Nҟ��ȇ�<l�����Z�]q�,�P�>\ Y�N����攞/+�$VS�BA.�5]MTo�.�s	>"a3¤
� ��d��No�?�_Bl=1�T����.}p�S�'X��3��DRl�+�k#Y�T!Gs��������p¶v���vk^-T;yzY}�HM��SR��~���������y)K�E��uMyi���#�QC#I�X!���b�ձ�6�J�U�*!���H���9��	q��C:&������e�8]T3n���=S�i-$Uy"oI�s�۬'����G�飑�B�!=l=�8"#��,�8@"r��,�Gmr�<�3�{������ֲ�ܟ�e����wm�rA�g�r��+aCe�!��?P��ۺ8�{�5`x<2��X�w�n��4�4�!�<ӏc9�������w����gysr?e������]W��.Ŧ#��T�		o-�M}8��|1����Q�ӨT��z�j=S��3��>3g�����?"�5�#g8�#�.��qX�~�N�hG�3,b��DR��`r1�������ɃE̷�m仇�l� @�*=A[{�e8~Q����1�K��§�o�X�@A����ƚ�ƽ�`�f�����IOG,�c-��i�u���WP43�9r�������X���[9��˩&��E���% ��ǍeS��,Z(B+�l�Aq�B�6@�����c�Ô�B��PJXN��l������"w�|��ΗB�5Oc��1��=���g7R��{��a���X�,���
f2�=s���К���z�?�j������~�<{PDQ�'�b�F�
���%i�5@�!@���_	3"j�'����q@r)[�4�_��8�k^x{Sz4�JX���Ժy����R�w��JM�b� 6�1|!�X�!��SH�g������{�
e�d�8m��K;��F~�[��]Y�)[����R��	�(���ыT�IQ�,�N(�偭�D��pj��F�1f�n��&�$��lѤ��uL�*���ɮ2)�,��������x'J�(Q�z,q� ��� �T�fUW�}��~t䵃�b��7V�����%bqzX# 
�NB��m)j3�C87_��H��5�xe�xL^�aR��وL�F�����F2����}~��"y,�i���_��~B���@Ua�d����YJ�����1����B� B��%�hr�@���'�����v���%�b��-����Y�gwZ�M�g�7����ҨH����B����j�n�tD�6��$`(��D�g$䲃R	t]l|F!������#.�~}G�Uױ%��ͫ�1��+�Mi� �o�,�:n��3����/��z�9���3��7x�O1y?\j&L���XC����6p�5s���W]i\�{��LCn���Ә%�s�勹�� l�3�AԊ��
Wvjx�JJ�U�_�� �%î9�g,;�G�	�n����j�ɮ<�b#�c�:Q.�ۛ)f�BEy�0����hq�_T��6lG!l�j�{�� @�?����G����+� _�3T��ͯb�u	�Zm쑲�|t���r�Yւl�B1	P�$��߀,!ڣ�É=?;RK�Y,��VɶP~���f�1���F�Ga0wO,��8�iM�����ߢ��a?���+���ǆ:�FC�������,���.Yu/G�[ۚ �P��B�k�ʛ����h� H��b#��Ɗ��c�ډ�`\c���Ě�>�_�Jk��7�9�P�3�g:��U��;NYn��v0�^T�/_tw�2�uv�%C ���k{��ر�����ay��lpP����]��E_Z�l,NA�g��F����`b��L1d�Wa�_�,:zA���O	Ý흰bn	C�#�?J��-Kj}Cj���J�D�|��®�.���}bXoe:�2z�%��>��tpQ.����׍�n����b�>���ҿ9R{u�03:�܅:��B|��{���G3\;�<�>��{��j�����k��~P������9��e�|7[�c����ĜW��[L6+Ԯ	��a��g�h�VP��O�����T_mv����z!C<57@
M�"%@�ý+�5��l����(J�"�j#B�lw�_���1�|��L��ܧ٧�t����L-�旽un�dV{
!/����6ݥ�rIuA� �7T�X�R�㦩�^Woe��Cb��jߢ�P�T'�A�TasDz�X򽗼��7��g6���1X �����2��]7mSU����4%�c·�{+�Yo��ܔT������|�(ia���1r�J�1"{ܴ��Ǌp��K�Z���ܟͤ��F�<[K�+b��@a�)P�[�����!�e�AtMKb"��
��#��N:����ke	�'-��o2Uvt�_�����\ê�-�	O��Y���Aۼ-�9�'�'���\�����"���T��Η]^Z�@����W�/q�^j���Xe^*{�eW�Tɹ5�կң�����0-���y1z6�c6nz��E��0���1G�\	[]�]�۾�]U�_�ؗ ,t��E&z!�a@cx�j��~"�p6�6�В�C���撴`H�oԳ���J�jű1`��Y�8�XL�� �aFL� F�_������j��ɓ�A�˫G�����wZ���!��J�F�PWbզ��"e����<�[�p�!�}o0��bےS0k���1z�:Mf:x�\O{��:��y����������[ѕ�?8W���ｉ�r�L�����'֥H�T��Qa�^�V���8<�wT]t��xmy 0���r ��B t���-O8��|��9�R�<�|u[�/��/#���[��YM��T��2���YVbU�ƍZ�ү�0J�~��
O�� �[`�a����R \���#. �zn���_b�U ֢wy?]m�}1#��>k�{�&�U<�'1����$}��k��= �]����L3����H�/JwA,f�PPO��|U��^g���>ϫ`t�T�m�pEt:V�����Ҭ?B�J�N��pW�\ʐ�c#&_r��=��Βc���3�/�^�M:#u0�l;���屬߳��ض2i˕7u����$8u� �F��A�5ph��֔�QЦ2�1�x�?HS�v��w�K���2����W�GFb��-^��5�x�x�d0�^�%i�L�e�y��w!{�[T�gB��U��͆.TEё�b#	co�Q^�c�����q' ��p%�pR{�l� o���+f�#F�=�h�����r��ay'���gI��ڐ0����BY�l�p��f��5^q8?o8�2̥�S������JK*�P�w��0|-2�x
8']y�	��vf����-�y|��OS�{r+j�,W+��om��ze)����j��앆w��=�}7+�^�ڡ�D�z�R.��I�%�_��iq�)��r�b��:X���rh�&9(��L�oL��ꊍn�u�Q1��D�O�e���bFr.P�5���&��l�����M|��5W���յbt��sG�{�^��e���i���Kw����kVQ��v������}�|X6ҡ��R��pk82�j<�[�
0��V�b�`43�-�k�ZL���w�i��p���2���)�����a��|bE��QFq�N�)E��<�PЕ�s�g�_��C��ێ��c�W�$$�g(�R(zJ��cS��uGP=XOr�.O8>ZN����Z�3mk�T}�ی�nq#��D����߮s�����-��Kp��ecsĠk�4ɫ�'�m���MȽ���B�%Ų2�z�&s�t�&�zP�/�rQ���#}VT�b{� ��%�l��o�>,�Lr̴��mSԣ%OX���_�VQ�2�U���/��V#��!��_b��U�.$nc�a̘іkξ�B�Q�g
�LޙG\,9�k�F�vP�y�L_�z�@c��D�T��s��������±W�Co��%�B:Y�#|��kZQ�	�T���eYx�ʇ��8"Ў��M��0ȋ�yN�3G�L��+�d�"n��2~�Zm�9&�ψ�%"���
x�8�����������_�g�L'Jj�!���y��[;�èUE�%�Π�k���1�Xaڑ3�����.��h�����1iiP��:�>k��\9�z������r�R|��� �P+BZxZ�#���s��^�,ԟFP��Q�Pj��{%z�h��p��f�|k�x��k�ߎ^ߑ������ݩZȭD	Ɋ�7�f�������GKG�t��ځ�Y�=@e8��#���B����0��c
�z���@�4�F�/�jZY���Z�2�������b���#۵�J�+mF�F��f��fi�����ҲT�ŷeGm&0G�v�<�4�P���9������4�0���DK�;���V/�b�G'Q���z�&�*�@��6M����B��B���|l����4t�<{bo���'n��
&�7�?o��6�wѳ���q�0�*�c>�B¦&���I�t�t�S�8�������5ou'��C&FG:˘>G�����ڪGCl�i-��W����E.:���-y.�]HH�.�`zhċ)���"�����Ւ'��xΘ&�@3��=x�!���^i���*����g��x�ٓ=a���
ݢ��ES�?R�+6Ꙗ1k�
ʊ#�3��+��$e�8_$�HR��Q�)H
��"�����n������ְ��:;g/�6N�wyq�Y��8���c���Xp���/#Ĺ�+�����鼕�w}LL���4a��J]ËZ��d�<ϤU�kI�'��w�9����g	{e�t`6d��"����jy�����E�Y:g���x�\{1Tc0��m�	����� bk��)x�U����y� �\��U��?�J>Fo5#d�6�.�M�lw���W��L�/z�K��E�����"S����C���Y�7�Y 
�p۔�'D��3�&�oa�č�5�O
8�)oz+�q±� h@�˗=b0���$2I�۔�o+
m}����c,O_6	�V�sP=P�?���7N3�$��Oj��jygc�$��!�j��:���En8�����E���޷c�m�64��yy1'8���ӝDln��#"���(#�
�,�RXv�����+���R��K*�uC��R�+��~�1�7[ �|i��,lQ�g��V�� �¹�@5S���>k ��ۯ�K	��ȯ���'�U2�R��A���֍r����T��	A���؊�1E�:M�̥��|�ŠU�'<^�'��d�Y�5�E��J�82���.����h�6h�����������[�Ey�����8�ڸq�u�n����<bw�0�k!`���_ '��mtW�y��U���0B�⃢�v��3O]`cOjrl�<�1ΐ�y��G�)���ڃ.0<*�\B���Qci�����!O�}��uS��P=5R�ǓғLk��{"��*��x�=�,���T�<#Le\h����ꨱq|�¹l{��W�͉{������ɓuU,t4'M�	b�����)�VW���sf[l����w��愓��R�Q�%^׽�no(
e�<�W WUq���T�N�1����(��j%T���Kc���⓹�nQ���*	gy4�u�^�?M��@���Іi��[�b4?xzMӺ����6��@Y�K?���D}��A}{�H�@��щ#be!Y�A>\)�}�V�g��gh��y�fC{�8j�X- ���b���ĂY�����_e������{ş99���������u��-���ˮ+�g�X���O6�gv�y���2f�}X�Eu�BM����5�R�����񦈼c�ݸU�Ok�zDlG�s�E�2�9A���4mkP$7��UǗC���Ü�҅n�'�T������a� �S��}m�gّ�K"�J	ݹ����N����aY��������Xb����<.�b�)z;�g<od�;�&/U!�s�A�Bߟ��$��G��Q�Y�%b1�1���CE���m&����}�r�8{����P��DRm�;b�<�I솛&��
K-f�*`�5$�r�s���v�uT���BԾ5�#uW7a��~��%�s4ʥd�9�[�@}?��㮿T-T'A�W�q�4���";;�ZL��,+ِ%
^Ro��'*�~�}E�k�~�;��0ݜë�����4H����F^�b*R���P�#��	�\,��\��V�4��׻�}N�F�?y�<���c5��Oұer�Ҭ6��:P����]��@�
��jʎ��{��]���K�tB|߼��]w�ig���6p1,>���d�T=�5��V\ ��b ���,L0`��sg��蓦f�����0^��>�Y&{SԨ���L 3 _�;�k�~�'�R��5��͸�}���Pܼ8��s�LN�!wp A���T'�
��#G��K5�p�Y#g1{*�z���<������!n[t�in�0q�c�䞼���u�j�f�WY:���:�]�ڿ����H���>` ��
*�I�BO�zI� ���$�Ç�H��Y�t�[;=��(�Ĳ�6��+)�X��(+.�q��9�^�M�D��M��~-_��JؘË]��)�x�������Ȏ�5�*W�1�I�qf��p���4V�0zM����P��S%��'�;1=pR���e��ㅆېu\���(]ȇ����#�y@�rV�~�a]�]���9[V|����G�"D3��:���Upk"���/�v�*��m�B�-"--�Ќݾ�ɢ���4�yʱ�����Q#�C/3gR�����Hw�;U��\��(�I��U�κ7���>��x�>ﺹ;p��n<rE�eC�_u����4ث�oW��a����IL�y�+��9�x�e6B�PK��jf<Q6,�6�7�룕�{�"�;a���J���;��t��F�^��2��f?�u��6=�v����a�R�!�짉ds�YT �J��-� ��m�o��҈I�Vt37�,�ֆ�.�3hJ�Mñgq����ˇ�[�Rө�$���Y���K�Ӗv�UƂ"��Z�yϲ�������=���p�o|D&M=Ï��6�/����i����V�T�u�#O���t��4�M�9����
F�$�dA�ޅ�Ylb(�l�{p�	�@��}�5 ��B�j�d�M�x	D��P��!�c���� ,E?f��d_`w�.�8�����Q})����_'��!8x�UƙB;�mߕ�? Rf�����C�u�E��!]��WA8P]�j��ol"˦w�S���K��K	�~�����KWL�����-W]�q�؇�����O,fj���q�=�*rD<��ol�ޛ�&��H�p�2��-M�)�Ar�e�K�6:���A�CGD��1v�A��� �`���%ru�u}Y?eh<��	k6q!	X%S�U��!����#�]`�RB}�1�
���7� �뚧��p� �؝�x�ͤ��j�w�I��@��L!I�n�=��F|��v�)��Ė<�tɜ��9��#;�ctܐʧ���i��S�z�+�j����R�)�Jj���3�-0`������_a[a����'Z;��z��GK�qJ�VC(u�d�Y�M���a�4��qc����:������+~sr��(v0=�-�I��]L2|��^�7s.��s)�r�Y��r���҃��ɖI��m?��^Ӡ,���,m*�/���k�n5ɟ	�:*4�}��쟃�9�ɭ��@���-��X�?F��u�H�>����V�:��G���fq{�
|�]�,k�ч�/�x'�Goo��j8��1�Rׁ��}	U1�;��� �CS��U^<�/5�����Ml����p�=�"�:�3�e=��H�8�7����Nտ5������n����q�_#����+#V�֕��l�iY�&S������~��=��TOZr�%7Vbd�ݒi0������H��9�� /�?���+B�X��k++Cɋty2Wr����?�4) ��\ͪ�gP�Q�ڜ�Ili���Oj`ۑL�K����a�r9��&vb<׻���7��{�����Ң̾�J�@ʞ)�1�E7K ������s�v7����3�����G�T%C�r��z3I�?7�P�����_���|�'NWzd~���M�l�ǎ�'4т8{N�-�؋��qk.jj�����h<=��?�6������@�Ďєd�
��i�S����o���T���:f�	�-fs����ke)Dr���s�/I4ݘ��L�(ן]��h��O�~�ѽ*J"�YN\yGM�_0�d��ͥ�l��F]("K�_iP
R��םe��s���S�,2��ԛW���7��	�k��4n��دi��c���J� �"鑅E�E�GcC�����Mi���9}V!�2�8�m\�n�o��*֣.u��F�Sh�3
32zdd5�]��ЗL���6��=�^�LJ�,*	հ`M�O�׃���Æ��#!�����o��]��f#|kx�(���q�&*x�%��ˆ�]}�U�xw��Kߕ��b��.�76�a��JR���� ��{���B*�6���	��n�s+���l��Q��-�����庙^���S�y�)�ZQuSt�ب�	����[^�H �+��&U�A��o��\�|7��ͬ�q K�� �)�?��O��m�*5�u5ơ�!^�����%���oC{�SV;��M��3��� ���X�i�<恏˘C~n�5��Gֳ����`�A��j���W��(5�0�S���d�+!]�4��#�+LY���h�g�H}����(��'P�dG�������{<;������:U�9��(���Kd77�1r�;1Q�|��hWg,"��d��WKIŔA�y��E�u�"M����4;�L�!�#H`ն:��Ir����Y�5��C�O��IΛ����ɫ�f�c�\�);-�,�;'�*' ��)5�i6h�D]Q���T�F�����3�o�������.�WBQ�L}�����'~���c������J��!�M
N������R�����ւ��\�m
1n��&B���ӈ�T��L��P�N���@o��l�5]�����}�[ץ97�/�
o��?�
�(��˔w�]�7��a���";�\N�L���>P��6"{�1if�"}�F�e�;�6�8J�j(��}(��"�hPH������҃�M�af�U�a��=�,uX�7����a|��E�����Rj!�H���N���X-H���"�_P8y����G�8�%+�1�У�e���B�cm#�]/��<=����&7�_�q�/�) ���^�b���Հ�1��ƶ	��,����*f>`�Q�\�iIDCA!�hY���yC�,�Wn��fr��N2�6���8@��뇔8�vB�?��˝�-�q�>WHe���`硄g�'���/��J����Z|��m�(e�����Tt|)�4c�>O*�T���רk�)�����*�-���T�#���m�@\�O|�!2��i��jQ ���P�*,��ظc=��T�C��=jY�?]:�'�u�W�g�ϻ�a��.d��nЈ�[o�<��Ϛ7��^�(�u�;]T�# �����w�_y�T>BB�a'{�HKDy������Z�����m�m��ƈ�����(#���z��qj�}��a1�e����{�)geG�l�i��Q�;��%���fL>��6J�X,¤[dV��de��2Z�Ĝ�E�mu�������=���H>�9(\g̇<zlT �J��BB�vˎ��e��?��RS����&2�F�lh��@�Xxri�؍s p��k���c6�o�}���	��p����l+�_����1�����
-�)�cs�JUOv�#dF���+�֚����X�@��� ��)�9�0���7^�i���T�֪7������K(l�+�
���^�;�M�m�VOX�tm#J�Y�Ty��Í��y	PU��"�����M�|�?_3�Ɖ�GeB�}K���&�|h0L\p�˚��"Դ�l+4�$^*�čT=:u'�	PM]mAF�\�%��&��IۭTB�A���7E��fO_�m���'j����Q��f�a]{�.��nਧ-��cs}!?���/eW�F��Ybk��j~�G��Tئ_0} 4��<xGk���wx�r�
KD@�x��Cğ�
����l��Լ���	>�&i�Y̺���1G�A]�H��7�4@[wE�W�}h�N�R&��j��t��Q�<�%Z���4M�8ꦡU+���C�4|YKQ��_�0Sjj�.[��WϦr�V_�;�{�O���݇�����\���!� $���Ou���L�ew}���(��²,0�T�0ET��D�ǆU#���.�֛��m�v�ŖNiμ*ս����J��c�k�����$h�ė};�D��z���H���������isGrnj�.L�䧋�(=(-O�t*>�?*�(�C�kSt�1���*��^NЪ�m~Vp�>�L�/L�)�������l���>�]�*I��j�uS��#���=dvs��+$W�_�%�T�Y��� U��t|��w��xo�
��V�;�
��ZNi�=H�_됌5�m(��	�6w%��xp�B��l�r�Ѡ@�dHn��_n�6T�k�S<}�q� �P�A�0PU-��C��#��ߗ�j��^�'�AJs�1��%�Yvӏ�������3�P_7�A�[ u#������ԋAϽ�H?J4��ȴ{��)�D����,@5s�ɔ�]�o������,����9C-t4T��S���Qt��WO\��w��w2��欍��*ߠц��&�{��"����ڜ���l������A�����q��q���0���U	���ռ��'؅�C�0��$��
�fCX�]��~t;�&��ZP�U4��>`�f�փt��L�?�ˌ�`oAc��Z��=n���<`�A��FJB����`�w2�!����V��!Uq�\R_ԄY׆�s�O��2g(��
���'��!nK�g�Z�;g��}��4WI3~�W��g�hI+�<C�3��R�>̢�I�d�$����c*5Ə���K$�@�ܻUv�Ҷ�U�����P�<���Q~j�J�B�MW���m�3z �E9��`U��^�{��캿M�)2�Y�b'ü�_�"뫱.Y<�
,"�s)����2�̙���������Խ__[Cܘ�ػQ�X��ċ�n��G�s��jA�?U�5(�/�L��h��t�;ro�M����=rN^@�/C�c�8�[qغ����� �h�jJ�j�j�]	�}pߔ�q��p��2�`}F�"<0~�����OT������vŞ�p�<���Uz-V��_����nJ�7Y[�ye;͂��|�C���sJI2*d?��4kȡ��P#���DL�.��X���҅�I�1��)��!aR���V�4L�i[,���yn!��՟��RSB�UR3���_��!8�WY�D������֝B?��3�2�I;���v���f��4�N�:X{�E�	{�@^j_E
�F˸�����g���ݾ��U�Mc�����1uP�E34��T����S��[Tڶ��	-���նސh�oޟ��LZ=~�*SA���n��r�����/�|6�O����Y�tK��.7�br�JtS�pg�毇wC�j ���"���ۼ��1��Cu �D������4j2�o�H��[��h@YYDU�7%�s-nt���������m-��k���=(7���8^�7K�d���W�Ti�E��n/�s9���-�O�oM���Ŧd�k`S�>��=d�"<�:����g�(RE����ڣ��67�I �̼R�7u���i�� ����9�r�K+�^)9`��g.�m����6��Ƹ�Uշq�ax��N=b�ʤ�l�R������7�3�m���j�Nl��:bg8�N�	 ��0;��p���Sj���������ˊ0�'ϨCT��{�b�P���{L����i�c�9�̈́tL�1�D�!^w_�ls.s�f� �.T�d���P�@�+#ʪ�a���cG8���S]��<����!]�phn6�O�K�"͝!���^K������;��xJ��>ZK�-�q!Lx���$vaX��VS� �i��� ~-Xgzm�/� ������<�̻���?R��d����oA@~�
��(rM1���E�+?���tg�I�-��7��xg���T���T�᤬������b�j)<'D^�ΐ:�y����Ւ��������B���x-%��$G�yDrP0p�J��Ӻ@���P�	��TKi���4w�	��� #�L��n����GxȚ-�/���I�!�-�}��T^��*nv�����)�s0���0�j[�v���Nz������F�c:��k��(`x��ŷ�%����l\[�vmPٱ�"��/D�T@�W���8�"c�:��m˴@��ɞri	a�P⃯��C���{j�fF�����1&���L�Ք7Ex�\l��W��Yx�����|��a�.�����9UR�����i=1@���V�Zc�&3�9r��.�>~2Cu-]�t����o���[��I��D=�y�����$Y�F��H��)囕�6^ɶk27$�GB�Ɇ�C�*�V�:�>�u���X )Uq��'��F���g�������FG�!��C��V�&�܌;��:���Z�L�$�]k�"�������	=���ƭgq�ei�A��m�C�y��%�ݟM����u~�ڂ$�{��,�6��&�r�W�w�I�q��*V�-B�iYʩ�e�Ĺ�A����G��ˁ]��*o\;�
2���W+B8ӎ���-vd���C��X"$�e2�����ꧧ�T�*C�o0*����X+�~�ի6p]�l&�r5�7%+�P����:Gԋ!������ɷ��#�ƿ'�^dRܰs�Aeǚ?M��o��%ʕ40���r?��5w�/�#���C�� _Wi��m�璑�F@���7��3u�N�p����`~�$�CZ��J�х��3|={p�fp11�ғ��S64�q�_��*��<�8�l�����O:�Kԧ�.m1&�KU圫����=*�5��C��/�s�S8N[�J|A�O�V0��wr���[�H}��Z0m];�������K"K���|;:ı�A�TV����Jc�я-�Q���f�m����z��Q��yg��Etz>����O|?��B8���Y�(��U	g�p��Ű�.�`OP=��閲�,Ut��ڇAijR�U�D�w?�|��Q��L�6�Q8�ћ����KJAc(�RJ��M��s#����b4�M �M3D�ч�|ji�e��P:�2����X�׭�GJ6�����n��4�A��ҶJ��yO�-/A�ֲ��U*�o:�]e(ic��:�g���\O����$��b�J�jԌK?s��̼�g�A��M�S��R�+�-���a���c�n�xXY�U�r.Y�Mm��ƅ%��<�������f�N��!x)�^����ɼ��5�51� j��jV�u"Q@�.fy%�Ρ��a��+g�E58��8A�/^[5r��7� �K���z�f�ܖ�G����b�ݥK)�D�i���,?a=	�5��1J��4�E�r��.���P�4:����Jf�`����GG��Gʾ�������1s�fL�*$�\�^%Gĺ�y���50����l�"�N�A<s+8W�$`�o��y�VԄ����L��&��C߀����O�x��F����F��M���o��2=G��7�_E͑d$ŏ�H�m{�Gn��~˾�V��%�r��rk|l=VB�F���I�=ո��VoX:�9�|&�6�3�3�9u^)�H�5��w�Ps��I��8T�	�A�q����!���"7UU� �o��QH���ǣis��K!8���Rw���	4X�铌��9�������"�q"����m�9���>�\���I%��3����I��i&�B��r8V�fpQ7�Bb�Y`��ǯ�ۦټ�9Kl\�(�	bآ���,��*�Ō�J���ϙ�_�q���{<�K������6� v1r?�����Ӱ��e���
�j�����yS����&m�{;<�������V.�>��:��ϛ�M��::1��{����!��� dSh���k��&��(Ɖ�
�]:!��墜�VU�)�v\`��3�2�mZO��� ):��VG:-���5d�yN{���Q{��k��B_}������\D2y&��FzaL�L��|E�L5ј�hC��������5��_aj+��w?�rU��� �V<iU�.{��( hWD�h6����%�&f-G'�r ԰nVy�Yl���}���r��������	�C!��Rw�	!���H���G�k�	I���I�Tؠ�`��������N�����3ޥ����l�s�, ZX7N�FV�p^�I�<[E�w�HB��]C!�o�^����<����:!-�K�N�-{���u�~=y���U5`�����2E�3����!��p细�f�⻂��#���v�{YZ;�!E�IkF�n<����h����y��=:�iN�NUE�VV�O@]Ry�,2O�Wޡv�mո�%1ԭ�" ��B���y�2���yu��ueJ����??�m8����fsȄM�j�v�}��N��۳G�&?��i� �R�H�W+nX��av�xqfX:�a�����ȗ%�߹����td�Ϊr�wOQ7�Â �#�p}�	��=g�IM7�ט4Ѝ|T^v���P<3$/�f�k5^X�"��w�Z��Lں�?��U?@�
D�4s���)�)��m��=ӛ_ �t��Yvl���/TX���.�D-;���=}R�gGw�YQ�E,�0�C�E�`n��OC��eII ���j:2|��}�U&�i�zJ�y��c)�i��>���=V�D�R4�'�
��4�
��H`)gָ��(N��ҧ�(�X6��)�K�`�vڜ,�s(ge��'��;���=���r�C���T)����0�HL�k������d��9b��,/�.��ng[���8b���5.�DL�{���Ǐ��̗;�l��3��$V̚4'-��(V�Dġ����[�2$�n��U�p'��$��!����6��m�v=3@�5G3�k�i��I�9�~s��P5}���lv�
���s�q���c� � .I63@^���:} T���%i2[��˘	yX��\��l}�L���]�T��ȱ��"a����h����V�9�M� �BkRJ��.�̀/mEs��#�n�*��7{�̱vIP3��/ ˕1۾v}1��F]U%�m.2<��&��h���\V���5��8�؊���>
X�q|a<�;߮�W��X�k�|h��Y�r�dߙ�9y��K�WT��~� ��۠�Uğ_+�h ����WfmB�?��O�@��b?��t�LCEj��k^ȶ0�(�~x����h���Ov���~cm��R���wߩ��Q��~^x����fшe���"R���J�OZ%au�c>��'i4(�?R�
[W�Po@�Wt�*fS�Gce�es���`މ
-�l�q����U�ˠ�tt�n�$��TՀ �BD$0���z����C��%{�X� ܞc�����?@�z*:�w>w����`�+R��F5لQ�o�����W���<U.H������B6�Gϯ'Ek�x��>g)�["%�0��b�0�k�jA�1�?�P�_N�Fl�W!�/Uh��<���v�,t�4�œE{��ٛ������h�V�i��¾	��H�� Akn�E;���������\y�=����*mU�%0w��|�ERq��U���[�f��}}�����V1��J�X�9��g�Z)h�ShYo��3و+���3O�oU��aT��P�>c,�Ց�'�Þ���fyjG�<�htp���-����D�:q#��q9(V���B�t<��H4��xU:9�ɔ�JhR����vK�Ɂa��N,�^���4}��7?�Cf|Uہ<����b��Cw�K �>z8Qh����|yԩ-�V���(q�Ɖ9��X<%�keD�G6Y�(��e]F���q$֔Bߡt�!�8ʙ�>��+�QyR(� 20o;�p`_���i�Jzr�+9�F��de��
�؏[���������{e��K���'
��-� �%^��G��_��?��cz�k�^%Ш�5G�<�����:=F�������{��R��ɻ$t|]��P����:^PR+�V�X>�,�ŌAJ�1hU��	y(%`e�nU��v@�Ҧ(�ܼ��CflH=6]����/�$�QO�����V!R�������[&�{�Jh�Ƥ�LE�Phw��������7��qyGn��
��'�k	qְ���v�@�`i�?"��6Pu<Q2ȴ(�͝ws�3��`�<��"�p��9`��:����C��Xت4`�I�M(�Hвe.�l�۪����o����z����S�rz��a�f����1;��𜱨�c��dԖ�r�U���[œ�K�=��k��9��%p�E݀hr�%S�Ѵ���^�0~a�`CX�ԃV�/Ren��I%3�7�e����<7(j��3~p.��$T$�5�X�������@��	oa1-�o��?�y2�v�(�^�%�ַ���`��~z����PJ��E��9|���7�m��BF�/��َ����3`?9�ͽ�ȨQ΂��XS�� ������"�[�i��O�$M�"L�5�� %�Q���W9�ݻ~v�wr� f���8ۑ�Ҁ�;x����L��r��n��u(�K�B���������|�>Z�(����O����)T�+f���:6q'�����AϾ~d4�X70O�^���WR/-w5�^Tn������k\M��,PI��w����y������˪.hp4Vd}(N ���:e�v�'mQO,~�b�����?@����34����qĤ�Zy|�<U6�09�DmF1���B;N�5	 �A뙍&�A '�hs9aT���B ��]�����n?)��v�c'��@��}����8L���]Oi��Ŷ�]�4Eh�Ɲ6e�#PF���̷]u������?��|E�6�X>j��?�
�{)�8+��4���-�kղ���\a�/}����&����.�CU$D;��S38H]w�8{{����6vU���ع?�TsTȽZ��䂗U�&/�I�0�Z@���+ F?�h���%j6��Ta�L�ʽb�d4�[K~���d��7nw�W1nW����)��16
�K��qi�k���5�v�e������:�q��#���Uu �RC@)�P�3��c�h�:�XA�8���2�I�7Xb�?�Ҳ�5Jg�����T�-Ȥ�<m�B�9�ǽ>���-���g����|����iG8$���z���y���b�L1ӎJT�|���:����(9l�p��"�	���Y�����H'���ZuYϫ�@K<���
P/�
>�Urh��?NKb/# �v(���x�L��c8z����n�G=\����C��E�0�Ix/V�i���c�����)o�&��z�48i9�bE5��z�b��,��' ��n���dR���V3�ԏU�u�V�_��A�e���PA` �ʒEoC���(l|�x���#��\����}��B2܊C]n	'A�����É���s�3�e�����L�i�� �:P��V�uڅ�� �����hc0{)[t e.�iJ����:�˾���V�
(%�#K/��qek�0������ �'�/#OaSe�.M��W���A�[N������F}�����JɊ,D�5�
��p���^%��W�C�ݛ���	p�N-�)
�X;ʦbSu����K��i��J�v{�o�7ͬ�v��EL��?��_���PJ%̋��j�xf��%j�#�Y$�񻮛��Z�V�Lkh��:��j��>r�(�/k���R�Dg���.괠�? �}�?�S������u��7$���4��B�p�DZ�{���.v�$b�8�%W�t2lR��X�F0��TT�8L��wT�	�L'��Y~vi�e����#�<2[�+�����`��z��G��yMD���0�l	9u��I������|'��fʢ�H��\�X��\*�a�_�󪝧T�'+�R.#��:p^�{jCl��{�"8z�z1{�
�w���,s1����8"jXK¹��9����%2�)�4Z2[A�74���e�[����Y��tJe�\��.�t���_�j���41ѹ`m崉��2��ߐ7��s
}sm����˥iГ�c{��wW��/��]� ���z���˵��`R��_|����>j�a��7����8+��n)�>���4CWL��;��l�Ve����YC(��3��WI�j�L�ٹXECS�C�5r�%OG���%&&�>:��$����޵���&����sҁmi� �����Vyf�����h��=��#b,����4ޘKk ��ǣ��1�9T������Ǵ����)�����,�������F.!�����}G;�Q�v����d=x��?�Ā�n,:5�",Կ
���j����8S5�8ݔ�w��/Y�pVy�'|���E����2h:kZ_ODlA�pCTV"2v4$�*�����k6��yE��i���ҭ�"y��Gb�J�wݜ��sK+:�*�a�����8fL��Dac���o�g�����{��~f��1c��ӯ�����3Ry���AE�uk�+��ӢMN�p�LOs��=0A�@`��SƁ,�D;���ViSE%t�(Bt�,Y��p���Л2�pC��<��X%�`��P��4�V�f፽�YVA~�����%"u����.]�����/���u�����[9�Uq=�GJTޓ�VB"7|������y��S��nX�z��?��G��a��!_kĎ��&��ᤰ�t6u���ЮO>bv�V�Y²�P��o�w�3{
0�����mb��S��
vl�g}����?E����p\K��>�����m���Zݝ�e�pmN2Q7��fp�8��16�`^��;rM�y�w�$��>I����_�7���nH���ץ�o�^�3�@S���Iht�[���i��~/R�Ɉ+�l�i3�ԝ����	�j�3�Bd��4�@����v��7���gqi1#��A�E�r���pd�%,�
�}���NJC[_>���{�"�U�iplg�J�U m�֩�-'�ˠO/��Ϟ��C���)�t��w�;ɏ��O.�pvSiHxa{���%�go���)���djB�3���|hm��`��?ڴ�9�`^���{�XE��W���v��yI s�T�O�?������/"�ߵ�7�.9��Z^h;�4��̯�n�P�l�hٶrcȳi��3�#�������c�d��IR��8����0\!�W���K�V
�{\TBO &�<lPY�Y�!/3� ͼ��%�E�=jS�Q����ϥ�$�폍�1�"1��%n#����A��V��'�����17� K��@�)=)4���x�ԕ�|V��=.V���X�^����(È��{�9�ȋ��"W��,� %т��."+_6X�h�$���i��nq��5�<�����
1���գ���R��!�H�y� 2��ʎ`�2h������"?���c{�ؿ#;�����贒�'k�z����¾Y6������s1�>Fܩ��(RӘ{���"�0�+�""��GE�۰��T�r�|�sĐɸ��"-��m%�Ơ4�k�/�ɱ�~��'d��%ch<�1d
��:�o[���|�rj9ŀ .4$�9h�SsC�أX�%va��?M�pwyF!y2�wtGx 4]�p��,�$��Wv��� �'�ל{4��hL��tL����Z+�f��fa�6���Ї� �!��5�UƤ����^��#iSn�.u���d�]j�������Ў�J��P�GF:v����C�L��z�.�8S�hп(PRm�� �Fҹ� 4t|�H���b?gT���۾�=����4D��e=(Izo�ޙ������?T��o_-1���+�%j��G��+���x�SJ-�� ]������+�0�W^F�����c�?1F�&K�`������}�߾N�i,�;O�C[��M$�D�ưM�)� �<�m�X�DY�ޫt�<�06>Px4q�]���4rf�2DD;����TabU~����f�yT�E�I��#��#S�7KQ�[�@�mGR�)�sK-s�\��\Ii��؇��St�������w� H?Gg��W~��r���{>gN�U�i���8"ڨG� @���Z͸��2�*	X��-*�D
Q܆�﯊Y���������1��";L�|���3�@|���9;lbq�ϋ&�����.�=G� H_g|��@��08��b�3��^^z�O�S����8��B��i�0�5Q�>����������b��9��.��y��<�*HX�!%��>I�md���NiI�b�~�Yh"����Y����,Э�<�:��%x�&���h�ofC��(]���HK�SYL�B��iW�,�މ�~�p��� 2� �k�����d�G����3�\M�q�̗��U��^��,"��W��5�$j5�x+Ϋ�(�^]"�iIW��Ni�j��E�o��^!����3�\�=�u��
[L��z��v�c�I����ڠ�h#VZ���������ԇ��,ۮ�d{�t5A¢�魓�DNX��g�ӦE������YՅ���W�It���y�z��q��l���u�Ղ���Be�І�ЦK>��G�M� ��xغ�d�i�����	{»���Y:��aKd8��"-���g2f��. ͻ>��"����������Fn�jʹ�t-���\�mE�mؐ'3�50����OÓ$���|^�ګW�~�DGz�T��E��(�4�g�p���uk���m�ɩfb$;��y���d��s��B�a�X��&"�����ӃrM��#mK��B'N�h�i&+&��(�������3�ੰPyRj��k!�ӟC&�ņ��-��Fw��1*�T���O����[d�3�<�8^L~�2<~h�,�C�6=�6+�S-k�D�W����mB�z��7�N�vsV�`�ψސ���Mly�Y�yT=IlW��Qt�H�1�!$.<$�fZ޸꩛�b��
S7t%m^�%_\�|p�DN�A6�ou\��G����>�{�E���tYB_��S���r��@�����D���ǥp5W�5X��֓"�Sʔ������Z��_ߠT5�K��\�Q�����5`�|��U���-&����cԕ����u�Y���!�y$�<�����Л1�`oqv�vO�R>�:d`�c�K�M�9���5 �cz��=�W%���eZ�_���I�{c�&D���޽���+Hm��9���R�繿XeL�Y��.���c@:%��	�������!t[�Z�����і8���2���Ȁ�W,Q@Bhr��><�5�S�U[�x%�y^Bڔ:����]y	���!UA�wA�f��eU̱H/x+Q ��} L����S|���Է�/��j�l� �c��Hւb�X��EQB�V�T.<�Y�9����cì^HѩF�=�ȰL��ϱE]5�W�+R���٨�p�ʳ2l�
�U�UcbPzf+�ճ��Q��+����>�A��Cpa���q�J
�q( 4��VL.� ����F̯����Ч�(��-x���6gR]O�L����, �T��� mÚYp��v,$�}ʸ�J�0a�䘞�|E��8V���eǀ��s�K�oE�U/:?��r�d��z#���lP����վ�Ї���P�o�?�$O%4
�t�Fn\�,%�Sz�w�N�
��N�M��~�ya���%�w�'s#jpzaD�iazC�z��_���D7�Jy��ɶ1�Ë{��j�&q�W�b�-�v�V� ��m�
۵��HbZ6��@�sh��ű�l�L�{[Svh# �i��g��!G��#�6t���x�������=s3�>��@&�d�!�B(|˃.Ѝ��%-�i)��!%`8��'��K�*�)Į��A����]����d�{7D�=�^+�5�4��Þ�d	�j�d����.�*/+�%k�6?E`\��(wGBqJUU:fָ�̓�=c6;r$�J���r�Ԭ�����˨�R/n��P�(�����\	;�v;�j��o �����g1z��aÐ���"'��`�:;���s-�g=x��p�5�:�X᧹'z��{��4�_G)���Z�ur�ݠ�gC�"Z66T��>��D5�˱�7 ���'�۪�b|���L�e��[����j����~ڒ݈)����������E�5��SF��@ ;��)~�˫莕��{�{+C��Lo�GA����c����0�Q�A�ԥ)l�2�����湥+�<�w�^�m��<���>��c����ǻ�W�An��b�y��x��J�Qu,�X���� XW��b��������%p�p�KQ��N
�D�CW�Bm�x�e8�^<���BJ�ӑ��+tJ�;��a�s
ӯh�����s�<ݾ��=��E��X���a�Q�%^9�v�Fy�����pZ�&]c��{*cl��w�'ſ�t�����@x���Q�K�mvTv����KM�7���g4��&�FUf����+_�$�����l�M%v��$��V�iv� ��M�H5���b������50�cNIlW�S,�����_�hDIS�7�̺RS9#���N'����B�KAw1��$;!!P�.�T0�����_��P�-]�Uz�J������k89o�xw��
�]Ҝ�<(#z3��ّ���t� �%�gU�x�KK��5Wv7��<u�2�_{I|�ؚ��m
ӿ�^�Q�<��ݸj���_���� -�1d�s�P �S��ѐ���[��:�plx��2�D�%9R3l����͟��H9����8��bqhz���s}�wfsH�]�ę/�҇P�""�X*S1@���7	Ei���T�1�S}�q�D��^D�^�J)���g�����F5LTE<>� }j�K���)�@cō��!Z�H9�TW� &N��UM������,b��12�1/WL�%8ƬŁ$t��Zf��¤$B�C�v�}��
�@��tj��/K:Y�m�"�q���o3�g�L}�J�4\�T5��ZHP؆�H@~g�ɻ�Ao�[�}
3T��	f'�kq�m�d+/&]���}����e`qqq�!"���S�&�γ���3����d�߈+�)N��|�e%�@#|E��Y�m����ꝙ	Be���#:]��e˙�k���B��=9����¹�'�q%�y��w�� �$y�W�6����v*��l�D��Y��b�7�T��p��wn���D*}�uβ����!�5��6�b��F7-�RsQ��Ǟ��y�i��J����)��߬�|d�;��W�'�,��C������L�k��&���UvMn��{��̽M'`F����*z�D�@~�%B|Q�"O���
�N�잃����|VM]�3���J�U09w�������v�<��T��vXi{;�	>9���a���k�Ѵ�eOh=-�����2OU�Ā��T:PJ�D!�?��|^}h��	��
v�.K%U����E�3y�x&<���Q��$�e��İI8����?!`�6.{76���-Wn.ǽ�x��S+���S���H/�T���ӑ�e����w%!��B������
��vL {'����D���P����Φ���i��s#V�r�b����@d�G�5(������c-��l����N]�_\����C��>�:�^b:~2m�U��������ު��2��pǮsc�lĈ3#�8�z��h>al��k�t$϶���?ys�����Z�`.6�'��c�N(�8�4TG_����~�~~�0��Ճ�z���A�`#�w �fg�6ri��td�\�<X>1�&��^��#��4���-h�I��y��؇h��[�o*�/9� 8�
��^=���J�foz\P�	XjD�7��=Q��P��tg˃Q:t�Q��
���u����$A�\�G��T
���nR;�>�� LwZ�tl��{�m�ĬFdT�P<����|�b�o�|A��>��ҦR=���H*<�r#�Bx��Z�}E^ϔ�\�/-�} ~1�^����rnuBӲ~�G:�����F�@��#Z6)!b�訑(���VSIz�E8���*��G��Z_*߯���u������ˏ_\,��+�2/�;��3p�.��6H5�di���:�<��
S��mʵ�z�l#��ٞ#!yu��p��|qT]t~�ߘ��Da�0Kkr���� U=��L��e�K�r��a���bC��mcS������k����:	&�d����dp�"?c]E��ptb����Tr����=�¢�7s�uXp)�Ys�BѨ9~�i ����8F]<�q�t�t+mNT������zM��ε ?���l�d_��UgG44�8�@�hn'�|fU��n�>ȫ�&�Ƙ��j�>G��{|���e&�Nt���g��r�AK�T�!k����H�H�oW�YTiƞ�=
���;'ZW{�A�jKI��h�`Tkfaz�1��瓢U�-C2��
f�lm��A&E���w��䚚K8���wg/2r(�'X��BہmNR@jY5��?�Ȓ�w��d=wF�uU���D���s~�Ǹ��^
Q��OL~sOH���$�2K�p^ܴ�;a��t���,k��Ni���!��s��>���z'���%M��Ae���8E��[�����TM�S���Pe%�%�_ou���+$��}ԉ�d�[��QE����E� ��~1i��"��~�4�t�v⯟y��� 9E�Aݙې����Q륾�v:)��0�)BrM�����8�IP����xօ��~H��?��UOQ�%�'x"��w�|���Ut��6�O���ࣽ����x��{w��0�`�������g�K3������1��d�f�G�g��*���s��m��)C����c�7p����@����ހ!$��}5���z��A�����E�lwvM��`K����xi_�S���z����F��K�ĭ0�r�t���fJ�o�ʜ�e�g��?F�N��5��z����
��L��m�?N�L�]C�V�����]�>�x��o�d@5���-u��%���4�����曇����v>^2T6(P�,hx�t��նM�:bz��'�����j�*�:��w�޲x)w�K.'q��`�5�i�#��z�Rf=Gi�l���b��{:��A�����t�$c�w0V ,��,�s�J�6	�.*���!f��T9ŊDa��w����k�����|�@]لa�Cʉ��"��r��ʠ�S �}���ejeu��6a�g��������ui���ݑѮEUj�\��F`~�C"��q���M'��$�Y��w�8�T�*�����X�n����^���2`m9�t���s8���S��ݡ�B��|ڀ��H.�2��-���
��9���7�H^�� Kok�=a�f��z[֝���Sk&�n�*NU3)���1I�;���&��{�;���M+�'����&�r��Н���}%��l�~�� v����=ן���������^ �c�~-���xzvf�뱟׼e)	2F���̖��ܒ�hw�4,��}H�Ⱦ�u�0�WY?*���-𭂩�1��в|�wi��w{�}!��wQ`��w�<Q��+��Z��������=A��93��
�s9���ayW7�e�����E��*���I\`�[K~es�K��OЅ!E�e�����,]8���g�Y,XJUքT8��V	�	�Yb����Ҏ� <;�g�Ks�j��3���)��7��
��ԄU5�����:,� x��Ix��������t��A��������k���p�xO�e|��[j-C��E�vS���(�X�af�홸�U~�b��~�rLV�{�uq�2ܕ��&����S��NVp�)���������{
���;J�[_D��v5��0\���N�K�6{!�M@=M����t�X5���6 �+~ t�(tgs��0A3k�v�[��#=�Q�\�őj�[���m&��D���!�ᄉ�������V�m�Bv�yt�� 2�߹'8YW�dd��kfV�WV��_��Z�o�H;�|��2�p�p��A�T�*�����x��4�wF��mIͭ�i�+��r�O�	и���:Ͱ�yg�K#��v�~@�h�)�%�\��]bخ�"[`~�}��[5/����(�¤����/Cؽ��]4���yRb�{;�yz����T��)9X�a��_m�A���9.�G�Rz�	�;�å�.9���07��-��yR� �R?үT}6�F��S (���4tb�9�;���6iRNi��E�T�1˙9<G�����$�9S�?y��S<�=����>� (��#R�`�
(� }mn@ЂA�S�ܱ%�*J�ܙy�>�0I���Eg�,��|2�.|Za�w����$�g�.�Ie���c�x�*�/���y�W7�O����ꡢB�#c6�S��:�3��*��6i��4P	��ɖ͠(�7��Fcg��2qfx$�|�Ļ�������˖��[U,\N�6PS�R8�HJכ u�g�D����n��Vs~/V���v0�A?D
y�v$
�UM�R.��5��5[�|��m�4�C�E:*r���9�Ht�H�>��DT�����i�L�?�aMtLK$�)wn���%��w��m�Mn��47� G���Sc�f��}�0�ȑ B�'��.$`>@ Rۄ9dG��x�y�������xy��Iz_V�߂И�X��=�:Z��|�ײk�*��bu�t٥�m������c��>]�G����"\�'��F��`�7>�Ծ�8�cN�����зt�ӟO�h7�����j#e��_�w�����i���3��6��.兲�i�����<� 4v� I�O���ȏl	BQ�O4��X�!I��Cι���&y�9����*&T�l�D^)��鱛q$���m?��Q���T������ɕ��5v�׎�{Nƥ�wK��I	�=erY��(��z�[��$��񆗠�w��gd"�Z���n�6�S�!���ap���"�?XطI�j�զ!z��HaN���(�I#c��tӟ;������9�WZ�34����[�Կ
�O�+َa�,��
�c�0\��"�'[#1^@k��r�@�^�1��W��������
ဧٯZ���I���#6iWtߴ?\��I*?<q�k�[A
xaAy����F�+�h��,�.��������z�\Ќ,�&�ҟD���i�Q���*x�V�����Ee2�O��+X�$uj/��D=�&J���.{6b�]���x��������θx�������� 	A*�+_��J��"Q`�t����j���U%�����m���O�q��v�#/e�	��2qw��A����ه����@��L	ժH��-�
)�#�*r �:y7�դbb�n/�2�����u��PÖn�S���' �����(Ը�o��K��+��_f����H�na��;TC�F'i�a|��f�TF4yR���w�
+�_RKL~y̺�60��xy�!�ɤ�����U��aK�u�xw�(�ܖA���Y����w�U7��͜+␅�2�r�]�l `q�� ��X�-k�L��B	R�`����Pq��"z,��%�[ ��6�6��Z���������c!�;�ϝ+[ը ̼\�\)8�7�Q�K�!�R�BHwsDi�SԦw�j�$rQ��7��*�	"�%&�V����:�6ԙ�_�?"����g�yu�-$����g�:%S�g3��z��!/��e�J�ǝ����wL-��Bn�ҍ|vl�@�itE8cޒ�:����q�#�����Ϡ|�	��-K�0��Ӷ˲>|�*��o3������F ��:�į�q���+oA]�%[>2�A���O�!��s�&�L�����p��0�A~ش�A������&�ܲk�إ�)�f��|��}I�̱��*
X���/�7�n͵���mz�	�_ ��S��%B,�`j�]$������j�od�,��͈��@"~�g9(���������7�m/^V�4��V�?���i�P�����?im\)�'$}�q	H�z]u��f+���4��[��c�%"ԏ��J 缺�S�jv��5�/����M�h��-Y�\1���e�\]����7z���U���e�=�il�ha������y~����
�`���F U�l�S&b�ؘ^z����;���@D�"@j����Ej'@�E�yX����@f^���K���aDV�����y�F�=U� �oϤ���{�xe!�Q7������=L%��^Ƕ���5��u�b��g��dGZ;�WK�l�
�ڲ7s���s]�(�5����-�x��]�ע���N^�j�q�(
`Z��)�N��Fе�����X�������0R�D��:�3����l���+'ʫMV�ŧ�K�T=^ߞ7���*���0&i�)z$�Yv�XSm*1W�1�� |Iq�T��!4��nK����0Hx����C��Y��/S.��=��w3��v4t³�޸z�%������N{���UV�r��q��4h��ⲇzi��Hި#�Rx��E�xl3f�*
�Q�{t��'M�V���C@�з6�����u���v������;K���4�y�xA{Ib�!
]��x_;�����gKB���\U!�տ`4���e/�����C'f������ڣ���#%%���S�n;���q+Y���Ӂ#��|������V;HIpyMl>�������b;O���F�j�Βŷ[�fptB��T��Al����La�:��1MLӶ�-�w�	���\��Q��ͣքw��[�8�Q3��p{�@"�X=V�p'Ic��x�Wú��[)L���*�Kv�X���/��۠M?����������֌�p�ܩYݦɳM`ϻ=��~��t����������1�]�s��8kgR{��~h�T��p���׸�4p.w��������x_��k72�=��̸�Y.��=������g���Zȗ�m������QRGo��_�!"�&����$w;Fx��=�L	%�p�RJ$MM�74��>~��~'�Q��Å!�����h�]P�57��"���VhOk+�q!'`V»n�tǃLu����x�w$����A�j��䋇���fq�q�J���.E���b@4,A�M�9AJ�*/\��yr�#�r����צ����5H� �F�(|P�`�h�,li�:HAwZA�'��(E�D��=�/�J��CŁř`�*D<*p�v�mj�gD>..*y�.�hO�!��߅Y��'��m�Z ��v��5�|W��]3�2��t۰�8K�W�|2��"�Ǚ�sB�a�BvJ�ٔekq����|X�-��6{�f{j�KJ�S��}T�32��x�ډoT!qQ��H����<ãL��i�'!��ŖC-����@�u}��i1N���Ks!�4��;&��ˇ��rR,�/fg��L��|�5���՗���Wn�mժ>�U:u���aò��X��#cQ��yvb�`��E��_q�<��w
�?���j���b«���<q�&�
{��ߏ�,3'��%Uc|���ɨ��<��p�-m�d��Qh^k��ԸX�'�֘A�+��� 4��۞ ,0�L��C�L˴2)�ks�O'/�|'=}[�*��T|i��l��_BDzί��L������2	@���.`ˀb�t��ʋl�Z�$fp�$%��a��A���|Aw�SWD�x�r9՗'�\�̋��`=~��*z�MrY���P�7�) ���Z9Y���hS�����U���Yɍ��\X���(�iT�)��vvݺz��Y�O�.$�Ї�td����W���0,��)���;�}��Ӹ_���ߩ���DL��}��{�+���ӹK��`A$�˖\�GhA�A�B��m��s�Ԍd؟�(%@�SAMz��S'�&*
���9�l����HK1A�Q�$z��*L[f�u���Wt�֠x��k�?�?������G'Xu*�*Qq:�0c��si,�LE(X��en'��j�sA�x%gV� p	��"cɺ�=�uz�)jr$J����^�d�-#+�G�:ƃ.z�Z�GcqE�L]ES;�<weY.'o��=r�}��h�-'B(:��WK�9F"� ����h��ܱ��59��S�(i/#������T���(�(��#����W5���H"=�+��2���1ȇ��}���z?z���Q���_$ ����?ɊM�U|��T�h4B�u�����s��ܐ;h��,���nf�+'J�ĥ����17�l�b�G��\�m��3B�5$��%��(<ҧ�5r�jB!���o;�������;�%
�43�n��:==���O�T����r�Fa�$�Vc�iAF���`I�J�#�?�}��5	�ÎIY��Ȧg[jbc;�pQ��B�����;*�݇6�=O٨���ݞ:�E@s3|�(΅tH���ț�Ԭ����R{���g~��J��	��4��Iͧ_�,4Dɯ����I��t�Ƿ�in�>l#M/���wទ�n��˪��0�o���8T���P������_��\�2���*U�StC�_�8I��W���Є@�ԝl���
HN25�]F�����q-������{z�=���cՉ��"
��f2I<�%|"��{LAQ�����,�qp� ���\Z�mY�����b�"���!?��4@���WAc��r1 l��	��o[�gf�D��R����ݖRk�c��%6%��L"�G�)i��* �4�X�E�{�\XE֨��?��F8�eص5t�
J�6�n1�Q���1� �Q�$��IYt3�$޿�F��#)V\�S�{6���7�Q�e(��n5� ����>���
 �Ɏ�ƧP��i��=�4����E��+ Pޣ�=����3�=ߢ���C_+�	�,u�W�	��d� �[��$F5��o=�1�o��J8I��!���@uiivqj���͔V"�5���M>-��&8�S����[�̪xKY�A5`#sqל"��s�����x�܎%��k�g�]��Ճʻ���>|���n̰~̱�7��S�#��G[*h\�7g`6	[#��U���=����c&�{xl���h+S���C8�£�3�=_�Bv�w�NLnI����e	A<����/�9=@�+�Z�{^���BVf๞�Zz���1Ǭ,�S��{�9PfZw�5S���5'h~��?�o>ʯ�R]�~���8�L�;�ʮDF�>�\���o����9n/�:��S�DshQW�"��h��-�Yo���Oa\8\��������k�2,3K9)�-��X�;���G��|z��.��eY��}�6p�w�������p'���M��y�/��<tS����!'��k�l�jթ҇v��x}	�S>�o�����c�w:��P��BX�	e�	���S����K �Y_�[!��{���[��ԋ(�����yԩ�W��C� }���ioc|֣0f�I�RK�A1EEy1p���_�fvo��<�'�wq�Gx���������ׄ�Q���+A~٤D���Ok:��=��؃���^�N7F1�����|C�ݙa���oL�<�R3���RL9@{���I�[���Ftru����O^̍���򨖍�Wo7�J�aau��AӸaQ;�I�a�Mj Q�w�&eJ~u���-��3[[�I>Ybo�x�$��}6������Ǿ����u
��ߋ����Y��t�}(ד���q�*�A�+�%�խ:Sm͙a�n�S�Y�_�������Xi6u0-� �'�"�LC�����O�L�&�Q�����T��&���/�(�|17l��J����)�0���;)�w��xj��<� J�':��¡\m�8)'�n��|��䦈=_�f�J��R�e���� �c	���ـAkP�$'��[%\�t�I�S���8�	(�?ɮ���&�
�ة�pbe[?oE���@ )P�*��GzM��k��4hX�B����'�#�#�}т��_ h�PF�n)
��\��&
��"�T-*�4G�O�nY���K{�	�JԄ�G�� ���z�}�zvλ5�C��@�p��P�4��ԧ�2a�=��́�&J���D�k�����"c�t<�c�fG1OӺ܆W�za/Ra_�X�p`���o��V�RR�PT�n;f��?����Coۇ>�E�vT�n]1�h��H����[� �_���t0c��_k,l�@�.�<`�����(nF��D�L�g��9�)�7{F��']G�;Z�LD�~�)����jq- #Q��M�!>��U�p�oo_�.E�5d<W��8�-����!P�v��g�m�!��	^�
�p"�;��C ����`��� q�W?�	�=e��*�����Z�R��m3 �v(D��8����RF�U��U���A6"$	�C�[���6}X8��;���prj/ڗ����K�YM�U�3���R���19���}��������$��������Es�x�e-������.2:�~�w0��\Dfג�,Xom�J�E��qϩ��[���z�q��:��,t��E��8c���!�`�
`5:�L�QT�HJ�P�b�V��7�A�fG����2�J|������Å��m?�H׏3k{�M]��J��\�܎�zD��Z,��1Q��2e�r9���X�ce��Y��X(�zI^]O�S�u	_.���ެ���"���B�#���_���Џ�s���޽�$���-?&l"��PD�9P�����
:�����y�9��;�w �4�R1�؝��
	F��Ƞ������f����O[ѥfSwFz�_9�aҿ؂�>����a���*JaaPq�z~�-�:�0����躧W�B��V���a�Q��W|R�������=�����O��}uo W]ӀF��6��X~?��(��$xÏ��a�"�����3��&���؛���fH�xJ6��D�C6�}׏����t���	�ab y(�_�p�x"�j�o@��?���&�P�r���${i5<��ߑ�=�Vݳy��xps��uysS���<�
1Cp�s}�S���y�!X�5m��}��Գ���6���j7ԗ����8��N��@���nn��y�@/ŋ=��"�aGx�.rq��h�y��Ϸl��fP�����V�tr�����β�h�����^\Լ"@���(�9*g&�8%�T�,�M;����SȌ�ԟ���&d��NE�ZLz��K��q*1��,��>F�:=s�m���d9m��vM��'�҃5�f`8"g��s*������aO��Vo�� x��,F�w�W�f��gT�
����ͬ����}���ׂ�5��\�:><��)�r�RѷC-DT�6�~��˃��ƸG�.k/]�'
S�����}bxF��Ս����ISF.1�O�K��f��c'�x&�_�%��NJ�COf��SC:���؆X�~q�AK�)����1�^b�p����h�15��CV����<�_�U�����F�ׂw�����G��|>4�+1��=�D=p��-Z��"��a��gB"������39Q�%
��n7tW�C��d��a�xl�4]p*��G=��q� �6�^�F��Y@�8z/ۼ�O�{�rT�����rl3�W�va�v����5! Y9*zN��2�rܴ#�G���/���т��y�#%l��
/H�?Q�?�9�{R� 8�,�e+ށ<����O�0�~b�a<���O�%I ��UH8=�9G�[ē8������\¾d��ێk[���=�%!���B0?����g��Ӓ ��� ��I��O9�oTe�$^���,�CD$�=r��n@���P� n%Pw>���S�*"~���Lh�xO�D�Ag���2��F��9�υv��|�~���ɗ/�漭2Z�)���Rb?��m�[��:���0���"��o)�*���$M �p ��N�C�_Y�V�6\�$OHCδ��;��4�k9�轕b_����˩��5TJ��szR�պ������x�m�M�6h%�&�O�?tO(J��Z�}΀b�N�T�Eq�-7��{a��A�{��%H~���5��_�������D��><y�tNǺ���`Zw��GS�n�����A���r���r�a�a,ZH���r9�D���Ff����h%11�PhÏlR�
'&����t��������c��U�cF�W����ٍ�VQh�������!�
Pl��?Ν۵ֺx�����,�Y�xF�-�z��^�4z��\�6�hA���k�ۻcW1����0�,�Q���>��V�`h��� SR��t�
���Ǧe���������DP��0ڴ�}@ ��C�j��u�PY;^���E��f4���M��I樹`B9{f=,��>&`��8"��C^-��'c�! ����*��M)���@����U�X��@�A������,�U�T�<� �x�Å(w����`�\���#J.���^��5����j
/��2��g�Y����� FZn�g,j�v�.�`,�]A�߂���찅���[��|�8���]^r��٘�{�ܞ��!'�ǈ�
���=�4�{a�hmG"^��L��]w:2��)�����s�MR@I�H���c��3��0|�x�/)�S�SbQ�8ʩ���'v�$�Fn;�j��$/��&=��a�Z��J��-����$�Ț3�X��;iyה�T覌PD�2����m����%@:�f[��-�A��%��u�S�d�.`k�U��:u�_��d��^����	a�i��W��<dp�w����D���ԢQn��g��������B�f�����p����:R�5?��1#�ʳ�r %��S�����+�o��B�@q�q�s�a�%ii�l�|T,L.�+�KFg���7p��z@o�L%,h@tI7q��}Ξ-�5>�,��z�d�����j0��U�u�'�ZOJ��VS������~���膄,E��i��+�,3)D�$Qn��J�$[��ju<!=|$�n���	� �)fΈ`c�D<xw��1L�[,�Qy���� ݐ�
�ya>�=�PE�%MB禒�;
�)E�b����[�b�Z�Z�Wq>l�gϢ�mV���� �7��I	$X0�� F��!��#A�[v����.�g�!+*qL�_�t'�K��vT��7 ��M���͟[i���[���*xT��s6�*6�z�k��V�y��
�=3�1 ���~{@&�B�e�j8�Zlf���ɥ�� bE������XA�r��a~��~wT��[��'>CSH�v��?�zY\WW�_�,�D���s�1r�6�>b)���F��3;2d���9��!�N��c4b��U�fr�d�m���C$Uv��:�]GW������Շ�N4U�r^C.چ�wAm�?o�,16�P`G����2���N���䀹�Ίr*�c���M�@�#�U�B��p�^�X�1�>���^i���VӶj� �t/'�(_�?�&�� �H�Qa��'é����w\�	 ��Y�����~#�`'�wx�M�~A�y��"`�]ԟ�7jLG���1�CŃ��y��zy�O����G�u)"n��"ݒ{!��Ak��������l�m<�Ҫ�ڹ��?C7?����\���E��zB�)-�J/�F3Θ�'�G ��pCy�wacQF�0��>r��Z᩺-��Е��Zq��T��m�n�ai�5?��i���5��h���[�x7	��,���r4��y���9<%/�d$��7��*�f�f�#�^]�u����':U�?r�?<zZ�~��>i��#�d��W�oz@u9Z�{�|���`P�[�R��d�[ZӺY?q~�r�W:>�צ��2�8����� ����"�N�f����T����l��g�Bv��)��O���}P�t$�4�� fe�{��(F��_0{�B�D��{�spJ�G��H;į��xSP�\�9.�:ޜj��(���c]��2�N
��dQZ3E��vR�F���lOs�Z�F��uX���x�0C�
�")jd�A,����P�������:�n�YoOC]��G�䐞�2���30/������z�:�����茄���3���%<�ٞ�`���ۍV���k}�xǥ�� !w�;^�s�����j��r�{�|��5A���9�6*�3�9�`Nm���F���4�`O��jW}#��ĠlgY��},2�u�􊨫�ӧ��))�>w��v?G���,vg !=\)����Rǡ3v����&�%缎��5�+��ɳ��m:�,�����\ ��ic�[6����������$�n{��U��eX�z�+۞��t���?`T#Ψ�(��!��n1'�6u�g�-[����!���_T���w��xm�E�P�H��:�w����H-N�d��������������1���y��b:MTH���w��<�º�!:�ZZ9�qn�;�gOi����}�^�TX�H���n�6�јTS\J�⃹9?=�!��G�8SRZ�~�3'��8��]o{�����?q���F~�6qE�Ҩ>V�3W|�(�1�6�e8L�y7ů1��W��;`��31X�ӵ)��ָ����x�c_)���,� Xqx:n���>:xs6)���;����d�n~�l	����;f��.����V~��^�p(q�������e{�Xq������Q1Bü?%�)t&��H�liN�,	�?�/d�#��\ 
�F��,���$�|�OH��l�+z�. �H�0K�ZF�o������Ő��,�b��d��qL�_4Ž�lo]#
h��5f���钭P.Ɇ�X���P�ᕘ�H-��oi��r�����qׇ>��XjZ �E�� �M�+��⥾��J���dZE⴮�<���C��,��\ț?�;n��!�*�RS�/w^���u������\�0��G/��߿X�wzE�Ӛ�3�VҜ��g2���(���ϗ��y( �Ӈg��1E��=RM��҂�`�q�� ���ݫ�u�n	i�fRdM��+R(�̻|��D0e�vf�KT5����[�=\�X46��s�ż:�gsTP �{]%��Ů���x����2�J�76&�-ԙw������C� Y���/@8gJ��w{��Y,)k9d�Y��ݮ���&�\� p�9�56��&�O��_��_+�k�����<ܛd$�^��m��g`d������[�J�$?�$Hf��[���-��I���!s��]S��3o"M�ɨ�ӂ4�M��y��l�����2wv���r�`\.)HP���!�Ѧj|���Z�)x^�W�}��#��sk���H��{ո:��6��s�@��H�9$��^�+_�`cK��j�E��g���:ߣ�ټ�#�:�֘?S�\��f�?S]��!�`SH�|���-Fy�OmX��7qJ�a����˴�x4�ޯ+#J�0�k��s�3�I�f��A-�|�	0����m��xO"ϴ;��˃)o�*{O�����fυ�L�Y��m:A<��J�3iS��W ʘ���ۙLD��1��K��ӳiO�?�PM:Y�JJ��$�Oٿs�KxHl�F�xD���uK��o��~�'�y�q����Kv�;S�/?�Rq��L���f<���-��STN��>d�½�	���m�v��r�2���'�cQ����5����{ȶ�Sy@���Yy�&��#[u��]�!>��gp���NV�t��as�Y֭�Xoβ��d�.�"%WW��t4F\K��Oh9�z1|��`���]��f��^����Z���g?_.�l�5�w_���z`3��i�G��&�X��������Dh̍ttăO���F���F�7=�F�2r����o	z��~I�@�H�u}KJ����*a�����]���g�q��T���UQ�D�4id�i��jN�S��c�D�w�w��_�,�qK��y��Hs�����z(�P5Jl�"Gj :��K�~�v�d��R�νZM��UW�X�����ZTa5�������C�o�Aԫ�^M*�C�ϵ�Eˣ�5����ь�"8�S�͟�A$~@r�]��
>*w�u�ok'�Z�γ�_0T�͓[h�����0n��ƶ�	[!R�	2��7�diB��K���ωC��z�!��'�V��R���v�ôU�v��L/=�q�s��ؒ�yʒ�^r��!��fS�K{
���xA�s�%8��"����ط�D������D�I�-�h_hMr3X�xy�晕���뚥c��v����vISb@xt�F~������qWN���=��͢���K� ��'o#XgT��j,:\S�BB1�Ff��ؘ��"�$MY	������R�K�;x|q��!�~���AO*i��\g������=n��6���s�R�/5�qE]@F��6#��6VކL�e���=6�pg�?����D���h���<�4V�L|���R���$?��x���&�\��~���q2%���+�[}]ݜL�ډ<��P�$t�l,e'��ƹ?��s�t��*k��!���hj jeԊC�L��tXKu�aUDz�0�ѿ�����l�-.{����i�E�+��L�,��u
��%k��3dߕ����I�_5��;1"rja���D[�j�zit�5�.�ʏ5�딢�bw��h%]��kE�0���x)^���(�
> fl{���EU���rP���v> .�3]`�'{j��=��A��2�}���AN��9r �e��$yE��#�?UrȘy��Rvg����@ޛ�{4'�$Ї=�����]�M'k������Y4��N�	#H!]L�8~��'>��	���p�7����w�W����p4O� 5���#�i$:3~>��~�:������� �W��fK{%���'�_�$F�M�W7f��
S���8����ZG�#���ĊR}x�<�K���z)���.���Cs��"5s~��x��� D�q�?1�U}2�@�y�h��/Ϟ��w
�ɿ�����#�\�3f���W�@I��B�׍?)&f7r$c;�}\p����j�H:��a2KՊ�b����y����rD���{I�F\Y��i��|�zƠ \�����<s�z��t$��)�$
��/-�����H���g��}��V�-��ԭ'�<�(�GQc'��3���c�aB�nۉY����~�X_
c���M���l�1���K��vFp����d;Q��%a�u�B݅�Q�cSx5Q5����q�<�?�z�v:�Ӫ�b<n9�"�U���Hj^�Ѵ�P9W�v�s*�F���z�`0�C�Z�zK����#_B�����S�R����<���`�,���[*ʦV�$6���?�����x�ӨTH�ٱݖ��)���Q1�*DX����Ѷ ��S{���&�&oAa+L͹��e7������kڵ�Dk�+�8�}��I���#��*f�h�'�˾bwEU�E9[���[�&'�*���m���Wv�l�/�m�+�����A�@-����^M\r	&l�P�'؄�VT��&��.3�-y��~J��iV��X�W]f�4i")࿞o�*K��=�sr�$Dg��xl�d������UfX�e�a`X�)���y���P4'@e�M�,X!�4�j�e�|��Xh����(�e��hF���h�y�U:�'h��#��Y+�N�i[���p�l��*2A�p���l��ɿ�ߒ�%���{�h�����T�%��\��2+p��W��m��Ke>�x0�.i�s21�8���U���b�8$���h@<X�%D�x.���5��"d�ص]��*�_&���= �7S��[`Xs[YÑzi>�&�X�i��rs������~���2��uO/TK�p��(Pk�t���7"�7]"�T�l�&kw�[�&7�B_�E�|~0���.W�HL',���|���55Iנ]e���AhY]0ꈊ���n�W�����MZ�1b~j뢆6��bmdS۰d3����X�_� Q��˽�0�[�X�{i-<�כ�&�0S ��;�ųK����c������	X-� %�����@3I�/�4Ar�`x�=�p$�^ӽN${׬O���Б7��
i)�s3�Q]ZZ��]}��ppZ�&�U�����.9�n~y"���KQsbʩ�ppQ�9w>����N�#DFml�'vl�٭���D��e1��S���@�⣎r"6�>#,x�,�j���BÓ��,`��ȵ�Ujs2M�h�=��K;��=5��5�r�5omȺDog���c�\"m@�bۏc�<�ޔ~hڌ;���R�;)�����c��"3(��}�9�=�S�[^�8�+���lKl��D��i�k_�D�0�;��K6�阎a<��Wg5�k�1i9o�a��M���3`�+�m`��iה���2>??F%��9��l+2�/���s�4dM����z-OW�Q>�N��R�1S�!3ȶ6��tj>�0�\hT�����Z���O�D38G��xz�Y��#�/6�������Mw=-�ܲ#�k�3Q��x��Q��p?.�?����@�0=K��>G{y<$�N�"Ű��PD�vBx�M��O�w>F����T� �����_����&���ϣՍ�'� (>��Y�WP,oYY�2^�m릒�Z�X=6��f5K~�*B7Uu�l�ͪ����O���#���@A��5����1�֪W8��í+�m��DR��278e���Y�H���>�p��ą_����_=�j�x��F��n%"rh��G�A(<c���8�C�	0��Z��
L6��j(�)}T.%�� {C�s��4FL6�0z2L��� °����}������@Cd�;�*�lb)��t	[��&.�U��JH��p<�DS��@���J`2�S����W<8�aEߍr�ŵ##ZikUX�e21Ċ`�zr�l���R��E�m%O�O���X�Aqj?��@ �n�?��|�{f_���ԓ�1�T@ZCyQ�b��!�/�K��Ѳ�m)�<;s�ʹ@$;կ%f�� @mKgu}>�d&��L����ɣx�&T�a�^�pCͷ��J��u���I[��l�E�H���nｃ�ˑ�T����"�rgV8��۳1H�82��bT��@��|��}�R�����|';*f�cd���b�:����$������w�"��e�Ph>�G�2��ɒ?"���R@��#��W8���h�hq=�ª��l����\��U��q�ag�ހ���nu*�L��g���_A���a�,�3Q�+Q7��n�eD�K����R��*���6K���C���̱~~�Т��&j>׋!4奤l���]i�Qq�^�6����n?\���	����W��:D�:w<��1��ʢ�r��
��i�L}EI�>{6hbV>�]c7LVBb�������-W̓�0}Ǳ'ۊ�~>*��Q7��?�2!��\�?����oa0nŸ��ZyO����d1{;�S����3,\�RBz�l���92�V/1+x�c7�t�>���@ ��d%w��쓡�+�G�/��Ě��LY��uB�8r������[g��f��3XŌ`�Y(��/�{S�*'|w�n'���(C���vd�&�2�Ѫ�^�!�[R�;oJ9\͈����3X&c��T��^�m=2�����Ζ��k�h��b��*���83ZL� ��ˁ��SǄ+0�����u�cߑ���Zf$�݂��O���c2<b{�a���H@<n���\.��r�~�|d8\ؠY �/.w��� U���J�|��j�C�W���d
~�8�
yt��L�Rr���R��]�46GZ(�8a8MC����Z(m)Y����]~!E#]V,�#��3݈�ĬNq�A�߮^�K0����u~� �n�x�dەj�Q3N�p7���$���NJq��6
��y�v��w3�����^CeYe�'!�9.Z����TF|;ror4[��z��N�wQ�ǀA��"�u.�E�7׿qTW2
=�%O�/o���ܻ|�*]��bI��,����};���`W|k)�]��0h��,�=3�h�����Y���-��n��h�:Y�{�-�L1��O�xp(�y�Q�Ǯ�������yS�V����N�A��?�e�d�_D�3i��T��T�=@�NF#��S�\�O�y`d	��gE�*T��)�.Y!���Y|�Rg{�u1�q���-|Y��^*�)t��ޅn�Fx��o3&�s��A� ce�1����`�K�]P���v�Y����v�jˑ�؋�o#���Y+���{����iU=Sb�L]Q���Ú��DP[��Y�i���Vڸ�o'Q����F�0h��V�VZ.��'��#5g4�V�|�oa�,�	n@�Y+��5w�,e��'1_]:��J��bF����AW
��ٷ�Ƴ=(5��)#� ��y%�}��'��$Q��@K�O4ʕu�5�[��eq:��߸FR�-��^�I�JH��X�z`��F@~^IGE?�=�hw�� ��!��Z�������@�C�x�������9�Ay���_8Ĳ^Je�8P]�Y�c�.��h�{n7ǂU⍰|n�_3���}�E�z�S�O2׺[8�|�y�p��c�O�h���}D>�0�GxF��.�z��l7i��&��]3���w�^��u�{���r�Tʩ:���;X��Z϶�;����9�{�]h����xLZ��=��'ku�1*��]*��YUZ߲zɏ�
��p�s�@�La? ;�b��������g8�Ub�0E-�R�����_�zk���{�$��`���~�oh!�WL��-s߷��k���~L�³�@��d�lW�Q�Э�+aKqT��4V
�����9�J�ޅ>48t��@�+_��غ�M�u����3�-����e#��qǑr���("�����yH�G�@����GY���Pg:�{����~#�y�5�443���1}}U@�c�n��[��WMO('/��+�T��M��C�d�q���:c�ׄP01�~Q��%M�zK7�BOEJ��qu	�����qT�\�tc2}q0!�[�n��k��i�ۊv���JJ��V�/��?3��ر�wd̓e�_u���^qB�o� �$jV����7�x�xs�ҋG���w�D�t���ҟ�Q����|��1~w�S�)��а;����l!�Ь�]��i{��[&},KGY?R�2���3����k$P��4��)䥓pjp�v���v]��F���y)��5B��E˿Quo�S�`c�!-��B��ѯ����ms�>�S�\�L�$A~|g6�jMH'v_l��'�T�^����/Q_q�w�f{a&�6��I��ld�Mԗ�J,Y�>Q�d��ni�"��L�6����	]�o&fT=�Ep"����{?|/!$M͚��/5�����)�4 ()��I^���b!�K�>6��B
�0tE� ?�Y�y�D���Ԛ#x�����ݏ��b��^���x�������l��U"�~����m8��mË�l�\�3,�*/J�b��xDpR�b-+]����l� "F=���*ѓ��h��؍i]�Ǔ��MB�'Tz��=3�����ls��PpڵS���#[���8��X��K�ѯ{�b���ʰ���s���I��)��,�6�������A4�+�m$ፊJ����������r���4�)LcuCҚ5l3Y����|`�;wJ'&�L�uk9Zjٗ�g���EҞW䯐��_����tmB�J��;��zf�b-�R�um���i��f�) 64�[�8��W��K�nu^�$J����;�S<F�/�S���������D��d�L�/3�d���n����&��v��Ȗ˂"�ËsH]���rb��8��~Y`ϔ����Md����^��8���ԭ_��Rp�Dj�ͱ�>�e	Z]{���K���H�U���Э�O�j���~��5W�T���EqG��f���葽pP�$��i��O?�f#�}|�[�����6e� �x�����ۧ,,��KέQL��%8��Ʌ��fAR@
գv�8J1Ntk#��(��s�蚊wV ���]��]`�Z���։�� �Q�̀��9�\L��S���Iu��rx\Z�'ΡT E_���枙qh�[r{��cXa�ż?t����3����$����Q� ��R�	�ۯ��$�>蝱�DQf}�j�M�X/�-S��wW�_M��ۤ7�A��46OH����,�� *��(v��x�8�X������E\��{<�����.+�ۦ�P�8�u��G0�|��;��@Ђ쮉���>�/1����J�!-5dy�8�\�5�
o���T�=�c��R%o?Is�>@8�z��>F眲b��b�X'|_	}�l���RR~^d�Z���}v� #1���}���j#��T�	+č�`�^ؑ���-��A�\qS��_��IH�����u/v����O�Q� 8E��gw¤�O�-��~F��������c�H|qds�]8�����J�K�6?�š?���E ������W��dzOo��m��e�D�;���2.���,D��t��1���~�}�il�L<>�^��kȑp�=p��u��/���~n���:&/��{�>�Z�p�3-���?�ú@���f�A��8y�q�@����H'��@��a%)͝��/2�ܪ�3��ؓ�P�[���N�P���Yi�c3!��Wn�7����2�B3U��>�<��*���9��kq��Gi%xBԟ8�� ���χR����*�nv���	�c_#�$(�-����+�5��8�BPǡ�H6�O�I��F���6�͝���Pa�9�����_xbYY��2��j���F*�>ի2*T���_4����v�:T�'$D�u�����74pӌ��@�*j����B���H�d�T�%��\ϐ��8���h��.�v�p+�Cp8�L�FˬXz�c���`��_� f��h�gܐM�Nn���;�"x@���~���\�~E�t�m�����d<ad���u�'bj���(��BH�A��?#�N�z�Ɍ�ݖ�d�g�`��,_%�:��t�ҷ[�cJ
��� Cy^�KZ^o!ĺ�q��36���;7Y/�-�Ni�*�fE��A&��Rb�e���1=}��|�Q����U�.�<�Á���(M��V��N-�`S¶��aU<Ҧ��/�O̲	�Ye+�r�[:4.a�=�AU��2ū��z�<� �D7��*ކ�j�&�0#��߿��t��Ts���<ހ�H=B|�a~R+1� �f��%��G���.�@a�D>n�w��gi�� !�h<��w�ǘh��A|��aI�G��p�v���4�1�A*���\�UJS���t{C�jY�ҁ�aǒ( -���rSbmҀY�gAWJb���b�����p���S���Iߤ܅6l�|s���	]CV���-�#^l]T�N���N15�	mםb��hY�F�2�Àձ�
�<�k8��*{���������G����n\�a����a�pp���:���h��L���D�����G�y�"u8)�*��u�N��t��FK�����l��T��]��W�
�F�_��q�_�߶.��l��	�e���y�ȂG�w�/u:��Q��1�yɰ�Q�!���a���V��mK@R�0�7/KA� �ay?5%<�Zd���ف
�U���r뷷��%A�w@����ۑ��]Kވ�M<��"L���*jxN����vk����ل�e$-7�	��]��9ۗ�� ��q�y��T�ry]K����E�@��KT�.�||R��Ҏ r�J,��"�6�ߩ��� Bx���B����>���C�5��Kc��k��o��U*ݽĻ�Z9$Ǒ�}Mh����d��B��;�~MpBZ��my��9;H*6�ƃǠ���� �K���N�ӄ.�����/�c^����a��PL�u���b|j�d��+J,�"�.*5|}��Q��{�n�l$�`���M�V�I ��GH�}dߐ���+?����p��"_pޙ����:��hI��C���d�f�t�9*u�Cu���Ul����+�S�)��ilV�:��pD[e�b��<�T�1���ĺ�q$�-���3=�FFg�j�B�H��mɡ���.~��4ߴ�X #W%\�o�����?B�~	N�������Ok,�2v�KVƭ����%���G%")�k�1M��0�Je�G�u���B'df`������0^}�����fI��Q�qS���`�K�}h��⧗T���
l�ý�? �����
��=�=���ch\��ۃ켞��c�9�D�D��H���C�R�/�:� Fy���<��	���鬝=�ى|�{���{P���
�M��'��.ḕ$		8>�p��'�d�f��C��]ѳ�X�S@f��4�㪷J��A�<*8Bxe�� 	�6�V@/eI�?g��FaZG�:�_lg�LV�"���S�n`��e/ʌb�[�����Ͻ#�P�OS320*Dy�:�#7/��{f�����b�U��j"�~��|bN�\l"�@��A�✊�l��y�C�Gv�M[��p�96;��,�8߲ƾn�7m�˖��!kl_V�-Z��Eg�m�Aő�:ocl����u�����o�����1����NJ�t^i�!#2nǀU��J�o���0�[�e��
�	�����ݤ�$ILV��A�w<u�?�`��(���Q�\A8У���c��l��C�Rr��n7�Ģ���ef�� �F�{�� ���|�n���M��:��2�"i�w��+vgJ�b ?��d18��<��z�b"��_��-�6G�ٰ��Uj�k���w��#-����ė�E/���hj������������{xb��݋\X�k5 �Za��!���Q�uTI۲��h��(��
��O�j�z�G"z:7��͜��, ��1�1@]ۨ�,���露�l؇�B��˜D���+rxmc���p���*�A��UnÅ��9����m�=�Zdn3�󲈎��c��N�[��C����s! N5���NطO.k���]��Lu=ּ���]I�Z&}O�~zqS�r
��}���a^�Ҿ)[�C�.c���WjJ��bf��]�4��B��Ե7I��n���9��j��<N! �-�a��1 ��F�0���>,}����H�K��[� ��8�<v��j\ZK8�I�w..�U3��l��p5X����Z��)tE�����W@�]s$z�������kR|����2�{͝Wʒ�Z��Ɩ�L}�n(��)��'*�E㪶F�(ؠ/.�j��C��a]�����[x����/���Nԑƚ[�s��,;	L��績д��zތƁ�������B�#s�y�1M�@?�_���%�茎XW�C:F�X?!�	:��K4�X> 5�B|Uw  �S��kU��G���HX*|�@p�[�Qq�>u�]%��BV���z'��}��ɤ��\&��U\\`�V
9�E5� C�[�(���b?�ƋQ��:U�l$�y�򳥗�\A��ȤBs������g@#G�8�N�u��%W0�?VL86[ɱcɱS ~�������O���68�ï�X�0CW3S'�*�C"*��~bB	��u6����V3���~��婬�T�d���`Ir��s!6���l����ڄ�P���ٞ�8ıZ0�c��GҎ���n=�Kx� �����zZ�;=�{J����3'���ob�1����TeIs�!LE�[�X��q^������q���Q��l�m��ٸ����Y����/\)�x�T���8(�~/6�-g!,���ٌ��"F��r0>��|��a�#l�p�B�/!�R��]u^���F�q���Y=��J^�A�;���ޏ<�ы杘��� Wn	��K�y��i�'���=�~K�ӽ�۲��e9�.�!"RC�L$;[ّ�ײ/O�G����!I�튔���NǛ�ҽr1Bg����:T(*;��|;n �  n
�7��{�f���>�d�p���G������߭7�#�z�����:|о(���c�K"#V$Ka�����h���wM��t�
n����qTp��ɥi�_���+�Q0:7��#�+8ArVq9縈J���h����CKf�� ��"R���/�C.�l���N�FW/8 S����D+�Ɛ���Fȩ#�p���Q,���ni�!܉�@2g���������>�lLzH*_A����T>����m^�֋�ċ��K ����
ջ��d{_�_�8��:���N S���JѶ��d���>Qr�����0�?t������U=Z�B%�1<Pri;.�yG^����iW �?�-lJ��Ct�9��������'��p��{"����_�h	:�$�.ud	R�_4���۞��+��JA��T�ž�j��d���_�!�D��5��jE�G�¶�T۽�k�xi��v&�b�g���T���=���	���d�0ƌle��Τ��z$�5�g��n覻�e�=,�]\)޹^98ɻ�50�]�8���&�����Ş��׼�5��b�%�Ԗi�5�fB��.V�/��`l��e,����xh<�K�T�c��{�wg��h��'$E�:6�$���5�2dIc�{��|hoom˝� �A��V��@��P/���O�����^\�C:���j�!fY'��"�=x���LGn&�G ��:ɗ�?�����NS�[ P|t�ɔ���ծ	NV�u�ȹtP�@��ʟ�b��n�MY �T8�)%/�q��� ĚB�������	�N�_����cP�`��cM�s>�.��������O-_;�����9�y���e�هӉ�C7ʸ>8Xj{��(?����t���|u�Z�"��:1��_$�`
���<�z\�A /�)Pn�73#�T<�x��tw��6��F�n�LL_Z�¨��m��щ�݈����b�4��  �	;�Xؖw�LԵ�N!�9}�� /�-|��N�t<?���xE_��Z�Թ-Rg���hF�l$�Yzҟ������l�?��[�$�Y�3N��,�M���8Ztꁰ�3���;�r��"t)�q�
9P���9g���aٽG�2JB���a�ڛU�B̫��FXݍђ�X���h3h;�w�n$��BA�@���s^ RK�; z��8q�"�����q�V/sێ���(��,���<�F��ub��xQU+d@��Y0�ë="�k������a���κD�l���xe�y^�1+�2M`�v��z殅FJiO��6��]�p釃us�0���u�E�`���S2*J)���
���V3_=�Mq^8*R_�*җG�RH7�/�h�c�)���{5�2��!{����F�z�������������>���̫�{q(SŜ�0��0)����"P,���7����Ν��_r錼=j�#-��B�r��|1c[�꾳nɫ�R#פ���?K�8.�=M��*|մ�|'�����/4�'�O4FT��
�u�X��݆�b*��0
�A�9�q�QX�����J����v��0��ޚ��bf]����VǤ�q1��
��v�&�gJ�sI�$�e��Z\�0cy�̑2sQ|�jݖ�Q^$�1��-�O�A��Aq>
�G��03��V���k]Mz�e��Nj�����������r(B_��0n�b� %�ʵ_�5�����=	ǔ�<���ŭ�e��7�ת�x2�  xUj(�rU�F���n����U�o����U�Ť��@$��ys�JQ���T���2�)e�ԶG#�%]Oɾ��l^�BTZ�ko*�|sd����c�ƌ������^�k�V�����*2��V��.4I�('D��&և|+�'�Tv�Mh)�;%;?���0D�+8.*�} ��҉GG��1f�rSe��.W1<�~)�	�������L�|&��;z�1�.������1p�ɐ�������4qbH��q�r�x�}C�r��D�N�	ql�~��h�������Μ�
��a��m�z�!:��	02P;/�}��5�Qp�*ڻ��[%�[�K���9��kZrk֨��P��F���0$3�JV�S�Z��g������KǖkD[�<��Q%�5"�$p��j�{[�������I�m-~��\I*�LG�ۙG��Aw�Ϭ� b�8��[��|�A{�M8*Պ7��i�
��������)�k�?�Ґ{9K�׷5��%�`��$��1�8�aE���q�&7)�.`�"?��`&����	Gs�κ-bV�	p���p��Pz3����A�q�N|<ҍr�R���\Aݙ����b̡��C��sxG���EeE�z^��*�����u���sj���V�MP~�#^�l�� os��1�s��R�D���V�,�,8�'YK�'�owڼ��%��L��k^�W�З��uS4�y�t�U�[@Ϣ����S	�M�{Rú;���Q�w�v+ʯaV�Y~/?f�i��u�C8�x�F���=>Xm�q�Y�t����B"�͚����(k5����:|j9��; ��O�)�-6y�R�����ԙ��s�L{+/&ߚ��m�q45#�J���i1�v4���I��I���s�CKWi�J������%-��&r����`2%��� N�n�7Y�{�r���zmե6?~_�4�����j���/Z�^k�hD"�au���6���8 ]���h�2^[�!p���.��f�	�����S����8�ӵT���aAK����n`���	���'��Q���՟r�C�";��Fh%z�����#)���k���s���w�e�9XB����M�S�ޫ�ȧ:�b���:s�]�:wLEX�ځ�\{(4o����8O������׊�M��u]�q4��p���')�	'*o�8,��8���@n��?���#�5����Z-h�i� �y;[$p�נ�F��T��`�7������Jm�������E���1m��A��-�O�L��K����u����iNռ!�z��s��(\���L�d����`�yxpz��r���0?<��U)"���:�_�bow�h�ĕyخ}Lк����M���:��uh��ό|�e1Jb
���Y.�7/\�m���q�x;�?��`n?� v�;3t:���r�P���u\ēb�V�������ex��2:'�����-sg��8f{T,���_���E1*8�y�:s�Iή��+�#�����uS�'����L~��YQ� Ʊ�7͎Ƌ��3��c��j�|�~dQ�@:�,�|�����Q��b1�¤8�������?�����Nj$���@��u�wt��!x�%<��9/��W�Hbk�V�EG8���%����g*U�h�q^�7\w��9��U{BS���4�K+�Z���Ӓ����j�c}Hj~n������0K�o�~�S�^�~���إ�*�X�����tX%�w�,�����';U;�m�*���]׈ �3��G�׌Z��rp�������Z5�6yu$�������-ҁ*w,6��=
~�#��9'���B�����hƢ���H.���I��6��7�SV;�oQ]����$zYx�s$.+dA3h#����ڐ|�~'�TI]zZlS�Z^1� 7�2�Ͼ�E�ŋ��9Lz!ߖ&��^�L�JϾvj�i#��|���8�|�ل0�k�c��7���cN��'i��uy� q�XjIP.�-�Wx�ןb�@�m�S0��Y��423W��m�!W�n(\R�{�פs�����U����!�e}L�B���E_i�_�h�o�����XS���z{0鈙HU�y����@��ks������:�04��W��m��F����P[0z���B�5� GҮm5�w�څ����'�?�ߌ���7�*���C��}i�i����x6Ⱒ�
x�-�����nr�|��81���6ν�WÅ5�ҷS��F�
�ǭ�{�wP�윪f���T���=Y��ę��L7��+�����3!����R�$V����a<<�:n�:�eU��i��r��~4� �ԑF�XG|u���������ӏ;��2�H��"IF���ے��?�uw�K ���]�DY�?�Bb�̉j�;㘃r���v}�h@�s�ۘ�������Y/c	馝���}p��єC��!���Ʌ᭬g��ŏMQ�ԩ����hU�.(����m`d㒩gG�k�B�B�A?��A�po-9Ks��# �z���=#���x�L�����D�G�m������4+8�o[_Ѽd%YL�	������r�P���/󖚜�|�
�f�:��w�֡��4����aX�Q.�a��w\�zCzy����ԁS�B.����V�%��������x��%�W���>�Eb�T4���=;�O�f�wQ��[^�̈"�
��lqhJ%`Y�y�ĠQ�%��/{�A-	dn� �+��(��<D螪TV�.]�.��r(Z7;
ՠ[��J��4N���(i⥰�� ���[[N�<�5"-o)8PhU=����E�R�V�Q3cx0����W���֠���b�¾�xw;����R���� ^^�u6X)�5瘄�V��l�������L<Q%<��\cL�U(P[�g��ER�3�����-�7�#�S	W86i����V��61�_�y���"R��Հ�x$�36|��ɣi���FސG6�e}���ɇ�m���t��Z�DCn����	���!UB�A#���s��l��^,)�y��?L�1�~���j4��D�l�X6˛�Ď��2�с���ꤜ������{)��%�Ú�/X{[�>ưya#��5VzD�P1g_��T�CiP��Ԣ�����E�z@�@�d;?��)U�0��Y�J�X bK]]��툁���t���f��2�@��I���g��t��p�D�
�QA4n��L�]q��F���K���Ӛ{��}O���^��SU{A�W�ܸP�l�8y���G\��;aquo��Q��%P���nU��)?�ӥ��H_�S�Щ�Z�BH���
'�i�3����1s�;b>�P����١�xnbO8f�!��}d��&��n�:���b;1S������	+�/��cJ׼��>iE��=r�f��(��;CgH���K�c� |�����"�%h�4�t_'����q�!Շ�����(c�N���󆅠A#Ń姢��bW�B��N*�8\)E$D¼[O���bޮ�	N>��je�@y�5!��r��f4�. [��p|��Z�������*��w���|z?���!���<1��uDG'�y�`W�|	�횶������t�ԗ@�Eͥ-��=��M�~b6|�X2�4?ےw"��}�g?�@�*_V��˒��C>��9 	����T�<���������<J�:��`I`�C�Zx^$�E��L��Q�]v\�(^3��>��R��v��(�yE�Z�ZQ�V�h!�|�\x�G<�?D6K�wE9�]�A�]Y������J�;�ȠH���v����E͛��:�MC�V�m�9Ip��)���GX��HMXY����s�Ѓ���������V�Ͳ��E�g�!�kߝ��P~j�fI�a���%�Q���7�a�7:4p����/'�١���D9q�B��� 9�,k��9qr�f�e E�1����#r�LI)������&�mȸl[T+�G:��Ƹ"!�n�/��Ф����קG�w�?�*���<��F��!b��T�����A�1�=��_��0j!k��Y�<m�WݩN�Z-�Qe#���U*�(�~gA����#�q琻�J`a�z��VA��<f��%�,��I�d����j�v�f3��Ė�1NnӍ��jsR��B��O��r:FB��l>u��������x���"O!4�ǚ!�;����[[6\d
���[{���,V$���³��f�|��6�2<��?�������~�6n�5�	{7I¯d�\�d�Dr4�,����(����вT~:�.�_��`���O�H)Ī��'�?��M��T��p��E�佂!<��8Rh�qK\���X�df�����P�y�c�F�� u��a��#G�b)� �8���ݙF�(��f�R8~AB���m�[wĪɗXtN+�^��y��C�>����A[�cW�r���}�K��5�ӹOĩY�| �]	�O�} #V��֊���ur|ӱ���͚&�c���4ʾPS���@�S@H��.<@�i��a�d�@%���O�m�g����Z�+�l�g�&����3GBt,���xB�EA��Ѳ�n6�hIɄh�	7����+�+5��3��)0k5�iCK&�<���#�,ɹ&1�iY^�#���y����o2���J̊	J�ph.��@���n�VI�p�6_��?Rħ���_��(.|9	�<�5	i���RVy=C�Sh�u���,ɐ)�_����V��|�*f0?�XQ#1�4r�e˘SA�e��Nb�^��U2q��l��?֟S�?#ET�����C����&	�9O��2��?�E1�Y���rC�;
72 J1C�~��W�a��Fy�|����������_��ut��H/M��'绺4Y��E�c��D�WaYN�l��-w6�r���ddzsY}z�?��D�1�+�L��
4��#D�o��J��d5�|m��Y�q�	�Q�*��w���[/��/��?,w� �Ĵ���AuC�s�Yd�h�$(�4�)_�̇��jn}�;^�����0;�5�(l��R֠��XV<�/������������������	i�L���&���}�+�ťǇD+؂(�K��6=�!��l[�2�1%�\1�!��(?�ʘ�#u�`�'�^w��_u�M�ac�O< *���Q���g����"���l˜P7�l���d��7$�S],O�SW��]�t��f�h�&�k�ɔ���F��a�v�����T�������8Gy�Z�M�䕻�h|�^� FA��=�R��v�5��6�(��3$b���-01�x`=�l
�Eh!b4꩘���J�քO %����(���z�Ca��G��&��>�#�Gd)'ϙِ�(����0Y�M7ܠ �&�EeP�i�wbX�]�{uq)NP���?� �>�KN�_��_r%����T�m��
��&1p�2���$A3���+#`�vWfIA�:iG�Q��u���v���z�1��+��K9GH�槕R�q\�!�Z�㭛Mٳ���a��ƕ>�>�%
"�[��;����a�IQD�w�ie��~�W��+o��lTܼٲ��je���X�v��P񧆑tI�����2D�R�L�]�F�3t=%6��������	޼M�^3��������0��[�d:��*�Wkj�8����+�Y�r��@>�=<��+� �_sёKCZ�~��K�hRy��/	�m.M7�'k�qQ�G�;*z�<]��YFSm����-�I)�����W�H��@�r���fOW��9e�fN�">�"Q\3�P >ںD���)�d�K� Oߌ(.'p/)�q�=+t!<���x`lor�z�f�T�"xUU]�|�"I�B�-(P^گ1�� B�����T�����w��A��	�)�Y`��q̲N�V R�uRڝk�Kt���I��bX�����}H�s���z��F"��:������K6s�k�^�?����גԶ�.Më03�
��B�'_M��N,�ujYM0ɱ<j�'B�SN��0�(z4��=yt��Gؤ�#��aG�󞳗>έx+.��ȯ ��@�\l�{���:g��{�U,iOw'��W���/' -�Si�2�����}��ڼYA�|,߁(�c�
������-����d`:��!�����7<#�yG�o��>đ��/�N������gƚ�pr��<�:��<l��j�	xz=Z���������z. ��i�=�MA����U�\����<�G"��Qp;��fi?29��}���C�S1�!�)&�~�X��}��ieJ������^5���}�Z3 N�����x���Ʉ�����A�b9�?Ɓ�_�-t�q�q�?��с��/4�?�X���GV*}�Z��`�I��)6%���	eN�y�Nv=�L�����&5ۑ4�jA��o�ɶ��<(?�g��#��A�}��U���`&a�K<a��G��D�1� $6K�|�<_`�_��,�;���]�ҕ|C�Q:XZ�V�u����&�í[�鍕ݽ I~b�Sn����h�>�#�����&��R�Ŏ����}×c�Q9.�ZU�2@�����p*��`jeja���u�hl�(��l��:I��@�.4�&��f�dP}W6����)���\�&r����Hs�U �oLfI�d��T�ʥ	��*�c���5��w������s(^!p�g���h��H^q�]( ���q7��1+��O}�n9��X�Wp�'O�6��01v4{����s�.���H,"d�R;�n�����`�1Ћ���җ$%�=In�l{��I�3����%1�`ԛړ��πe���_v�{��z��Pq�.~!���&����ǐ�y|�pU�Ԙm��p�I���Y~z�9Q�t�H�ёe[�!�T%�	���DYo��ր�'Ȱ��Z��c�Ⱦ޶�TtP��R����Z�����x0�;�E�:@���8�Q{�MX��]�HK�8�ur�p@;gı{ b�F�B��<��5Y~|���z��_�n��=W�Ƥ�o�2��z�?�W)�w���25R-�l!.�_�CGNVh��	�F/o�7$N��l��هZ�J��Lr�Y�/N�����p���?x�}4�syu7������1?�Ÿɢ֏mp�~~�>0��D�����o���������B�-udT������*C���.VAd��/ၩ[ȓ1�b��������Մ�|^��h�$�A�dqM{��JIE#�:�%���F��^doB�<J�msG���K���*&;�M2�`���&�ay�r��^��B��$Fa2v��Gu[���"����gY!�x���'M	�z�B���F&�>�q-��PI93n��Q�A"��V�z�E�eN[�n�����! 5�~3���'�� �
�ě~ǃƖ�\���e 	%c��/7�����}�Xx���j����s���9N�hb�]��:�<r#'�H��zJ�1%�b�t�!E�SwQF@er(c���oɦl���%��X��~�gtp���uw���!K�F�l��wgk�E�^�́d��D��1T�C/`V�x��8�(0�u���x��W����Ej\C�z���BXwe�����S|2>rc����Ҏ����{���ĸ�c�͵�;�u�L�G�a)�,��ga	E���F�rv�x�0M�������HR��e�0�>)5�F���{�[(�a�^W,% ڃ��YR��wU>��ی\��Q:��г5���@���Իwv��V8�}�{g�|�&�6��|�+�[ �G�ww�(K��~4����ˌRV��3i���#w��E�L��<��-u�����]�ԃ >��<�(��x��騔��0�ځ	:�����i��ю y�`tf�Ұ�n��(�	r8�(S�q�M���	�$bX��x/	����q�UЧ*��[� ,`��c0bP1����F�9��TY}��ڿ_D&R:�"���$��-��V`�����CV�Z&�qܾm/�c��Wq�B(��V������j��$��2�{��	šSТL;!H	
�#�X1N]Ώ�������w�O�h�����zpNqm��ڐ���υQK�N�QY���^P�^��x��dǒt����^�Uv9g��<��C��߷pƙ�ybc�e�ؽ����r>'�[��B��h��/���¼j����L�=�VfN��ެr��(��w�d� ߖ���N������P+���|�<��.=丏���1K�;=����	�����Z4xZ��)C���w=r�6�SX�"�1*�[
��v�����v
<��Hg�s��|(f.mv��4z�0�����K<�M䷪�.��`ǝ	g e,���P!�;��g�h��hnX���[{�k�l.S�4�,��f�rȟoG�Y�"�&Yb��T�{�����N���t{�R7�p�|*̀.��g�r�'#Bivű��DiS�C|Ґgq=+�ﰩ{9S�x���1���U���C���E�K��Y�:��B�d7��΂��Y/kwݓ�@h�o��P�1� Z/���p�*~�Y%,��[�"�!�l�in>g���k�SQ�?���ʭǌ�9�[���i�����;{�ª>'_�F�D2��P�覆0�%�sO5d,ɷ�s�٢�bS�V�K@�|	R�^xP+�u��H�A� d�,�� (��;ԓP�����uP�ww�k|Pv��`U$˳>/���N�]�Y�+�P`���%���>�06�iC�S�񶺹}���Nq������3��N)��h*����_\��M{�F�:3E�&�����1��q ��Kݨ���.(Uq(��N�=X�����#��� Z��9�K(��ئ��5�zJ�d�9M��L�"���}js,��=i8gά����+��i&�.��g�_*x�,�|�N���9��h�X�
�	��"s�ؚx@�BR9ӥ�%�;*}>]ن
F�r����|��;�~��g�ۢ������k��ih�ր�O�>0f�ʑ҅D��hǄ9��Z f_��@G�Ȥ��d��L[C�pH��{ٳ���v/�}ŹPwB��^���FI�oF^��d]f���
��v����&܆�)5��P`"?��bP|t���-e�Ɛc� ��^NjE�H��m�"gk3�;}#;�i���N�g�}�f�8GܷJU���,���q�?��:�HҮJ��̥zD��=��F�`�^��C�=T���]�<A��p�X�5�MgR�Ӥ���y8G3�6Z����D�ȷ�gη�@�iG��ly4�\�.�>k\Ћ��]*���V�D�Z����R�m#\�Tn�}�^-c�$�bَi`�h䇭S\墉;5 "������+�x[>�
�C!�®�x��(H��B�фз/�G��9�5��e-�߶v��wR%a�5�yUY�:�Jqm=Y���`��Ǆws�e�+�~�(\�Py�Z���k1�����i����p��R�K���v���[��r�l�^<��V �������8Z������M�����Q��䬲ʹy�R�X0��eet��G���9��&L��Y��w�zn���F��ZRmKІD�B�6��|�6	[7�V���M/��F}G�N0����ɶk�׷b�T�S�j��X;D�ι>��������֪�g�q���iL;���Uo�B�b�P�7�>cɆN�v�-9�=-�S!�$�o���*�.������Mw��\���n���@_x��%{H;�)K�ZU�,��o�U� p[S��iE�"R<�j�c}�����6F��&�K�́/H6_m�C�=&��Q��T}��bi־j��E�Rb��T���x�d�u�[fk�o�.�Á)T����Gy�� ~w_�`�07����j��
���]I4�*�ڏ�@��5��`����"C��K�4t9Iݪ�(ڇ�����v���-�j�����vf��1s@tk���Pv�J�<(%��4G�����J�i`l������w������QX?<�5:��Z��e�
y��pz�Ġ|)m����Hҩ�.&��������ṴѠԪ�]��J��tU�8�_�U��k̈́���������I����gRYɒ�r��(ph�5{��2x�e5H�Ϯ:= {ɣ/A�+�;������n<Ɛ$XU����o˚�S�-�;v�Y�U.p���{0���&v�v�d�^�O��w�t�gܨ`��@A���d��9tߦ��S͜ĝ�!��u]�f=e�#���	�9
�&R�B0u�������p���r���oH�6O*|�x���ԗ��[cr����:Z�Ͱ�7�c*�m��<Cݣδ"�H՚:��9��jƺ��+�9x��N�!�؉B�K��d0�x����F����w����`1 ��}u�ab� ��3|�L�#��_-�ˍ��](�
�|G�PfN�M��Q�T8\�9�m�f�M44����>���*o������̒�����&�4�4^U4��@y�}�/m��r���YS����F^�N:��7ݍ�[���<oP.
�o~)T2�D_1^�ds�f�²�$��o�b�&f�jiJ:��S1��)��he�"�;��5��V��9��m�![����E��g����N0�[�)*g������pJlA"A�mHv-�Դ�Z2������v۱|�?��ڈ8����w8�9�\���l�B��JE8��C�1Uz���9�L"�B@.��wY�2u�����O�~ ,���T��щs2���-@�^aSui)g��	H0�����/���e�Q��ᱴ�O�@�P�r���w >}Fo�i�g7��5�_�42�]�u�����
N�:P
6j`*
���,�P� �#���<)~FU�ͯ�>ڨ�i�N�V��?�8��EF�y��omY���Q7>Z%C���5��C�p��RC�7��(um7��3w�����_
���3����X���/�4/����c�l�dh����@?T�
�^_��&�WH4����ˡ4��[��}7QQ��Ĺ�S��.ϥO9����#Eĉ��'�R喅w\�i�k�B��q���k���v����|K�6�7~�US=�`�'x��1�/)�3+����2��*w�0�fx{�.���� JN/zl�c�����h��]W$Q�o���'�5�&�G�>R�������Z�.O:Pk��}nد/�����0���M^�^�ٯ���°�zz�"?u��knk�m)��~�ׇ4�J`������y�[@��0檵�\��s��(���:g8�[�J�*z��1,6��@���Pݥ�h����B��p.l� oK��2ˏ��G�?u�k�ێ�]�Өl�|t��'`^�`����c��4��E�ҡb��Ef��?r��hŇJ����Dq��:0cc�lV�F�rCl�H嘰^�THX�;-{a���A�t�����v���n{�
��E��ո�S'�a�Z̻��̈́��B]+��k	� 9�?�'%@m☸U=s�c4��z� Qx�*Z1s`�E�l�����8qI8�
4���)G�L�K� �1��]�U����-�Tt���������=i��ש#1��+xsJ%�: �9!��RG����GP&n-9^�(QUэ����k����k�HX�0b��İ@;���[B�-m�~����-x����?��B�owo�2���}��sN��6G��軸sfQ�>�[�:D��]T��$�����+�˞F@�Nǡ!:a�!,F�ϱ���۽ɢƉY��*jM���OvA�T��	�|�f�I���Ddh�@�:�fNKDSϼ��ZA�H��+�k����b�Wؘ9��mfeX-����m[v�­:`2k����^I�\8�E���� M[���f�>^�k��&2a���������%�ۖc�\ �i3JA�(�[^���}xV���j�$��p���@̅��`W�=.�2�E�%��ﮣ2}���&�7���U\��:��Y<x.�7�L���^�~���f+)�uUM���;�R�"�5�L��1����נ9j��1���&V� -�q���yDG����$�~�-��(�,��v��󳏱�<�#��p�ǙE���%&�����v��N��h" I����,G��;�9%հC�s��d)K�"�r�ȀUhx1�B�����=�.�׻a�x���AdUB=# sP�����o��1i�{ԇh�^�5�A;I��Die!>��f%'�_��g�8�+��eOk�^+bb�����L��a{���0$^���
�Q"�@�7��nt��_h�#�������sq��i��Y�f*�����B6yIq kD���Y6�^��c��:�nz�REաz�iL��el��51��Uw\�*�T���q460��ɥ�/K��p���Wk'?�Qm�n�{�'���u�2���b���8�_~�,�L/��W�_�{�����z�A!	�~^O�p�<�K��T�E�~�-�%�o�����f����������Ŧv�b���b0D����D���N�\����0vŐP���=�1:�0��x���⁉���I�'|9{$��9�SA�h�`�HX`0�|��v���˧IԔ>�_��Q�W��Z_����N֓�5r���Ou�Ns��k��q8���N�r�Y�7Z�<ߖ�ښ8S�Q4��
Cl�X��|�� �6������t�0P��Ń��p�Z�a�K;���+%��Y-��}ɶ�W���Û� �`�Љy�7,|��V�-�Ţ��s�#"�d�g1��t�O�1����P=h���O]",��e�\�Sp���.<��̢��R^�dS�ja�c�6��I���!̪�w0��ޥ�)��a�DF�@�P/Y�V�.���\��s�?���������c	k������[�<���U��ʔ8��_J�;7NT�[-CZ6��;�[�~C�$�����ERy���7E��pv}��|$�����I2 )gi/��G�0�ߥU��'x7���P�pAA��>t�Br�!f�v؍^� ��M�A|UL�0�a�����X42�E��k�ڱ~Lo�LBw61ő�/�> |����b��
s�����?����?���!�7��yطi���.W��p��$���'��3X�R�n#����Ye���Ӷ�x�N��T�&����
dĄ��_��r�5F�D�#�e��_FO�q7�Ӎ=&X�Q^��e���!���s4W�Y���]
����}~ �Yc�?cV���j��0�KLg��rGSt���y�C�şB���d]F�r��->.�6\����D�"y���/$�]^9k��y�s��`+F�y0��K3��vZ��b�l����Iax ���c�&��*�A�@W3���jWŴ���������B`Ө�\u�.L^?�Bg7	F��T��e�e�����Jۂ��1�`��Ǥ!��8�4'�þ�c���~@KɽcD4�S���
;�54��BG��m��B��Ag���3�<t�~��i��@p������6ƙt�S�eS4�A�$,Q���<��v����ŧ���"��'� �}%���ʝ�@�W|�����ey5��&�&9Wo�����r%SwY`)�����s����B� �&�O����wY�|��U�H����Op����l�jDJ����H�@Ʃ�FQ��rZ*���B��W�t>�M�`?v�]Q;r�u4>�L5F��0�Mk�Ρ�,)��U����g��/��E��ZC�W}����w��tO-�2�����	�HBFT��Nأ%UCW;�<�l��PW§a{��_�h�k��a�B��+�C������\�p3�����Ĝ��両����\8���Ih�oД��N����� 0Pq��i��RvHsLÂ��ɵ�!��h{D�W�(���o�t3�2���b���?7��A��!�Q�U�SK]׃��L�/:��'��]�8T��_
�ڨ��	���n�'��sa�P��1�e���4i�����U��<7;��l��"���ѭsss�2L🖛��y 7��e�J�����R�jU��A@>���T�/�t��f3,K�ʈ=ǯ�<`쮵����Ɨ��}m���^si(as)�Zn�X�_�+�t��V��ߺ�$E���Չ�V(���,!/W)Ǽ����$e��"Y~��Jeg0��<�
��|*n�a�\M�1'���W:@�k	8rot[�3��ij'�ٮ@�#G"�K���d�"N6r�*����#�n�ebo��
c����qL��-uB��L���H���#!�!��픲w��c*"�����u�U�ܼ}'�ж�V�,�̓$�=Vz��Btf�v�a��W�B��{��O�N&9
��P��k�%Ϗ���vv8�gY��r�h�(Sz�M4oIQ|^(y����"(������_ŉ�\m�\�N�xd]qw�����"�Ӷ)�� ���3{��kΏ�����x��9���mJ�h9kK`cWmOx��l���!VK�[��a`�XW�p|^�_H�b�$�������c_)(pm�E^vj�[q��-(r�<�H�ڕ*�:���G<LAH�6|x��^K҈
�~�ܝ#9Ő%�_�e�a�N0	BX]���U�M��=W	=�e&}��<���A��U���7�ϰ�i6<���15lmy�";�MknV����O���0p�ҬתIN��^k����K�IV[����B!9�Z��S��HN�/Mq�K���c���
 �h@��V�����qW�v8��o��Ξ�7��
k���z��c�z����7�(i]C��$YdB����/�����:���n�ތ�q�����83�l��	˃�-�4�VcTi�Z�=c����?84�k�pP%�a �Y����ID�������������i�LS��o�����/�����e��E��w�hH��5g�޴uЋO�U�������'��ypkb+-�M��S���
�E15�W	R���y��g����	8��,x�L�m��D�� m<*��=VH�v����07�rY��$�"�M$�]@�k-��Q^*+Q��Zw��djٗ�3Rt����sY�B$���G
vSZ�=q�2i��ZgVJ�?��^^ɶ�J�PL�"5��§��.B��%��@����@�\on����Iu�������n2K��7�Ӿ;�b�}L�q��T6D��\���s\aޯV�AΧ��ó�l����>>�;�jF��^29�W-����&�����YK���\nf��N�i��"ꡆd KF?]0�֯T$��&Ғx�W�OAv^�Fxg����~��2! ]���˺}�C��2�D UjIh �q�V �fϿ�e���)��� ��Rz?�����v���[_8�p�0�߀WA���Y2kL��}��~�Wǫ���p+���r�4y.�^["�__UB_��9�5���r����N� µX5
&�(����a-�$��.�74|J�yrΜ���#���x�}
�S�C��/pp�૶�c/��Q8����'�)Z*��	��C�B̭���������"X� ;oD7�H����/�X�e�x���B!@�:�k�ӻ������<���W��r���	�a���*��6�Q�}T�)�'��o��z0
L����!��L����:����K@wH d���X�F�zP�J���u�JbE-�K�v��
��(ϰLcx�>q��7���w��������n1<p�1`���|��r����`N���v�$����W~��t�-H����aU.�{u����tR���J��S�������"
1����ZrCT����ܫ3Ѯ��4 �����(�Π:*��\�TV7����3-��@#'�H�N�2!��g�e���F�F�(�R+[1����m!gK�:��� ��J�}C�r=��|��XvGZ�8U�f\<$�Y�~�m���
$��-�ڤ���ʆ_�YӀ/�w�TܣC�`�s�K�$0��˽��%A!Q,]�t;���m\�Jv���14��@Z��F�/ eQ����z�gX{��Q6�]�)�7�q�Q
(2f�W�*�biRηB��t����ߏ����ޗ��7��ܶ����2Sk`(a7���`}]l`yq�:G_G3������fz=]r�Yr!⮬>�ʞ��©t(f�w-Q:lm�7	��_���B49��7�J�9�����A֧�[]=�ʞ���%I�ѿ^�wy�"%|gї͵>��$I�Q�&�B�X�#x�,S��7m��8ּ"�l*���8 ���3�����+rH�p���a�Ũ�Vr�7Do*�����%���Bu�Pèq!$*���Z%Ys����Q6c½����4qU��l���%h��bV:�]�0�Dr��{����RX_�!ü�j,����Ȏ���9A� �o?�s+�ő�P�9�[�JѼ�Ytٞ����$�K���W[�[ߕ��Rt'����F�7��N롺�5� [=٭5���&���s���j�LW����7Ʊ�O���|��0��"��J�\�|#Y�0Q?�%�Jqq�mo�#+Lm�&���^v�c�Č�ɬ}��<m���F\�G��e��>��eSēW�R�K�V!D��Z��nE��������,���| 
4����$�1���b�m�.��c1�)ּ�ͦ�����%A�]{h�9�þWz:8�����'u{�m�ֽR:Ptn<fXT2���V?��|fz<�u~h�
�D�d��d�D�DPE���y��[�-��ɹ���v-࿁&�~�m�2����s�4�Ҽ�ͦ�6؈9����>�Lxy�c��ڿ'� Lch-�ج)� ӵ_O�P,`bī�>�d�KS"^�o����Lr4��� �	�cyş@���ŀ����ؗ�����]BFBG�M�m��=�^���р~�sj�B>�����iZ�BQ��K=�y�r���}A�s�>��S(�^�a0�򏪃���[����4��X�!|����,Bݨ*ӹv��Τ�vW���S�(MP˝N'�]�F��e�f�0��I��XiH0�m���IW�'�M����_gS�Ą�_J%D[-��G`/]1y�(�o#@��:��X{ڿ5��pPҞQ��i��<�i��Yî�U1��ҟ+;�)�6��&��K�8�z��#-a<)�d#߫���t�UD"���c����zH�%j���~�����T���)�$�a�uL�[�������㏓�r�s�����z�?N����Y��=�f��e8nCJ�� ɲzt�D�ŗɑ�3��m}-2	�v�TW�(�A��{�v:�9 Ψ����"�b%�[?��3`>���4�,�)�)��-Ân��?F�f��=� d5�)U��Z-�)��4���ἦ��c2����bά�_�Kf��u����T��5@��r[lrz��3L��xN8�Mx؎h3â�S�:=��H�M���䞂�5�_�]M��q:?8a���\�$�h9H������p �T�'�)=&��YV�g��	�g�c���@�r��Ŋ�v�=x�<�������{W�����qbB���Ձ��5�o��]�|P ��q/�l���6�^��EjuofW������ѹ���paG����?ߎ����_�#GNjU{�5ğ���l���M��WQ��0z��'N�۷�����c��$iIk�t�F*I"<�����jLے�e(8ͪ��M1f�Z��2]�BR	(d�=���bX��@CH�}��j%4�B�L@S�=K�3sA[
���З���[&�X|O���{��]�v*+���c&�]Y����!;�3h1g����{�lj�����N�/���������<A��g��K�}��6�"�6QYH���u���I��n�"���eb�-ߗ���3q5<��R�Ζ���mp	�m����k&Z�w^w�8�-���<�p#��2�LEǹ�i�����j�2� +���.D�����H���\B�|+95:��ǆ#�)�k-�|W�p��}�.K��РN�oڭ���/ �@�ND��f����|�"���ʻ�/��u�CUIy��֎��uQֺN�*iÿMf�;.���,F�}�-���7��F޻P3N%R� r"�.�n/�Sr/�0�ɓB�G�}�⦭XGW6�f>|
X�~q��X��ꇊ�Ҫj��X*�����.�!ZIF�6e�M�����z� $��\���������/�&� I��|T��7�o=��� ��U�T<by�+��6��wtզ=&4xE���V�af�ފ�Ux�qn+��������2},�WENɉ����Pb�:�W80~S9-����ܶ���#(v͡g�m��1�iTR`��'蹕�����Z
qn�:����oIC����p?ϊ�U�࿪�:M���=G��'��YI6�h�:��Hv��|��)��o�P�+����;�m��c�̮��qs���˰�9��?��on�;����P9p@o�8i�΅bHl�FHu`
�QOj��_�WTT{�۴;�=�[�\s���^�d�񗗌`Y��&�C� *iC�nF����!@�v@��\�u�����/N�E����?�g���60�����}��u���D�m���ZX��V��q�՟��"̣4�`ͥ@�ߚ�d�<o��i$���N����'+���2 [f�R!���� 7Vr^�-Q�^���ES*D��>+��{���zӖxU������P�4s���P1�q�Ox@Կ�̮p�H��|)P�����c�&H�p��|���6��������x�6q���Ҥ�q��n���yW�����(mW���f��_��&�_��QH�8�m��°��D2���$����%Aw*������ף��UN�斞������)�.�8�C�S�Ľ3G��HH݃��A�B�s�>��֍O<׈?0|+_�݃�����^I8$�{���lA���p͹�}}�����a�0�Nr���AװYdKd�Q�qP�?�^��"1��M��)cQ�dU/P�+�cH^�R�@�i�'ЌX�P³D��Έ��>0ޱsR��DYa\D�t_s�4<607��0��-�g�����5�/�Fh�" �D#�~H�y7����(m
؇ß�N(#_���\goS�2�r����gǈ�CgUw�-Uv"̦�������Ζ�+�
���j�n�ë���TK��i�O���C��C���2v�7u�q�������0��Yq/^��+a��TQ�dT�?F�?s~pJ��t:ԓ8~��A)w s�����$���4���숷;,�?T;#��T@uh���OI�HJj�X���LlX�)�uh���c'#1�:�OF2�1AbY>_Zxltfq]&
�e���gH*ᵛ�T���R��m!%We�r�]0*���.^��Qi�Z�"e��:�Ř1`Y������s���	�D'�vАj:���q?��57|�?2�R\;
��\Qs&��~��{�a��#��J�����>�����	.Z������"��s�{��Z�`����hH�앚�}�/��9��R�������UT�h���3
��pd��U"A`�C6�%���{`�I���K��SJ5�~[UA)�ri�N��#L*��_Bd%��(�Ҵ��r ���c���h��K֣RM2QyAK+�/�O�#�b�/��J5��۟V7��������Y�i���`��l��O�B�$9�Ü��ȸ.\9�a�[��h��-�ϮQ-�?�tJ9Ĩ�).3Oq�O���`���=�qK��Z��gy��Rb��p�ǀxae�ء �`�~j��=����ۻC�n+���/�_5���;�U!��D9PR.��#�hx�Q�UPhn��x
�)W�, �L���& �:�ўI0��K��=�$|�*Hc�;ȿ�����A`�2�����.�ENo���ZW�D�����֗�)��4׹�%��C.�6Fd��ن�[l�(>.{d͡�k�,��Y�$W{�_ɹ!n6��蛟ð�$	t����j�_y1�eK@����C�9HDd-;�m$���l�sN�bǌ"��D"���c�����L���y�}����粽����b?�$��3��sG�W>�����������%���[�?�~*���A%��:$i"�eɊ1v������b�\�?�Bn2��`5�ڭ�4.&6 Qkʲ�x�UEx�eI��	G�s׻�,��6�l� a�+��Qǻr��4%�)����La#Fڠ��w���u��(#�Q���<1gv��48D[pޝ��VH�-A�	����KL�׸�K"�6G�ź����=q�
{-t�ul1)�-J]��h�p�=��kS|V��`��4�St	���k��;!��_���Bm�o��Nw�D5.�DH�g�����7�>�e�$������ɞ��B{�y��
�S���&�_S��s'��m�G�D_t�/t�F�S�1������@�Ӥ�cqB7GH.�9	�Cy��� b��.�]�����F]%*���η򻧑�Fo;�]ۙ���������-�<|�vBj�6e�~��t-^+ݬ�ݷ����39Y�j��_��N]�x҂�L�EVqp�Tj��\-�ښ�J$�5��v1V���|Lqj֕~v]�{�ΰ��JiX��yPr�I:<8����8�TI�|�c�L=��[�X�|.�Bޱ�T�\���M0"������Ɣb�1ʚ��P�?���mz�{��A_Z�S��{�G��`� �k��ֳy><�%�����t�/�(7�.l'��Y���.�+)�+(z�_��NM-�,x��n���w�Qd@�J�����h������:�0Y�{�EN0���@��]��cR	ZV�C�0��g�P�f8l�5���X:�7Yl���_�`k�����~�rb�8N0����1T����(9���|MKZ���ƈ*�'�kW�։��U��%���=a\����L ��~5���~`��xp�ǐ��	������y5t�U�ɵ�ژU��g#�6O��9�] �Gq�K��x<-
Z�B�/���b����C�V�d�ے����:G���w�MKL�X:���u�c3}�ri:&f)�rTQ���=D�.4w���F�6Sc�������d�n�y��>ﳦ$�������ټj �ޣwU�^�o/���'��R�����X�-��_�h�~��o�z�A;�%�՝��"�)��ǯ��3[k<�~��!4F3R����;X��v��Bg[$÷�OF�,G��4E��|�|x�]��L�q�x��E~���Yt��O�KU�qBR�p�ۅ���ͧ'A�I�ŋ%��p�:�1�VM�P>�xi-4��)X����8����{l�6�L�,y�G�_L�ٳ�O�?�] ck���_Y��Rr	��h�� �"W�)���������Du�Z�=�z��l�n����%5����>	��B��H��~�ы*��K���4����/i^�f�)�4�K;nz�V�:� 3_6_�m6y�T�?_��I��ß߬��Z8��;'�����-+��,�o���!�<{�r$%�?R�*a4�໪�Ǒ�@ۚ��tR�%��/#�au��H�V;�����rZX�\p��Y�$���Z.�]r��W�s=�?SIвS��T�3�?���_yD�I]oJ,v�H]H|�ڄ/��앀̼����iym�K�!6��<=�|ʸ��\�� �x-E��!m�;�����Z�GC��5j>��9���iU;s6�a�����e���팝�@�������Ճл�E����+����kJ�����»��A�:�
KZ�Д�*3�@I���II��$���3����קQy����5��*g��G�!����C��3��d3qEft�mE9a�{��3��?�$�p�]�R��~O�n���].���c�6�d"ͷ5����L9Q����)%Q|��x,4�i�����L�A˪Y$!��I#0��/�x�ֆJ��O,#H~�ah?г���	��:�2�[?c�ק}@H�\#6l��0����2�V���fVm��g7���,>Yk�e�?]�I��W?:NЖ�w�7�4�Td�h�z��n�]��?���6��P "�O�}1Anw-�"�ҍ	H���H�����n�xXH2�����i^B�w����Р���xO�`�����xq��
|�Ԟ'~�u���YA�H1�`�pS,����$�Q�� D~���n��K���Xf�1.8�2�e5�X�Q S��A���c�^��ٱk�	4����c��}���(���Pom.���xOL��{5�&��m
�h�����Г�&���!�O�T,��nBt4B�����|��0�{T���'����1��{o�ɮ�67aH��}���x�q]U�W���}Q�RA}f	-Q�vԳ�&j-��g~�oD|p_+�y�����V�b�m��9oml�ljzVP �1�{S�5׮­$Q�6G�Y��o��4�аɑ�.L��v�d`�OF(e[%�:Qu�|r'�A�_k��:���F��^��ٞI�jB�96,�d���&�RP�Dn��A�?�O�#p���@��yW�I�s �s]�oo�@JA!�ĴPOZ�3\�T/"����q��>�\�t��H���b�12Ni/1R��mD�8��˧�w��94�S���:>1�c�"��d���R��m?��3�'Zf,|N$����؏G��f<Z�0���/��	
W�����Lc��d�E��^�e
B��#~k������� ��-��e���ʙ0^������
6ܑ�m�M�#S�tR�������s6l'�·��1_"���笘m�����������SS7�1���\t5���9!��O�2�T���(#*��w��񟱜�-�Q�׌��U[ړ�|^B�7 "x+�uf����Vm�dO>,ܯW;�6�C��������Z�,A�I����wm'�X�2|j��v�d�Ե\yD���p����Pʍ�l�����CO�X-#|?��Tu���O��s��?�#�,�׳�#��F"M�%I����#����@TVÊ�S�@�o�y��u����{cGZ�R�K�37�&�2�!���C_R%��o����Q�w=�ӦN��{�E_�G'G�`��Z^��pt FIz��"�fn Fs�Ab�Z$�� $e����9�,�w��i�����tT_�l��.�y�v���1hZZ���������}� l�}�X3
�3�ɛ����-�1��`�0��upHU��v'���]� :'Z)=�@v�3���E���J�6k>]㡅�K/* ��Jy�^�*N	p8H��$wĘ�����`������e%��V���u♈X�A����eL�hAU��V`���W��(Gk�.��_y�x[X�����05кY��Wց���D�~6uۖ8En�&���J�������b��Ql.�wɘ�&veql�C��[�"��"�I�2�6$��t[��w��m�l�7Gj��\��f黧���k�/��\_�}.v���o3�9vc��Gnb:p��Z����0�2��`��q+	�g-��_A{2�;����׏��Pɟ�����%�C�|���}ݳ��>=_��؞Q�d����y�b�(�&�[F�@�Yb��`ZM�n�3��	G��M+_T���a��}v�V�ݓ&"�'��
R�(+~��S���G��Ф�\���/ڈ��D��KB��A.��J����h��_M��}�3 �G�������{q8Ar˥ӐoD\��;MP	�N��L�%��9��>�i'�ʤ��%���=@~�㿶.�?o>>aip��k!�:��4:�?U�J�ȶ�>�{^0P\�*Pj!4w]����=*��#����.Зs���Ѥ� �Z�/Q��$���Q+x�ʄCľ>ȵ�ny�ϻ�[�nyJk�������aJ�̥��ΈBbF�?禢�ZgJ>��Vr�y�Fj_D1.�	���&:aڧ����.�Q�P�Hm
Q%���2�x-1Qg�4��⣹�cO��)����,�:�h��)`�x>{�RE/���G<�k���gwU�9Tt*Z��m	
����Iˣ��=Y��'�Ov_H� \5*������c�	~ {T���U̵���>��W�3�
룘�C��v]iҬ����E4ؙh�;��E�ɶz�Y�k�c?�N,\���1n�6d�`q�N,��z�����ghT������#o���`������������s��h��+��$V�����Mb�J�}1o��#�q	��f�F�Ė�3���Kĉօ�p�Rb����t:�������J�n��"�p̞0������ �PҎ� 3���8��5|I�E���x ����1]j"=X�S��T�sF�;&�Ѯ��ul�?6��Y��q#� L�-۔T��(�����HG��WT��,�_�-�i$�.kp\@�J��r֗_�@��~|��֥��:���wN1o�kiBz]'s�/�3=j��M��MrL�P�U;Os��2���]����^p|3A�r� 1h��m�"���} ���ވ�ѕ��J��a����ȕp��d�ʿ�����~A�b|�AF
�T6fT\;��neh.�}��&�ښ��NȚ��k ��묌Ø-T��#j����r��PW��ý�_f��x����.?梾oDe�+������s�������:�k�L�O��z��1������'( �d�*�o`���z֓xx���	R���$]�X�@�D DI���=$��PI?�֙���'&�76���d��f��U��>�K��=�p(X�ux�?�u�X�2����8\!�@Ş-�ͣ�/~�7��(ЁS �z>�<�u �g��(զ]f�ع~��=V�R�k��q��t�ב��&y�i�Z�%�q�)�pC�I���E�v(��\P�C)��澦�$%�kB�vb�"D
.�:ү��5�B���)��:�Y��x�4:4B��'$	��F���}do&�Xj���r��ĆT����� f�#1˚K�5��/6�k|�ڔv�~)w}����TN.F�����3Yl�^b�Y���w�tQg�hx8��G����b�tK�@�Ww�#]lE<���;�-�8�O�#����@�2�������F&��t��N�|B@����7{�N:�h�,J���#�Ӛ���y��5R��=��k���u��&��f*E��҆���B+��|�v3�l&�E��!�Ğʅ�d�{K�S�[G3���}	�T��¨£��y2ž?�x���_����x4��MS)f<�9e��0��I��?�kh�gG   �4���d*��)+u��ל�\�8�c��κ�SGa}�K�����Dh�� �J�=��3�7�Y�J h����?�`��LAPJ�U".7��pD��^����Qp�Ҏ��3���E��-��=hd�����*9���x�sD���Gt��ͪ�N�2� *7�#�����Q���C
��|�8`�/�;yk�c�'B��A�}�����ߣ�zGt.��W�����#f���6ܒ넇9�5�H�]��7u?�U����m+�Y@�%.�`���j8h��ȡ������$؉I�	۹���T(gtM�n9w�U6�yx�(Hl���d�)B����lM�^�o�/0��g���P���������r�1L^9Sī��u���T�ϗ̫	dΰ'�C����,sn��i�ԣ4����o�|cU�c��}��ʡX���x���#��.9��?����� g��Jn�Z
�c`W>Wm�(���H��}�� B~�[o�we����|X�_U`d��O߹5I��dN�|��������$6&=�P8�� ï�4ͮK�`͖��7����t�e�Vת�X�.�����]Ӏ����C^>�׋E�'`L)�T�_>�+R��T�m�<�ԯ��40��=� [�*�G #��&,���iކ�����U��^���KiL��6�>0�1�hO��'�ڼ W�����<7��1��Z��I�|����Z>��7�͡��RIo�H���z{�/��h�� 
z2��YLx>J<�z���r�^�_I<��j�\ ��eQn+��E��=�	�5�h.�a�e�
;=��w2��p|�1�3nm�]n)��|�����&z΁Mr�sz5�������'���p:1����&������̺Bd����}\�յ7V�K��ƺ�4���?),��/��\�ߺ��������K������r�Z>�3�s�yd��Wx�ĸ!�d!u/�%J\^Gl ��ӱ^���������U0Eaڈfs>��a-2���o�y���c�w�Skұ���龢fj��L�n��[m
��[#%�ޙ���r�:M���孥��$O�%���`x1=Z��#YN��~�[�wA�}X�d[��i���������#�EyL� Y���=2���+��s�V���gC)Z�*��6�#�,��~�~Q`��v���dڱ�b��;]��z���e	T��k.�P!���n�ja��Pk�>��,��+�A�V�'Q��g��$�d�o]r�v�������p֖��	U.ݦY���^�hڣk�u/$�	+�0�ӎ/�{��M6���g���
Bx��Cm�7i�X��U�?��I���$�E�:ɮ�1�:`#?�G"�:��M�@��3Y�%e�yp"�S���O��^2P��Y2�mr���i���PWv�e[��i�M乚�q�T������D.P�0Uv�'M�Z�s�=�%�ت.�@ �ɀ�E�A4 2�~T�xQr�+�
ܮ�p�m��σ�>��4���|�[@x5���}�՚�.�T�]�+Cr���/ӱ��3�/�4 V�?�Ӆ_��VX�������5n���Z\�B�P���%|��u�L�db���4��q�Η3Ze��h�%���)\�,�ܹ¥tN��NlT��U臅�c���J�d6k���p��dr2�pe����C�4�3N�$�[=�Ԍl��)~������R�3�/����nZz�)����-jZ�4)I�c�|���gs�:�SH���~�p�U�����q��$cm���.�P�@���f�ڧ�^Ò�zb��h��Զ�� i�T�~ӵ��[o�&�V���ìfrI1����O|���L<�2���A\7a>�����&p�
o��!X���o�x�ݭ�A��I�FJ�"��z��l��(fM?����m܌�M�`��%����O
*�PDf������<�#uT �ԛT�޲0�1�	���\'|骍v�xKO���yR�4:�t3���}� �ŝy�	�\Y�4W2�l-��O>�I)ȴ�EI��784�+�Ȁ���ia��K#���,�R,�X����x$����a�`%P�?Xᠥz���@6o���r.��6^��ϯ�s��*�T�c�V�fAx��J�\Xd�YH塏�P���K�C���D���5�q��6pd@����C�n�ҼO�S);���n��^��(��f�.uj��#-A~�&�-ģ�|����bF�
�&m�lz�sG9E�.���Xlj���"�����]A%��[�+��G��KU�UYEڏ�C��G��V�/"��Q���q�~���U2	c&z�ä�KS�%�����9��Ȟ-���Bj w�\���#�[�6sYS���s���:q���f�sqrA�T���L�TUۡ!��5e��������W�7K=Tǒ�����5&4��t��:u�$�:F�D����|+-�m��֋����?�镡Uue�V�;=(č�`ɷ�5BQ�B<Rh��עޣ��ƅ�o}/G�!���y������]e��q��7O��3��8'���f5&�j2�ժ��j�[-���'�Q���RO����Q\��4�y�-��3���Ǧ誮g vw�I<��z�k�ݨ�����7C�\��Ѷ�UQ`�6��`R�������X;�xo�B">����O�&�G&��A�! gg�3~� �d.�N��I�����xY��@DT�cLdi���Q��FX��3j��> Ft�Z=����o*&�Bm7v�!TQ5�+�<�Xc��?c�a����F���dǞg+��5|ߙ��dc3��}�7�U�UPQ�ܿ��%昀�Y �eN!e)��]��y��W �Xe!#��.�<��� G?��^,���� �����:������wg�-	@|�2��|�F���:�� 4M}D?_)�F��b�v��"Q��Y�6k����FVQ�,�Bj5Er�����2n���F�̡�O{�tu�F�o����rdo��xWH���BB��U2�]a���_�a�Ci�V�9�q���՜ۘ0�p���؛��`3忲L�Z;M;�����P�#��t$ђ�� 㗧N8Ļ��S8��87S�3u�Sm�f�Y޴���B;MM�T�>��Q�	���bJ#�?�p�V:\�5r��������Ų�,�Ĥ뀏H����������xN�]�x(�+��[���o(��bq��RjiTᚄ�B�?��̱m*A��0טO���^�e�͜������$���s�@MF|,=�\���������Y����s`�Z����e;�u�'��?RJJ#��
��F��pS/�-�V�?v��_�m�Τ'�UI�����!ڶ��&3d��ێk�9�3�ﵡ@F���H�x�/벞�q$f��սf�������b��C'�k�R"c�o�@���=˛����]��U�r��	fY׌m�J�]:,�Q`�"�{ܫ�M��#��1T�qgw["��H� Рo�HQ��[g6�O��<A�Ҷ������-�g�c������9�������d�o��&8Rע�Z�3�'u7da�� k�H��a�Z��S�(9i����r��[������,������>�k'!תi~J dO����l)�ELhʚ~�Ȝ&uR��{�ȿ(#�D�Z���XA����ߎ�\0F���`�J�y�P�Y�`p���U]<�׳D�{h[�kEu��nqE�Co Q��;�qQ�-���i�|����Y�,}E�"���)zޅDL�w��F�t��[�[j@9�YS�'}i��J[[�_��*�9�U��>�1ÛU�z����I�El	��j�,�6�%g���=a�.�������@B.t�EZ�.>�:�I�!xF��ю���v����Z�ؔ�����1r�EH4[��
��I8CP���xc��>�[���t�RNi�΀N��g�`��'d/�9`�g���]�_�[�?��൤1Tg����،�z��S�����5�b�W�XC���E矝��/�������@|���t}RUأz`�3*y�q9��W3-�}k�	�۪�|�8i��&�G��?��s�Os[xi���Ԅ}�Z(�i�����%���=�7�禹354 ���8�FvqϹ5�T��G� �>��J�^�*;a��ȱ�-��C9L���1�KF�-Oзui]��i!�1Բlu=\B�׫>��A�Q���������3(ﾼ��H�&�$��w1�[�Uf�.��4`� ��G�]�z��0��Ab��ּ�����_j�*ɻQS���YkI^o�A��F�6�ǐ$ń g�{�m�Tq���{s�K�(A-�Ͼ����N��^�ls:��0����_��[��i�נ%z����f�x-���vBx��	��nDX4`�(��"�nwv��%���-�Y����k[�b�'C<�Q�S���K��h|HK���c�1+K���Z���O�D���*6W��ב��7.���!"�~ ܯ#a�Q���i�"���oBv�~o�U���B!͢}��F'U����j	���7�H�`�b��6�ӌrZ���l�u�JvFC`P���I���	F�WX/W�a�K�n�xm:D���l���}ɐ=`�ΐə�y�ȉ^'���u��*��Ӏ�ѩ�
���$� �� �)�
v��-�H���RL�~oS�E��z��ܨb�L�
y��"���()����
�����՝�L�����ڦ���0�V�r �"�+t91��
���`3zi�Al�S����fu�n����x�F��h�EPg,rj.��
�sWܜ>�8�<y�}E�F�q���f�]2H�ݓ�D1DN�Sy$Q���|�d��^��9���	v#�a��T�_����+!��hn���)�i���M5����Xo���3��n}�Ǧ�E0�d�'�p��-�KJz$�nΚ.�a'^@8B{����i�w���ۄjK2�I��y$#�!���_W��g��+���T�o�	Đ^Zr�TN�K후L�r��ɘ���B'�����i[:�&�~�^��;�;�����*YG�"��uL"6�t��m�l9
�o,y0d���A�A�F4�.1,m'.�H���:葁��?�o(׸`��?&�.6�����k��\�=_5��U�p�>xv���y�,X�XG����d{��j�ϰ����$C�ANTZ�q�g19�D�[/��=�ɴ�\���k{f�@�n_��A>�Ї��`�A+�B�����k����W������{�����ʪ��ʣ���٬*(rcd�a�X���U@�0�|�X�7Ìi:{u)\�y;{"2ҘJ:�v���;F`i��%q4S��U����z�h\������<��T9��c�\�����h(L	�t9�bU:�S[ti�?�O} �<eǍ��L�/�߳��!+{�| �*<Hy\���p���X�J����~�N� Y�
<�Z],��(w�B��I�t�S��C[+�4���
�޽���ޣ'��m@����2��A3��7PR����'��%r����X�ɗϫ̏M+�Ć䆉=��l��Y[S���R�4�.�* �?�d^���Ԯo��G��d~�<dh豹�
��~,��j�c�Qeb/��Y��eC�A78���%�V%�l����{�oWЂ��%�~����]�}Aן��9���o��f^�B>�FF��K�;�(�-�(�<��9u�R���N��&����ı�B����gbid?����/u'l r���#2�X��@(�\Y4��G���ȫN�Luߍ��&�y6@�i�K�fH���5r� � �FM�`a�>���+%8(��)���g6Zb�����q���(�ݸ��Yުq�ڥ�+�8����RT��Z�\_G�D�W�'�k�Ke��޽�</�l�:���S��ч��b�HC�P����㻓�2��*�<�C~vM�$��Y�*��<{��tC���y�*���Ŷ��gϤE���v������✯���d�J�r���(�;t��t	A�/�E#x_H�9^����I��Dk�U]�E�-ss��ORq�.���~�T���]%�"yr��<�iZ~:ʈ��\:^���c�x�@��zh<d`�=��z{���d�Z�V�|��@d2�7s8�;@�޲�� >��+��m��Y�E�^���9P��YM�4�����2p�02��ۨ�Qr�^<���F�3�l��"��*��F��t�B��[�9)^�
�k�:��L��W^�T��}T>\������}�-k�%�]�-q/�/��	�X`�����t��V��)�vC��~���>��@��v�/ě������{B��8dV�5){ׁ=gO�H�쟹�^`�c��ǲ7W��dͺ����	e�y��0�o��'��EsĽn�5v���N�	�HpST�`W�����*�?@ffj�Οp%Ɲ@~ۖ�y`�1ș��\�7�Y8I(��>��ۦ���6�b7�D;X�	'Ĺ�l���'��}����m�G��0��a�����nkJ�,�I��N��D�~�."g����sD1~�o��3�m�aK�6���9W��*���|��)�uE�3���_M*�$!�r��^m{ޜ@�dA������4T�i����5_Ŗ	�ﱘx���[a�6��>0*k��w�G�G�b[#�ʹ��,��
"2�Nʜ� 2+��� ��A/�a�,���ȦwTAEE��V<:@�..���e�OM�ʩ9��v����6����
�*EX	ۥ�l�y�G���U"�89[{�rh��Nt��Tt�8����I����cѢ#M5_S ieXm�;vY2�~\�
޳$�>�~;5��H���f��ҫ��"�/�j'����m����������@��p� �NH/2�Y�o�1��I7[���E0���{�ڿ+�ݨ���
A���ȓHݠ.Cx�R�^�3~�Ȥ���a�4�s��o�2�
.� (aw�O�.sm����'������ދ�����a��9�eY$�J^e���	N�KC�xan�/\�Y1&٧���F�9liFR��jG�!�A;���C���#��B�!]�BP���v8}�֟���Ԉ�a#j`�ͻX�
��?�d�#�je#�_23i���D���O���V�o5D	:p�ͦ��Vv�l"�8�^�'��]K$3��w���h�Ё�<�k,z�W|�u�p�8��L�I���1�b���p�7���O�av��.����������ؖ�j����
�PA)�_��V�I���5��;[[�;���w�wy���J��d�������Se�a����f�����3�R�A�ɳ?}M>Y��<����K�����-�>��m4�9tI��\�?"s��������4�S��x�䠖~��e:R����2��i����dݳTJ��F/�ީ�	���TG���j�O�jE�<�kS7Ց'�|����	��:�#hL7�����/��h\���u{Bz$F������vK)���yé�r����x���tU�Ov��(�ma����j���S��ӆ#����%�����L>s�܎��cd\�p�݊���E�����O��(�?@� 2ey:���cB��abԀ�cգc����`Ps�i�Y��b�D�����}s�C�n�ѝ�!*��4�V���$�#�u�s�%�>7Jg�.���R��U��o���VK�]�,כh����
��i
�d�f����掾�C��@�D����x���&8P���A
�U�kH�C#����O:EA�$�w�*;q�$�0�AT@���	A��V�k 4"P0���0XN��\�10k��mN��y�z�R#�a�l�/���E�$.v����)F�^R�*:��Jr�h�2V�jx\"3�gk�v2��n č��S��l`O�[Hd ce�_�/Yw`��^/���O2���%�H��h��&#�b�Φ��2ˮX 7ǈ�Z'xA�$�tDli�}8�#�<�'�ċ������S�&��[��:�"��|��u�(����9vo>G~��>C6��Y2ǿ���H����$ �2g��^�aB2�6_׶�d���)jg��b����؊"oIHD�]2����>�7L���dػ�]>�^ƛ.9�f��
z��Pf������G$2�N�R���s��#�4��s�H�53<�/^2�=`���&5��;i����3j�m���!��v�</
��G�� W�����B%�*���%n�g�xt4?چް�d���@&B�^�o�hЈP�^�6'9�H���u���t���f������\�y��c�˳b���=�`��X�N+6k��a��a��g���v�"���^��E�`�|��:�`��&Z�zt���h���ݎ,[��-�pp!��;a	J����{3���ʫ��T��/ѾְT��h�\����W`�7x��K�t#>���-�h��F�Vf@�A2�z���D`���u�Y��A\��\��I5�����|NW��Y��?J�_8Z���N��*9Q�d2M������MtŔ߆h�v�5x3w�Z��ΔU�-�p����wa��iiL���<O���s���ݟ4��|q��؛A,z��rG4��w���z(�^}�ZW1$���=�H�8F��OMQ�3�>��B�e���P��u��kX� �~�<�[�u�D�����f�U��x�qׇ�05ط��>"A���B,(8m<r���V��1]-!����͇���xo>?���d�X��Q!�Q������^j���Z[(iR�ޡ-H����b�C���5"�/m&��靄w��x#�DF�N��������+��PG����V�O���ْpk����5)3ʇ�K�ؿ�⯓:<S��t��u�֜J��-�����W����U�ӄ�#f�x^" ���e�j����d��M�؂�pm$i��e�4~��Ⱥ^E����"/U�
o�/�7��Vp�j��W��īY�>#�Mb����|`�{��ۍ��i_�v#b3D�J�$@�P�e��sR�mp�����;W
�q���tj�6�B>�dIT�c�҂x7=�9G�p|.��9�[C2K��u1����J��\8�S�wջ3rN�����<��&�Pjl�PR"ic�W57�0K�pxכ����P7�Z�p��Y�:	��$������Y��K�#$<�1��!I�����Q|f?4�uo��C/��:�N�\&�c�������n�dqE��w��3�X; �^����n���DRv]ғF39gw���	z@�(}#�4�+wj�	��I���O��U��0w��40��v�<���Z�[ԣ�\`wg��f��Ac�=w����������IaL���Z�P�j�]í  �b��+f��"����&@����=n�*L�j�<�w�P,���`���!�z�"-�l�HÖ�[���A��T�:/�f�[���o�(;���M�r�i74��j�#џ�L��@����n"����%� /_�Q�*�f(xeJ6�D�z�c;�N\�����������6��0C��ιw D��p�`�[�g�j
疈PG�@6��������q��,�>�H�{m���ت��G�M�^`�C��D�"��O��0P$t:p�t�`�ϭ�În�BTK}q��$aA����r�x'b�
8��֨ r$��Q���?�>E@|t��qT%X�ۙf��(��ԟV�9 �.�1�H%φ�1J��q7�d'*���t1��6�'&�!�;���䣘��Y��N��3X������+ۦh�tC>���tl��Ҙ��O��& u̪&�g<1���B�����} {6X6��-�'\`7��M,Z�O�Im�$�{�r]/N��6]���#������P��wowO N����N�;0���������QEQ�"g�u�uB��O���5�T��-��4�	���S|@'�;
C��G�Y�s����JBp��R0U{��� ����6��d�vv�N�%���A]l�#���<�џ��q����'�!�f�!�S��2�I�˶癈����-�h�l��)�v��@Y
$�L�L2W%�v�#u��	��m^�/�P�V�>G=G倧�ڋ�C���c:��.)��tv���g�����1{\�Q��c<��'>S6?n�Og?�s��Լ+��&yJ	��l�I�𺪝|;'�c�$�9�r�,�	S��c@ꈣ��=+�5�E��큌Y�3���|��
ל�gj�T���U{�-m`c*�\�\&�cQc�!�:,�]��L�U�ƻ�Q�tP��#>9{��!D"�[���IFBe�π7��3�9D&j!>yr&�K��(,�lR��� ���>Hl�b��'��\���]$=,�M�839�:�� fY��>���X��9���BP�\�:>��x.�Z��-��Jǋ�f<\s�<�+ů
���g�Q��cJ�~�'es��T\�פJ�����8u�Ua{=	3g<ƽ��e��N�(򘸃G�����\*�x�_C�'�#�y� �=��Ŀ�[h�y��B�	��#��.q[n~G7!�<�����ihp�W��%����$��W�ח�;8	��D��X�c�R	w6�L�k�5�˰M]�FC��,��7��Mַ�L{�Ш� e�d����v󬒺�(����3q+*��r�Zj�5f2��ȴ[�pC��S>y�`״V������%X+�1�yVf����ģ��������bH���"�,Ir�'y���N詂.�俖��8a��ӛ�D�ڂ(�n�3�T�J�p�-����>��#�nL��ׄ?M���(��U�g,WA}%{�2Y�3q����@:oT$w�� �.Hf�9�Mq�F�#���~���Τq�,ԣ>�$�N"7h���{LS�@G��QÀkF����g�8��	!��Mw*�`}����A����j�?�E�-��>���h�(��ȫZH�����dk=_-�W�%��fCk�?�CRu�W%�����΀F9EF�Aᵀ*��P4O�����ZwC�/ƍ�r�4��}A�r�<�o��r�����W�_;Pq����_�tz����yE�������k�6��h���yd���	_"�F�i��m�
�G�!"����ƨ�3���`�Z��O��������eP�zG���H��M�#�|I��
�]����hg�uǋ`إj��\�9�J�lz"���pwIy�=GJV��$W�����ǣc�č/�A�d�����D�v�x9��ޏ�H�V�6��2����.ඩl�C�)	�kA�������Y��������GI7J6}�FA���Bk�� �$OxE(�<���{�c��]��t�=�d3K�dGW#hǾ&Vˀ,O��ݲ�1��|�gL�S�J/� Qצ<�B64�Gͼ��R��u8�_����]��h�BݖǟI��c��$S#4�|P����:�P�)�]+
�P���J��g�OM/�}�Sߒ%G��j��>�(�/l���z�X!�&�N��qvuG1X�2m��������!�h�x�<�}Q\O�m_�Ɨ=X�E;7b��%��u����mJ��b�u�g��j�@~��rؠ�83���µ���s�g�[�UUX:�_ڦtΧb�0Qif�����Ϩ����s��$��O}�r}d`⇖sn�]#�LfH3|�i˩�A���QD5��rwY�/�:���2�ǐ.������g%j���G���	]��P�%��g�'��r:���(B�>T}ݜ����w�_�R��<�3�ҭ�72��J�����
K��}/�⦩^�_��
8�/�ϑ���~�ۭe��KE�T_�%~(a5[�
j���oxWKљ����c�W��~یF��`�φ���-	f�-L�%�����f�:��tl};r�4�F�ъF�,eP5a�XA!B֗��,�!��7�c���1�UT �Vn�ȩ�EOƕ��S*�`�_)�{����X�#���W��G��^Ǡ�	��
��ο�y���huR��������^v�3�,����mBa�G9��KP'�CY�0B��K�2���v �����&��ݗ���1��]�D�9φ�Lj��:��LF�mu����������ŧ[~A�9�j �%��ؽ����Y����	���]�3�q����%ncjH\��(��/�_?15	I�7yR����n]:�)h�y2�߂m�tO��#��'X�~AQ��i��f�����W���+���P��\�L�n\M��Sb��"�8�΍�����pz�&����Dnw�7�Xd���hʳ������:��7ż��o6�sN�="a�i�W�5���~��>}�	,�ŋ��<P߂88����;N�5"�d�2���\�^�p�]�cY��w>�Z�	��������泅y���/���%9�	���sI��`,�4bbs��d=ľT�c�ߛn4QZ��f�ȑL�����i�ot�̹�m+�kz��B���?4Z��e��4������@���}`~W���(:��I#���4�o�#]ܗ���MvK��A|R 蹄�e�n�R�?�.(��w8N��I9�L�����/��x��%�?>�4B��<Va1�&";V�n����3<3���D|�Ñ�4^7���&�5�a���c���+�C�N s�l��ў��������ߦJ��*y�&��b��oZO��3%����DU@0?�qL�����u��)s�M�"'WJ�rL>D�f�g�c��;&�X�o�i����4�C[N�s'���{Q�����G{!b�PC� �(Z����DF��1<�X��#�|U�1�V�Jdw2����0�ͬ[�M�����T~�ŪDԁ�1��M$r�����a;��8\��Gl��&�>��a�+�y�K�Z���i�J���O��p��=�{p"�\dUT�=�&��tYX�!���z�X�Z���%��n���$R�T�ѫ��y(���r��ˆ#�렾*խT���]�w�kt��)ަ��^h��d�3�|9R2S�Z1;������1G��p����E�2%,�q�.0�ڐβ�uw`�,���1�oj漲�.�\)���C���3���ƾ���Awy_6�^D�-!���	�!Ie�H~��> �B�K�2�!"��}�T�ٿ�&r�R$w/�/���낹�U~�$�����Qc�`��ƑSR��2���uQΚߴ�.{�ŗm�<4��=�}7���,Л'�-$��4''�������r��Ǘ����!�>>�/����)s���]�'��\#,����lw/U�S�-��',�է�&�tH+͜L��Ȁ��u<N���Қ�.�X�|jb�@KS��S�[�BA�oW8T`�P�f��u�ߌ� �����1�8^���ɠ��<c���d�B[$�H�g��s���y=�~1K�&""�H���@�r��VS�~�+��6۷o�:#�]��ɌD8���FV���<:��<!~�ăJ$H���i�%��I�D�Z{!NE�[F#��IF�σ�7�A��dt�Cb�b���f<O<�<�VH��ٻ}�����4�k)��E��E:E�7:k/���_�Es:�n��}b��8c|���~�ؤr3��{�Kc�ƘM��S�ZQ}�O���֞.�繋��H"������ ی�ȇ�{ep��,���1��F�ˈ9��ˇԊS�cw������J͎�$���)L�)h�I��-Y��F������������gi��R�-�P���v/��DgEӓy�mPGZ��?\�P��������}�ȂS��St	8t�Fn�j0#%�k��V"�=��Å��X>���*��:�|:�n~#�TV����I��I�C�7A�{��̊��-[�$z�c�c������y��a�<��XI�4�h�)X&�%�ï�'��c���
����J�cE�4��eN�LC�	��ڃx-���C��Gw��L�-�s9�<�H����r8ʻV1�
�ٮ� �?Щ���R��d� �TwDwҬ���(N�*!T:|�������Eg���޳JkË��ͽ�+k5B=�HFd������ա��0�N�T�����#��)����)o���Ƃu	W|8d=Mc"���DUÊ�e$&U�]qQ��%O��+?+v��H�������`w���=C��p*��}��NV���
DG(M�* <.b"#}��>C[������E^'�^1�Q�$X��ۀ
��'iv�%~<z�o�!Z�����;�U��[By�#��*�PF;��'a���6cS5h/As6���'�o��mus3.���%>g��#��Uמ�/��t�5��g����F�i����G��������g�
ufpݪ��w�/��D����8Y��-UT�\���؄kȰCn���
�e	����c^9h���J7��6q��([��P�-�I"��ڀ>�����{� �(��c"����V��pؽ��4�����t��.I\�F��%�fJ�
�׬�]~��.������U� %�o���M�C��,��z��'��j�Rk�~�a�	����e�T	����1�nZ�R(#�Ř��WZbEm��(H��n�t�<y��=��e�.����ƞ��1�X�=��sV�_�>�i�ؔ���2r�;�1_}&�gc��!�tM@��U*�=.X�&t:��� u���o��J5\�	H�5(��_��=�����
��QY:�oh=�{��˒g&J���ĭ����^��ۡdT�=�ѵ�>�'�������\���%��^J=U�e0�HQ�N�ퟦ�F9H g�D��P��R
穴����眼��t�w�c��.VmCΰ�kK�����e��Z��\$���(�.�6�����1��GN���4+��BԲ�#�Y������y2Z��Ӡ��������[\��7�R�tv��Zß3�y��T�ӡ����a���\r&lw�z�}|�7 �aZ����F��S���X�To7�t�"�7�=} �d`���n��c'0��J<Q�2��'v�T4ׂ�c*�#�=���� ��<���T���s����M9�ayA�l����6\w��������Xe�

mv�^����&�<����ضm�q���9�n��ҬI��	qJ	^���@%�:HHׅ�a��FI�uS&�p��|�Uͯ ���"t�țM�-����^Ll�$�fZ���nP������bڢO�vY���V�:���}�d����hqm�T[ϻ�����d�/��j�����_�Z'��P2z�w\](�~��V��-��'_R ���;�G�����KøA]SWG�:B��5�9Jˡl��Ҋ͓���b�'B�ښ��I7󘼡�z��~E�,I���~����C�n��t�Вo��B��۔����<�aQ�1H�y�%��Hd�Y��."nb�ɑ4o�P5�������)E���g�6��b��(�p���c��i�f�v�rE�lB�%P�U�X)��3�@V0��3��a�
S��~p�uUGP�Fb]���Bjk^J��ׯ$�NJkD��'�Ȕ�p��W�Lt��[@똎oPÂ��p�r����P�c�kϯ�-���GĞ���Ҫ.���yk�>XיP���4��jx��(!S2����p��YlaB�����؇x^�_ƭ���6m2��a�󯹺h*��r;m�6pE@�l���7	nc���&�C���ĕw�0�g-����hˑ�J��ԛ �p\��'_H��;}�5�q�F� �1��IֺU^���;�K�tS��W2�� ���(�C�t�i�5��GP��,�-�z�u��N6<��6W��%~�x1�
�����}x�И�x�
��x�r�M�=.� �t��h����CD5auj
�`Y������e+?R)�}R�f���Wߌ �������05j�g&�<�L�8�W���6ш�� �r���8}ә���k@-/�b��~�B�9�_���3)��緋��w��a�Y�#�.Dٞ��g�-�v��y/Gˠ����:����k��Ni1����_;��Mc��s3����oE-v�8ҊGI�,"�95D�H� C�����4�O����g�x*ԡ	"t|h���� :K5�_�L�3�����yB�'$#�#&8��)*%{%I�7.��u��K��={�NsF9����11�L�˚��O	8�cmu)�.����ʩ7i�n��$���M	��*|=>�Ȕ��g碌��9"(X �������[�tT*]٥�U���̵�6��b�1m�_!�LS�1�.�ՉB��%��Ag/T��ݯ����h[>oܩÏ[P�����;�a��m��K�>f��W������O�u��{��N�.�����:F�wM��||&���'��]�Ex\a��x%6U��ݠ8�\:�q�/#r]�h%�[��)���ܴ3!ݫ��s���d -$��<ao�P���xùd��n2�8�O��Q�]a�����OL5kl�����nz�9��Svn�Z����i��œ��p��#�E��@={?/�:\�7Hsf�"�+��������δ^��_�৥�bfQ�����ܫ�j.�#��M��v��	������.���t�� �;}�=���?7'0����0|�xλ������'�zX��Y��=�ѯRgQQ�'�b4m��j0�7���%M��������8�p%�Y�k�*2VLrǀ�d�RN�6���!h����@��XV�H�#$9�y�q�-���� ͇�G�"�1=;n�Y.ǰ�oF���,˽�+H�u����>�3i����t)������"�6�Z· `�Ҽ$��g��T�s�>�\��0�n���ƥ�?�8�z�k5U��1�4�p�q5��V�,�Ц�	�{J���V��(� MxB����l��*G��.�G��3ܲ��nt��o�Mly��*^} �ʙ��,AT8zē�E<���"���a�vg7���M��cI�Rh'._.�6@��,!'�Cdiëa)J���@�Ӌ�����˅��(<�k��RH�w�\v��[�����=�;Ü�y�b�a|����J��]��u��&�?�y/=E�?�R}@�Y;�}���]`�#�x��"��6�G����pЮѳc�2��p���W8d��$�U<,��ۭ4,a��ߣ�?��ݘ�J[�x�G�+O���k�|�qO!SVސm9$���=v�����o�q!�у�~��\��r�R��]7�c�%�;��7�8�8���(�7{A�v�g\Z����!�l��j�dP�m'C݁&���>��S������OU��{߫�[@�C�-er?�n|^>�W�Y����'gO� �=ոo��C��i��)�ɔ-x�k'A��[��^4�D�������z����ʓ}����#�䞊�eH��'M�c����6=�d��c�$�k4v���l� ��е��,�<wB���AT+,��r��z�
Lad{��Ayx,��i�Y0ۜ� %]B>�Z�f��Ju#oQD�r(zG�;�ތ���.��E��rل��A-�R�o��A�W�i0�f�*�(�W| et��Yb�HCc�I�	��� �4O�~+��G�)s֣�}<�Bw�x�?����" ���^UQQ���)�#K-��=cd4��9���cę�if��m��71�wPf髭�X��ռ D��z3ӛI<���	3�%��]��	�i��/���h
̞?���e�l����h�As�k��\��Ej�<�!DM��l(Dׅ�0�ҥ-�ݟ�F?�7��HO�����/������}8e�9Q����>�Vq�C1)��Vg�td>��R(V�;�ϊ;a�W�ٴ'�T;��ڏu��aE������ݶ��E־��,�;P�B?{��)���G�Z�wy��?Hv������S���T�s�ln�K�"�J2�鹌�|Έ�uCV /�#Qe��r7�_��:h�L�+wڹi}vI���Q(���jRcac^��l^���av/8k~�G1�^}_`1_ZR1�5�����E_��ZWmg�{P�
���l �FJǘv|&˄��\��;��P�MsT����mc�9H~-�b&:�S���nh�(E�8���l�D������%R���_ѝ���#c�b�𶼒�4[Vp�^4�>/lE����gv�׈'�,�v	g�µ;ț�nDE(@d���ݬ�Hxh.�E���S��{"���`��#K�Yaa��*�6�z6�hFs��C�tSbM��s!qӂ�<AmY�@2&F�0s4����Q{̢�ʣ��u]�'���8�ۻ�j�gC�"�{����
�8cf1�o�[�C�_�I�z�	���	��'�6�Q�~�/��zP�Y�������g�`7k�h�]@��ui
��!Ϟ��7Yv�T�M�!Zc�v��8�T��A���2ޟ⌍�q��R���ɫ�u?� ��~�C��~ �uZ�z�M%7n�(��4�D�=��d _�L��^��S�H��\��wH���£��$��Ǟ5z�v�7	,SX?�>��e� �\�\���'P��Z����]�P\�s�����_��l���|h�Ƴ�MWWh
VR��3�Ԑz@���f�K��(���-��1��Lj��i��}F�#�g;����`o���Չ����
�#�)�����g��b�'0:�C��7p¼(k�P쮰D3������퓚sԊ$=���8��1�c9/��p�۟�:2�-yT@|�� �,��W���d�2Y m Ҷ�na @Ϳ���6q�}�j�1���d� �>����ݧ�3��m"\�G�G���u0��S��|=��ӔmB�(�7��lʜ�R��C7� <�.�k4���j���6��ο�dO�797g�
��;�7��Z<'��L%w<8�k�U
A��bI�_c�8���M��\�ް�Jج,9e����r	��MyT݁��`6gςAMŧ����&����ׁ�R�'���u�v���H�W��/ů^钃�t$��"�  ����F����>-*��P)]����~�����"�vPHfƞm4:��Z�_#s`O�m[�X�|� 1v��/�!cQ����`�k k.��6�Z�!=80w�P�%���tc�C���2?�����ק�o�n�=õ���ژ�l(�R,I�G�[=�4:cm4����q� �
\D��	���ɥ7��tv��)hB�4�]�
��ZBS�ٺi��a��Ht�)�������4����EZ#��H&����'|Qq���]���4�>s��R�܌��g�%#�w��6�� �Gt�T	X�bx�&�0�:% �j��a�,�Td�%ࠂ�p#r����C�����ܹ%�.�]��(�����M�_������W�1T��|�����"}Z�<�"����/�ff%�ΖII^�ZzʦB�.X��lE��5f]��,Ŋ�Wncü�n���5��W�u�J����Y��t�O�l{kp�n�|�s�\B:�R�j�����³�v|{�C����Ez�xI�"�zܶ�{����f���m��t�!.��J��?�4c ���lm�Q8UU�w,�hL����Wܲr3��zq$09��"���w���T���!d��X�� N�^������_(0m�\� [e����Kx�;�����B����"��5H��C9a��H�%��l���	"8�W�eم}�]�g^�4)O�~�'���2!�<� -!iG�?D,f@�	_\�A�IXe��z5��|�2�������J��l���S�]�.�kK�4���)ħVM�W��A�D��WӋ�n&t���r#��!��h��@��!��k�흟	>kU�@]�{�Q4{��g��f�+ɣ��5��;.�}������a��&'�EQ�%���X�x�1��*�p����O�m�]���68���\@�Ƣk!�̵J5ċ	���9�1t�ı�:L����L�׮��B��Xtsɥ�O�FKyF��?�J\�N([�j�8�%�����7X�'��vᢁFa�`�=���|ޥ�������N,�r���j�7�귞U�W� B�32A͚�;�����zV���$n�.w�[/�P����ߧ7b�>w:Ԍ��?|e+����l�T,m�Z��_���[+>ڦ5��]%s_�i�zX%[}��	��u3A|����D{��Y�w�� [
�l��!�aJ�-��|����,����0�������_�v+H�W����{�]�O�K��mj���U�7/�n���[0�Q&����ߺF�E~]ט%4SM'�X�u�S�&�s$��k�D��*7��᳕&{[�;�%�ۦ�A��Z%=�U��E�p��Å����_���uzV�\¾ZY��y�I1qs_O0d�46����$�Ln�2U���aWQ�p��;-��h����\�e�, Om�;�ρ���9Pi�����4=(��`s˙X�E�Ɯƪ��qܗ�V�]���Nh�t������R�ZT��]�q�� ��D�nV�C��l�{Gl
�G=�������������x�^���](�P�v�grK:K����˨��������0{�Δ�UB~�o�
G1��]�<�,f���2:�t���B4�Z�t��l_�<	3�(�Ǖ2��SM����l�?�����_�;JK�C	�Zn>TP�iQG�z/�g>aTO6J�`{�/�`�G���gz��jEI�%�
�I��U�-�7�Qf��J��a�K��0=�� ��$�q�ⳳϞ�yS�/�-�o�gw���s�2��pP�F�����~4���/�fR��U�=ݓ£��=�p�Yӈ��e�\��#k&�pWK̃��vIU�';����yi�w�if|	�M���c48Sᢻ�g�gPޗ�f���h��Hc�Թ��rnx2O�b�ƚ�j�6�MT�������~�t6m��Dǽp6v.��D\���y���0z^�X/���?�3LN�B<�Ө�/���U�2��\Y��WW?H�}�.Md"��-�рD�����|Cd3U�~I]z�ǉN�s?��HG�X u��¿r�Yö{d��$ز��ڽ�^�hrW5���F���c�oH�$#��aqϕ%� #[HfrQa�M=Fv�����6�q�<I�����G��ӵ0S�ɝ�l�Efr�A��䖂��rx)��5��m��Kdi�>!�[�k~��'������4	�ųX���|��XTo>5��T�:�l��V�S��ZP�(���%_VN~���R����S�e�<Q�z��g���>s+�#�ֵ�	8lG�UA�J=��� l=�dPV�<�y�P����ջ��u�[��);��GN8*T�J���m��k�L��>���"�ٙ/�5�OH���z�d�b�7��;\��1^���;~Ji��R���V:��F���-JҨW4�H��X�����_>8~Q�ŭq8���I�uX;w��/���8���vF��,���C���M���fo���'!�-jZ������;W�

s�|-�y��[l�����h�n5������=�_1�+���/zvН���^WE�o��8Mm��k=+��ǒ�@7n�wȮb�Ʊ�O��E��a"�W��X�/��~�N�&�j}�e�.Tu�~IX|y�e�S���4̏���:���TCp��#��#�Z��x+�u��$�'	N����~ZdN�%� ����־a&L���i>.q���?݃&U��.���uI��G[���d����U���(�O�㷦�ܾQf!)��c)N���S�+຾ r��\���D�
a��8/�-�[fv{��V������ι�_a����D�H�fj��؈��z����	�j���&���<�m����+�nr;K=ZԖ3f g����")�	l��,��:����$"��z������Nc��2[n0��]�T1ͱ2(�aA3X5K )s$�;��P�Ev#Q E�g��Q�?%יT��*��e�ws�s���V��k����`���\Hy��h
LP��{Ǒ@�a2�R=�xIqU���fvgXL0%+Q�I+�����K��@D=�!1m���#D��.�pz ,$�9��ⷂ��`����Q�/��_���6�0^��6��s>j�b�����R�� ��,��Q%�u�s��=A�B@���j>�!�-��#w�I�s�����Ψym��ݮ��Ͻ�ne�4"�"CQ�w��:��@�!���7p\�[K�LaI�i{��` F��e�����=�3aF��b^����Y�����_��H\�	�y7��� X��S�a�!5��/�\,+ ;�ж��?_�43l�:J��"p�'�.N�*F��u�Ͼ�{�E"]��~���>�L7<e���E�(U�㣷Q�YN4��	YN�?�2O�jàp'� �� dI��� �AK��,���Z�v��8�eԥ~��3 �\Y�jv���&��C���D>HLT���e6��i�����ΡDg��N��y��w�%e�=^C�-q�Y�jC�I�s��5�N��6݅�`�D��k�ݣDZo�Mh9�>��R�%xrJ�ĲU�;��G�2	S�#1��d݉�����2�U6��Y�3��@z{������|$�o��q����91a�z�$6�������V��~D���`?^Q�kWh�}�[Gؿ-u,���V�S��}C�]2&���8k�e�����gA�bZ@�<Y���qkZ���$��$җ�� P5�ܕ��c�[�-l�@s�$qn��$� =���z��Odx?�m�SO��*�0�����$I
��|n���O�ں5t��9�P	v��3w�(_[���#-a�t�I*� �����c0Ei�(}Lg<b3�E��H?'���;ֳ�ⓀK+<E"$�-�ᠧ�|�4�8/-��&���֦�W�i�y�h�M�I-��a�ΖAg��) {�zX䊂S"6aI����<V(����}i�dQ�"��)�N6@+�y)⴨*�E�J���c�C�d"�d!��u0�<6�Qf���.��h [�`�mg�Pm9����.>����m�x|7�JuVuj�D8N`6LJ�v~jO,�m����o� F�io��4�T�9ql�H��X3SL�5�+ޯ��+�'�6�P/Yw���{�~��qLW�D:P���1��S��QG��+�9�Bd��YIO���5�Nt���!e�����#�0�Qjb�;���v�d)`:m#�׎ڜ�M�kC�+������o%�:�0�n/���9n�[� X�����L��P@5��npm͗ԉ�ۤ��ɟ��t��
¦F?/;٢\�x���a�
�#�y�͵��m��@(��
h_&j�p\����P��^D�v_v�ϻ�.��t6��h�_Jչ���D%�I�»iFueH��c8�k�[�0��3C7%��EL�?�{Z�|w�.�0�����:,v��+��˕R�z��Vz��{8���#M�/QY%�:���^�,ׄf��/�1���q]��q샚�����{�z�����з���֫;� ��t�bGM�g��gm������I.�$4�g����rQЄ�Q���Ln��]_{z�t;���`�
q!��iL�;�aacU}RD�\�l�*r����*�X��	A����O�ģ���W��G�7�>Y+�yMZhjd��j��������M��u��鳣'8N�y�U�Υ��/5��;+d� ��ڶm<��~��>aDA��8P���L��wܼ���ξB�Os�Ǝ��Ԩ	��G��8*��=�eq� {�N��k43�����k�h(+��wdACӾ��th,��J%1�dE�t��lc�e��J�������oc�C$��7�V��a�۹�3��D�9.p<���X���ߖ���}V��]���ݒW���8��H��pYX/�Ǽ�����5PE�����,��w	N'����|��x����|4�Ӏ��7Mj��c�q�y?ߡZI�tQ���d��R�Αiy���F�I�<{�+'���x� ��7@�$��:�"@B{}|�Z��҅
%4*t�%����X�祍n>!�
I�D.v*u |AM	���e�Z�f�P��T!F�eD����`�Q��Y�s�78��4�ͽWr�ֆ��W��������\���۠0v��|Xjy7C�s���ܪ�h�[�}��Z$�����"ӛʀLs�+��I�7��Z%�5��-Q:5� Z�\�c��S��Y�HSv�^�x�P����SzL��8@��<��Ic�pY��S�b�	*��,���F����r�`��w݌Ͱ��cC#M��I�b��6�ܽ���$��i���Xf'jMv�qJ�7��x
���P,T=�l]���?�R'-R�H�}ρ�>L)��fE�`�
�r�>]h�@+tTb(_��}��G�9�53��~�{3����[�Qi?��+Or�;��)Y��7�MU]Ao�r��_����:v�79��V^�n�aW�j��ݰ��ۺ�O����2G�����z�*F��k!>���8L-�%��n+9���ٜጬ*ҷ�D��@��~��?|�����hd�@�M�Y�[ \ �����al�'�V '⺘�s��8���&qm�g��|O����CJ9 ��|�|��I��c*��[��Q��3
�z$%��J(��jXUk+J��?��X̖��g��;����$���F]<'�Δ�;W4I1��)�
y�Ѧ�E��xSt��Q֞S�^��8�T�b��w�%����2Dz��HNx!��%��3*���7�{y[T4�������٩��n�6��M=C�r��4X9e/�C��u��F����۵;��(���H��Q��1����@Û�l1������yv�_�ϝ�A:�Z�W ?����PC9h4ZѱR�������C�;�=8�Q�Td�/{P��њY���Fz[�r�Yyd��Z�����/�r�Iٖ�ʰr��4��q�o�������Yg�	C����
�}�F�kD~��3�Ci�H�@�r�N-��>��gR���ۉ?��^&��=���	�X�K-u>���F��1#<�ϟa�Ł��J	Μ�`��mK��
p����B���D��X��7U9���E��?P"�^�]�����K?�dd*A���BP�k����*KA9G�t��S����=*�cH�LJ�WV�o�X�"cg,��o���Z��m6�/�~/1���gR�P�V�U
�}́R���܀��K���x��8��!�'�",s즙��9z�/��x1\��[B�CGUPE�L�����5FqCE���
) �H��-��j�~��3�|� S0mͼR�g�D ^ͭ��h�O"}��jgvhah�T|"��Hg*�6K�^��Xp��؉T2�6��{ G�,%bL��v����3���;?���nMM�B���}=#�VH�vV��˝Ԝ�]�ǿ�b� ��٤݌�q-�(���2�U��ꔒ8�w0�XF٧������Z���~�=J9ks��gx�x�NH˟�}C���S��һvFk���T����S���j�~�|�c�o3k(0���K�t�QuB�lǎ�������i3D��J�a ��BO�(#�d0�bO:H��_�\�!���ic����	�KШF��"�=H0DE7�S��Ó.Z��������)WM�:G�ԅ,ڳ����������7�i���] ��@�H��,�^W��ή��X*�C7����Г��t��V�,�vŘ�C[��vO���_\˧��j`7xn�	�k�nz���ŰdWR2�$�u�!��O�-���G����k}Ş��)��.q��ȸc��HH�/&w�92�5�N�%�6��.��@r��ji]U�vV׮!��qrAdax&����nq�[j��܏Rt��vf�����C��o)��V�z��eG��=�uj�����>��b�fTѰ�IRk%�4���ˏj���A:c�h]�)f��],<Q-&��V,ȆY+ǚ��,�}0z�Ϗ�[�,t�v�ʡ�F(���%k,eY��Ŷew/��/�PQ�f��L��d������W�W[��~W�U�����CTq�X0�R�t����K��q}e�i�팂j���#�l��9��@6�>3�h�3���Ӛ�9�1cќu��v^3OQ�*��C��I\a�ҏ�s�~x�	7�r6̹,��6���s��Dc�ӈq���A���d�:�9�e��HI�Y7jd1U$If3�r�I��� ��0���ޔR[�u= �S���>.�d#�G!�x�G�~�L� �_�G�D��^UҜ�����|��S�Ѩ���1U])�%�OY�T�1�eB!%�CDj��Wg<;����V��~���/]���R�%i�Èo�&���n1H |-L}Y�r����z�`��+�{��p ���Ⳃ��re�x� ب��TeR����J������w�l�T�F���m�ӟv;	>��Zo���g�)�}KR1|`��<�D��aQ�?X�k70���xu����5�H�?v�4�m�I\5���uA�όY����O�w���Q<^AܪvQ ��Dt�w�u�sl�yy�E�7�Bxl��+�ш.K�-�/�|����a�S1@S����R��!�d�
����w���9���b{���Y�Li�]�,!���5�iC1��V����)�L����Ū �����^a?����-�o�w+��#�]� ��x�؝�oZ�Fdq�7�(��-X�)�D�h��Z(���ϕm@��QCԫ	��-Z`���.K�H�q��<�3m�Z��������H ('!.������|�)cH���e���`�>�5��;D�)>H��n��$#���������Q%�.Sh ���K0_76	�v6�]�fD�n�7�X2��Fz��b���a�#	�E����{)����mt>P��YE`4��_0v�H��5�^�ñ��a�v�{Qߣ�Sj��T�u�eX'��T�Q�Ko����C�ūZ/3o8�r���Us��L0�H��=W�1��:�+J��2O�UY�/�o�><���2��3����B2�f��v^�b�Aiʜ�#=V�p�b�z��F$���t�ҟ}�-���;>"72�J���&B�$N��������Y?���ii>��� ��<$~�T�8��e�ˠk7���W9�zF�X%ML����5D�ѯ�sKu���>ռAH�"�K\�#CE!Wj��>��bɌV!b �h��K�b+��h�4ؙ~.б��עn�pφ��i�nQD�(Z��i�"���5��l�B#�]}}&�^�� ��jj���Fg�?��N�h��}�.35Y��Z2%�%��
�Wo7�s*��Ծ��=9CmC�=�p��V^�H R�?�"��d����ݐ�Es`�A�b���IU�<g�UO����ն+Qަ�����P*E \.�ۡ �s�$+ p���~F^�S5�ogq�L����0mk�!��^�dY�<Ҕ�VH��'�x#�z$*񘯬1�T�/�1r�0!��Y� ZB�Of�Pm�����8ŵJ�6F5��� �˽�v{����"�`�ߌ�����i ��Y�O� wnE�f?xش:�0�+\�^�r�V��j�cz�%}"H���CA����E��b����V�P~�O�'�{���;���L� Y������df�ߨs1�%8�?��mԅ�CX1F
%�L�m?�j�����m�J$ź�KA��'Op�!����-Ma�'��v$��m�t�m�\�c�t�<+I���$�AY����Æ\[�z T\��%�s�n
N\�=�V��X0��F��n��fG�����T5&��V��"���F�*�ƥpp��ъ�U��� ����� ߙ�X�O�uqZԏ�k�����x�rx��F�1a��)�x2@ol�8�' O^(�[/S�bT��9����k	��T8�O���Ԓ�c�L�N&xZ�G��P�˘��K����I#�X���E�N$�St�>�^�?>����d�eу��J�ܒ�KWg�C��^�tʹ4F��^����Ɋc�H��^��Q;���7����1S��<�bOd��ψaq��3�s�ʅ4Am;e^�7����αt������>�퀱$�⌘9.+�%Ԏ&�[�5�I[B�@���{T�X_��Y�ڿ�(F���j�DEel��^&�ji�.�>���Cѡ������&]&E2�o��82��׼g�ゝ&���:��ڝ�Oc��}���'C��\Y��%{#|�����{i���{��.8.�0zp9y�Q�x���Hȑ�=t��U[��A��,(���Mv��Y��9~^; &�Kw!��DQlR�@*�i�}/L/󯠧T��ŪZ�jHۍu6�ybI�SM��r�-_���%دOY�R~C�R	�W�m�j؂�Q��8s��$4�� {S�r�`�����H˨)�7��m�X�v"�
#}_
΀<�,�1)�p�m������y�5�E�,c��?�ԍs�ulx�E�-���[kw�5S ���n<�}��Zc׆Fm�b�5�S��X<.x�蛬�ߠ�o��8m_�~��$0��D���`V,EV�/N��(�)gaZ�f��FC��f��[6��A
>��c���J,W=A+�\�㯇�"qrv
���Z`�D51��;f�M��^�ޕ��+K���#�$m,z�7�ž�׹�7آVj4|��,2#B)N���W���ev�٦j���u�Z�n\��5��M�e/Db���Bݼ ���05_�H����)�{��+�j+Jq1�V�}�c,�ݴ�tF}#:���V��i�;��g�`���ae��E$�Pv�[�QQ@�"�Ar2L���+�����TL��2�¨%�}C������̱w0�W�-U�Y�sSv�_?��L�?s*���iu��6o����Ļ0��������6h��L�����~d)���9!7�izmA���s��b+��z2��K{���е@�M<�)��S� w%�s,���$�/bX���|�)={fx�S��v��fđ���/}���2�YM����d/�?�g$]!��^�G,d^�J'���
���0[���˕�P,V��s�j)T[vI��Y�ޔ��Qoib���ǻYd�Y��3���^2���B4�b�k�n3���#�"�X<�^A�x��p�#c�n��/�-�g���e�C�A����է^
@��1�� ��?�M���c'�&�Lx#:�%6��p�=��u�-_Œw��1�7_s~3�mg������oLKK��w�y�P�/�Vܹ��i��?��o�u�$T3t�7�L���P9�䙩�at���
���xC;zmQ̐*��9�ȵ�{M��?+�d�l��Dt��[C��q��Z�8�BĨ�dq����q��Y�m������Oa0!ڼ8 ������MP���bBaj�,㈼j�Ԃ]��Nm�B�"����gbX�
V�hG�(3],�� ��	1_:�'�Ekq��"s�e�?h֭ �:G_���x�`,�S'��!	J�� ��Ԇ������@��7
���68��V��	ߥM�ѿ0�0�u��4�j�z�~�"��Ù�F&�f^�u���/FU���е!ubo-ݧc�*���� 0!�xL������	˨�b*��e2�}t���5�̉����b��7���~��k0wL
��LV�X�+�����w-��䓛�OB9FU��hi�$j�'����7�����s��]�sQ>�8�q&Ș�ّ���g���`v�v+�ɑ�q#�}mP{�=�c�"O�>M�mhgs�:!�`L�N{D&oT���*�Ok��l������S?���� }�;ڂKD�UѼ�e[����^ p:{S���ڵ��h���O;�`�C.�T��ɍе?c��n���D�ve/
�J����(P���	A2���W�.�����Q��B�'���1Y�zZCBB��"�N,����fn����*�!Ayi��d�lE�(���@�Q��$rAȌ��1�{��o�F�r&� C�vfM�YBr��*�j��PZf��)l͍ �oU�1�d'"A���E��W'�)y�)yucXSM�5ٺ݋��Z,�����i����z�4�x[�)�=��m1���R	�u�u�`{C�$>{���l6�����
�,謤��g� g�Bz���-��,c}�3����-��1��b��*l��f�,�����]u���d�Z�T�a��)%���D7�tAO{�lx
{�:g��r4㝛ޑ�gd���o]l�&|nG2I�[@@��0{T*�]mT;�/����-�m9�Ȅp����|�t�#*��x[��-Z�<�����Rf�W�%�O���h����i�������J�زg�<�^��)x˨t��/筁��H��l����k�����Kf��?y"�.�#� Ѻ�+ù&�����Q>���D#^֫��A�E�]�n��n?o�vM����f̼�;y��T���('�I6 ��4LD����FA/�X�YF����~���^]��4�.H���ߞ�*�#��3ѵ9?`K�8Ւ�F�?�9���0v�4�I�8�@�\$��!��^ἧ���W�jtԯ*M7������%�7������#�[{jWy*R����*�*M�tׅ�v��?�u��N�JW�߲��2���O�[�/��,��?#)1�f�
#�j���ث���ʭR����q��t��)�)������˷%� ��%G���Fi�-��_�a��Ѡ�fK_�%@��i���I���ĝaf?�Eh7��G��{fA���9i������b�B�ʅY���4̓�o��$�S�l�fRrL�4k��Ȣ���6%:�P�!��x)A�?��>RJ��rx4P�g�e[#���qB��g�Y����?������~I�zH����и���]	�qc�>�v��/)�Lg����^�1Tx�����i���&�����.�g�s@ٱ�q20�0��1w����]����޳�7�>� }�Rfں����`�����N@'��������p� ݅5�eW�<��n�^ #N�gS8'�~�E2C:�GG�Ӌ?�L���!S�_�MʒZ*.$��)�I`�t�X�-� R��bҝMY�>hDOGs	�X���@�+� �����hH�H����1��!�����de�bR�O��}<�ו;�">hA| �����x���	ye�HɉӞ���o�t���L��=�X��p�i�����1q�\X!֘zY{Ě|{�~H�ޝ���6�v�� �xFƻ��4���N[NS��`���
 :�Gź�0/�s�;8������
)`8<=&)X�kۆ3���]Y��K���l[,�\#�f\/���c��u�����m�]�9&��H��m< �l���;B8&���#xBcX:;u؁k�&��U�{��/+nX�<f*=����_J��.��e~�X>~G:c�dM�+F��"#�2�՘=�1��}\��ɯ�t��ny+I��h0)���n�YO��͌w�o������>�'�g-�n0Z��3D�8��������4b��n���5�V�Mi}��Z�H��E�B�(�Χz�����tD~�p���u��]]-����ӄr���v��*7��_"GՉi�ZW���O�|�dҒw����T82��ϩi��:�^��{�ۣE�'_b��`�&�9���0"�RR�D��%1�؀�7SCc���<�R�*��@#i�i�����fϹ����#�Q�:#��n�� ,V�����i��y���)B��w�gk��^i�+��~ZBĻ�W����f�Ctd������ba���yR��U��.����b�������̫�R�"�5��E)9�5�J�	����[`�ݗ�YRV�A B!�o�7@%>��Y�?�7Ҁ��@�(]q��Jw��W�-5�2$U d��{��D (<ʎ��{4��f�	J��|���Ѝ2䩎�,����<Q�z��3ύ�_(�)�h1��5I*�y�_q�Xm��(t��8�?�[�:�҆�!dJ�;p���{����~ٹ㩞>���B5F"�� N..E��*�gg�������V`�K(H����IAr�3��m��*IIaF�^~%ad��K�6{2�sW�=���ӘJ_1,�zF�&��pK�-�?4��F�h�3�&�$$H*�<CHŘ�N�
ҍS�M?p�P\e�
V�or��Ќ�n:4T(����׹l@�*��ә9.8�T�9h�}[���f^҉$\4�/]7���8TʰTTP��,��C8���[�z���\�f^���Rذ�{[�w���͠A��Eu��(١|�MRFTWLO�
�A-��d�4����􊻝 qֵm��u�Y�9�&`�C���T휊MT��uZ���Ȩ|�)�
��Z���z�ealDM�ma��Y�Ў��q�4���m�r?������ćE�H�ˡۚp�?m�!.�30������[�RVf�vm������w�5�(�`�%=Q�N������W̷��:�nʀ>j錝�c�X�����+m
����������\.�ß/Ӯd+�T�C��(Юj��U�P�a�%{�+�,�����s
�R禀����ˠ7��i�_�J�IŴa jɽ�R^"�Z���GP�Y%���	�h�S��� �v��-�Q��R1�-S�lС�Y>������Ӧ�"@�^���TR��øA��z��"�1Z���_��i����S݊P�WU6������41=��J�%���g�$�l���ݍUF���A�B�)5 BZ���5&ؐ�X�e�+z�Ңk��+��x�R~���\�`M	�3<��"5�q�J}���7��m�([�ԗxn]����O?	�����,y��r;Q��0sO
5����#2����q<��U�[(��@���#F��2E`�i�"x���w
54w��}@:�h��ZAbWq�̉(<H�V4i:w\Q�a���u{a�Yk���n�Tme���b�X̭̉�`�e下}�K5(6Z;� Y��5/�(:]�k�)pJ�$�$��B#�em�'�>�)�s	+T$�Љ8Ԫ�h'�LZ����7Ş��U�(6��mH�&X�"&b��$���#^t�=�%��;k���m�F��^������Y(.!������E̲/�w�	D�p!W�O%z���=r��UI�mz�$5�&A��U���F�8�QV�h�$S�OPM�t��9�w�1C����>��u=��y;�5��y'�{ڽqE�T%�p�'jS}<]��" ���S�ԙ�A��������4�Jo��N��k|U|U�������`��g&y+�C����
�x<n�q�ŏ�~����[G��:!��ď�w�Sʴ�}D��n��r�a.I������Q�+��e���/����|L<Q�[�+H<F����鼇�L�D��2^�.�ə�ft�@9�eT6g��}Z {�w6Vۣ?�_�.�0h�j*�vV�Tw����Ѿ4��`ji.e,4���F����, �F-�Y�O����(t ����:(��c�C!:�HS��\�X��CЍĐFI�[��+XYF7����l%��ƇJs4cX G7p��1ң^Xѝv�����֌I��R`��U2
��̥�{m�/&�|�q��S�Z�+����gTk\߁<�;k@k2TȈ������.u3���z�2�2M^
�*d��4ϲ������4,�"Y^?��t0��E)��]���je�KÆ���}��ʔ?)T-�&F��t��o�;�(�
2*ُGR���IB��^~�̓y�����~�j�HZ-J�����c*��n�.*L�������tD�WN 5�,^u�������U��gujB�m�홋9��ѕ-���1�RvN���,������`9X����J���5�菃u �Dz��B����N��Ǝ�I6��RLVX����|@{��+��a��]�>�^Dz�:�,�i�䄬�f��|���pѧ׆'�{ z����-K��y�dOl���C�A�JV7�.����P�rԱ)�ŉ��������[*�w�֟�nd��F�3�l��^J�n>rx*�/�7
@�"�)��G(SD$b�n��l����;N��(�F��UTY2����246^�ǧ¿���^qNy8�B9���K�.Z�ۦ��3�(.�).������j�e#���%,��W2�n�0��O)FP�����'�Z�7�8t����u{�N��n�l�+iZ>�H쒱�������k�S�_��a^��mJ��rj�/"j������q����8����fY���#4c8>��� �k`sS��U�ce�wг6Ep:S��?Z��˪���c �)E�&���*"Ȑ��~W��Jاm���\��^|�m��sxX:�}�5�c�d�qz1�s��y<��(���J�D�%)�E�"@��`���kƍ��9�X[S�+���"�c��hOe��Q�
�{/O��SY �M�=ϵ�5����R��Q��V8[w��A�.���o�ŖS��(�����lvtxR�5�����ԣ�A����%��pNU��nT,:�����7�|���OCK]Ѹ�r��Y1i����������G���w��M=��Xba�r����%U��]�M׊�\��Eʐ^�s` y�fm�V������|�����nܥ�q�&W�R�q�ku�$-�*��,*�l ���/��}�QI|nz4�g��Qm9��%�B��a�f{�����3��R�j,a�:���z��s4!�qQS�Y��`�Oɷv�$2�Wǖb�G�I�ᄘ�@:b�T�2�O!G�{j�Fż�Yq[~:C�P��4�D���v^1�Ԫ �O�7�Gb �3��+��>S��K�5�ڂa��07��(����hh�4���<�j�%q�+М��i��L�sp��*��6?t*��v7ٓK��L�L��j�X3���-Ƚ�a3�@=�Ò�n�$�.n���GZ%�g.��S�e���Eq?
�J*5��M+�U%N��3�ΘH��q��%h���GY���n����))����>���x5qڂM�+L?Jٯ,|�H�N�}��#�襺y	٬�F*s神�����`���@���TvR�:�w���,��������bi]�B���d��Brz9�$`��0��t����>�]��W1��X�v	�Q�~�&�!-�/��>O�"����k�C�����K�@�����?���0^v�B֩�i����?y�v\�ߞ�_ő��	��1���v��~�	iՖ��nj�.�Z+��?�#<�Y*W��[�hz���;�����%����@KW�Q�*oDe+�r�yk����=V�	����)w9� ��;���&������e�U�9��(�tE�F�UY;$C��6a��;�6�7����o�@��45
]���4�)�;%}ӹ�`����+�j�zZ�T�7��"j��܋����7]Y�b?� C����up?-�dD�x�)St0;,{��8I����9���
��7{x�����4Ө���a2M������E�1� ���@��sx�Y�o�ȩ��֡�h�R���e�*'T��4ոjk�Z�j*��n�6��G��z�������o0���=����S>��$��o�+�OY�G�G7&���!���Au�pW���(�@��rE �\T�^���6-M�uq{|}H���ޚ��4e""F���~n��c�h�Cl�=�W-0ƭnE�tǁy֠G��J���-��tX�U�-��`�9��j���(���(��Q�ђ�o��}�0}j�+`��<cv˼B"��LR\��<���N
�+m������r}�� ŞY�����t ]���Pn�֜>s��	K��	5�Aч�D l!�zpa��´Y��A�`��?s�xڂ��R]ΤA��TK�V����@V��a!���25����NL;kFW��K-�[f0��g0(�)\F�x����W�t�_��^"���A����������<�0�d�r���&��t̑�`�x����k���JЬ�S��}@�����htjແ՛���j�4�W�����َ*�=NP,��TP�'�ຝ;S'�!�]y\��;P��%g��ϼGd.�k���A�J'oN�-z(t ̫��#U����,YЎ��S!_�DaR��k���i^/@��>V�b��'�R�'�83�v��ay��wM7&U̮xt�����S��5d3�u�[c�Rv欶�PG?��'���f���vn�3Ľ��,մT�������-{ԇ ���i�J9��Oq�h[d�m����W�:.�unB[�F�n+ͤ2P� ��1{�o�$/�0�\O���J��F�On�`�K�Ӷ�P�0���G	˽О��Ĵ�9P�?Nv?UҘ/��u�6!O�-���Ca���'�B��������M��c�n���=H�:��D�� z�|:.����@3OW�⪮R���	TJj>9���ĤG��r	<Ľ��xgv�z2��n���E�����z�#"j�{�= �W�������km)"u,_h���hSK^�%��k�x���Z�'K׈l!�[���a��!tV�L7Wy�ce��M���n}�b^|��H��b�0�Q��cu���?�͑����M��gpS�${�MpZ��/Ug���d`3�� ef?�7MZ-	�yyh&�_� �jM� ��#��s�6z(�+��Y���B>��|���Nx���V�CH?���/]���_��5�S�l�D�U=�DMv
(��p����᱿���|zLQ���c��#&�>Y1QI/��Z��*?ߌ���,0�ެљ�>O�[��AYb���뇷8m7�)�,|
���B��Fq����n��p5 Rlڤ�<�������X�44�Ɣ����hA�}1&�r�y�����a��~�����b]p`i9:q�i����	�p۲.h�o����M��p-���sG���u�Ƅv�33�4a����;B$%�ڟ�˔�dj&d���hG�)̅�s�ko�6��g���:�ϓJ�w¤��{�$�)�0�@��>5K3Jrr����ҏ3�1!21��{�Ro<i��}��<��wUI&u8ֶ��3d=�E��O�ř�9;`+':�R+�"� ��>h;6~s$,���爂���k�t�X�^YH,	I�A�7Ik%`�V2���!�!7�`X����8]K��.o�h��4⺖\���2&�S�T��h���.�k��0[sD��ilJك����Bd�5gq ,�(%$�c�oO�ɚ�ɡ�K
��[9DZ�����badż.9,گ4���I��y�A��B�P�W���]ʆ�	Ƴm q@�$��s�dX�ș~�<$�6ؾAn����P��U͵�8��
^��Y�sm��ވW�d;W_�[߬���օ�%l���s5]�S,���w������4���2���,D��Q�cb<1E�Cp<�=w)�=Y�$�A*��r6))�1�f�k�4�{����+i����QRbg�?E�퀦*�lHju��K�8�׿��m~l)-�ּ6�ߕ%t�V�Uaq�o�i$
��7r���YX��DV\��K��RoT"+V[��\MA����rIb~%BQ|	�r,�`�J`z���(�6�]G�N��Ψ��B��!��`�2y$~�������^c�JF|�N}��Jvbru4��E|�}��l]�6d�7��بLs�<;Gf Ȱ�MK��qX�<D��0����-l�Vۜ��)��[�l|Cki�?��ƥ��Mo
���S�x.Qκy"��0@G���(�yq�3�d���Qr��0U��8�<ԑ�h0H�T���9�eX���޽䨕ӫ���/��/k�[j�ӡ�wmS�������׋G��i��\�T��&�H�c"�7���87M���S?���D����C8�7���/zM���f�0�"k�7@/k5�-i�`�5�A�q�r�2��&�+�b������������㶸�\�9��#S��Ȩ����C���j�B�ey�C��^%��HY����s������a.|�aP^N��a�QNV<�v樂����2m�٠���#�xj�_経ޗ�������޼ �}�ˈ���,8�/��M�?�{����݅�v���C ��$LAd�E;c`����c��U
��~Z3܏b�g�]����;�d~��l�'�m�ϣzHÑ��R[J�v2d��F
Ս:#
��u��O���Ȳ#�C��Pr��5X�s�J>M�Kb���S� �_���fc��C�Ði�=��Z�ǰmKT����I�$�I�����i�Iŗ��:�4�����?�����j���1�W.n(��P V;�!��,o��<E���Nl����ƃ�� M���"�xᢧ)W�c�`|�ݘ�VWM��SA�R��y�l�K�#o�~� 4ı��Z q����Gݡo[Bu��N����=�S.r�PDڊ�>.*#�S�H+w�!�x�=L���\Jd'�Y�l���dH��%�.1�(h}l���o)j�o��&��c�ц�Q>�8�MUZ��cX���),� �<^d�k��
4�'��cU�D���F��S �5��~��A�w���
(��ܷ��O�Kf�B�PrioJW�-~����V����L���CX]|���=Bƈ�|Q@�3�`R���8H��re;0�M�썃C���p%�J"��:�����j�&'@$龡?���𪖊����z������3vxd�+8�J7,��S��kLZ��,*�(RY>�(�U�?��[�����pbp_�N��� (s��'�ߵ�-��%v�<3�ܺ̩4�$ʎY�C���D/�O�FW_�� ˿�����â��y�n���Qbѻ\�`������<��A�v�ށ<��dy��U������DE�Gg_8�i"s�f�u� /�%x��^��)�Ap��-�vr��_�����)��)P2r*	J")�?�e�Ip;G���R��v���,�z��'F��Ip)����v�2�&m��Ha"�L7�>���`�t�H\J{���M�QؔDQ���s:�HA�u��E:��4��E3D������M�
5-"t��S`�8㪣��Z��E�f����:y"(�檿�h�\~k3��S?0�2��ߙ�6~�&�/9 ���š�j�[�\Q	��u�?����r���R���F���h�	PG.C���61�*	c����a��.a����^�ApzMC�r�Xc�����G��j�د�����SzU��pE��5������Q!����G����r�u��A�˝�\1�.�� a�����E �^E)ҳ�^�ћ�.��VU�����_门z��<��߃+_��on��A"��M��4�m�v���UQ-����i@a��3��N�[YA�yO$�'t��Nh�B@�NM�f�#���O�VGS�*��l����SN;�طA��Z M�lzd�<0�����	�X��bSۡ�bC�5G�8"Eʵ�bE�yQ����9��J�;Q�c�H�żN�F��;��܆Y��ij�0�;�� �wl���$����!��u�V�kx���K��s�I��t �:�x`u��[��Ǳs�p�^>Ʈ' �t���§��p��싮�b�c�p��B\y�Q�� ���dn�ϥ`{�|��W��|�Y�ꕟk�Wi��%�T������lF�#Z��_��:�ֶ����&�:�M�L�L�HS�����h�0��ÏŴ��6��n���b{��������&>CQ���h���۱�%���@N`�&:��{���N��XÄ2�@��KhG�"���A�b��3���v]�.
�b?W��������=��}ܬ�Qd�8�Y�� �x,��������9�H�.`4B�� ���E*޻����߂N��t1�由�Їf�df)E�r���<HnGT�X��,�B�T�F�D�I�iSG�(�k!}����i]Pd_���nޒ
����kS�,j�CK�5�U�k�^>�ǘ-@���f[�؈�� ���sKB��1�?�z��v��el��3d� ���Q�<&M��됤��_e����"��ӐB�O����,W���y_�z�}��B1�[��*=��v��eI�q��u�V?>sq�p�IR��_&r��,Ue�ŴzQ��\�4����T�*�^X��T/5&��V'�?ā�������>��2&YXQͨj���A��=UE���[�g�K�M���_�M��OL�X������΋��'0=���+����:���]_��+:�Ls�[޾�X�1����h�����*�D�n��$|%�+���J7�%�����V��d��MM{ۀ���5+	vU���E�r�_C����=���zUƄ��|	u�5�D�I V;�_ߣ���'^��6�m�Q�@���xH�Y�cS�e�)�E�ۅ�
#���XF��L�ے�B�-����h(��ͱ���'w�>ƫk�[&��**6�1V��6C�Ӎ&�c�[�Wg���&�� ��j���� x�b���Oo1ҥ���}:V��[�>)ؔ��9���-�<js�#��[[�r[Q��L�if����z0�`���9E�����bF��I �&&�99��PϬ!n���Ks#Q{�<���닩Ñ����)F�LB�UƾM	L�+��߹N�ku��3�R|/k �޶���\��2�H�}��>o	o`��S�T���r��Pd#�zd��z�5c�`W��Rt��?��n-���Hw�X�n�i�����/��D7�(��,-�̝Q�)9Z��W��`5]e�3JQ�M��H\��궴[�V�������=h
�(f"S�]�4
���Ǟ��~�������ɀ��\��`���u$�~!4�gM\?2�`_bzf|�(��K��^��:l�Z�7�iݗ?V�|�	b�Ӣ�W+L���O�z,���j2f?�``�Ċ��v)�8���Xf��mk
~UZ�Ӑ��'#�,�=y:E�D
(`�Ӥ��o���O�W���	dj�AE���`s�@���j�,�k"y�IR�AW :j* �k���� �*Ъ����y	��T���0H��a����ֲ��ϊT@�TN�`�kk@��N̟ΈV��g_�Or=�sk�_�,<���).FdB��C��YB��6��y��8�淚�Da�Q,�_S�ίt���.��I�����<v`f�v�G��0V�7!�
�ʚ�J��?&�v�UF�J�d1R�"���w���[���w IY��
!BA<3�o��/f����6����l��b%���GEl"ƶ�5��Zl��ئ��	qL��� A�i`*��t�o,��AڔE��0淴�*�m��֘�U��pQ���B��J�G':Tv"f����WR����$/^@-�۽Jc�fv�'��3�kM�Rp=����\��k�xB�@��7&����-_\�a����]ҳs
�zҺ7����u�$E'�j��
���l���P�$�{�=?���w�y����]Q���!0%�d F�ԩ8�;���	R������g��\޻�k��c����IфV�,زs����!'q�>ڐ�Vp�2/�UF@^8�A�q&x���*��Z�#��_xN�yM�;D�ܪ��=fFT�����27���qK�^� $�l��x�;'<�E ��%�0�P�Y*lJ��(����m1ޫ��c>��L�UK��97bV.����ym[���d{D?����./s�?~,�0�R�Ƚؗb3�("ׁ]y��2rߘ&*�/<-�|�e��A�u�%�
uK��'9bb���%�^m���Ѵ� ����啰|1�2���ך��zD��6�� ����oE�cg��}�Dw{(�SH�y0��RvA�=�Y1Y�݅�ĝF�Ƌc�=
���pE���ݫuZ���L ��R|��&�#����9��5�)w�g �ϫ�˼� RC�h����=������C�헀�I�h����E�cjD�L"�o�zgt`�!|(���(���8����pb/���@�C`�d1O�����j 6s��+j��X-�v�oQ+pCv�Q�N�Q�>|2=J:v���E����f�O�v�L\#q:+�a��}���2p�v�q�oc~+�Haw���ccy.r%<���W�%���������-�23�p�`�k��i���Ӄ[པ^O��PI���w��E�@�r6�BW�ơ�����Ӝ��I�{��P��?.D��L����&�ǈ<��~������9C�hܚpL�m�x\<2�6� Zg�^ٺ9�
:0b���sf���t�۳�Ǆ��o.���@rz�f�D���N\u�Da]2ׂ4����ˣU�V�FĎ_�4H��`W-�@<KI�'��LıJ���X�4�M׹�Z�>n�4Q�m��'��Y�~�(&ϨU�M#�����v{H�������I�'��OP9�L��Y*��E~r{�t���'���2�U��N�^��=�h����?�#{`������f�?r��[�b�FA�ڽ^󦒉������O�,��%53-�Vw@Wr�󠁒q@�v��p�3v($�P#�I�jDm�}(u��e����[���"�!�0�8>� K��#�L㟛�ɇ� ��:�'F	\{ P���g��4M�PH,��ٹ^b�x]�=
��P�~�
��V���Z~������q�Z���c $�r�ħ�i�0���-򳪙��6��8rW5>N�[)c�e���A�N_��Э{؞ַ�cp�N��8�(Ī�_<гK�����p ���N��DK���޿�>O���~�M�Щ�L�A�A�)��١�������=�� �O���i�z��⫟�gB����;�e��������4йZ/�M��f��L	0C��=۫�q�Nj-��5�J���0�����!%n���+���B��ƇO�h�d^$z����67��5/W
�
5w�D������'�8�;�+�On��D������Y�4��Ǘ5��z��a �0��� ���X~sCU��T�@C��<�q��1���h����2xW�2,X��t��X�ތ6�=���(���zV (.�?��ۅ"4�����5�w@�?�A��ջsMJ+A~9�>��/��:ڗ����A������GR+�4L�UP�����&�@�_�w����C�g�'��<�1���5ݸ�#��#���*d&��Y�^ ��'F�<?�HGYfI	+�S��iח��(qB����(�#�c�j��s���]�CǍ�d�4eb�!�Iѡ�cME���,}	)�d$����Ҿ��� ^�I�w?{l�������䞰RQsnEL�HD�(��[�6k�{�����Ǣ(�)�)�G�����lh~���wWn�D���$�`����!��:7Y--/yI$o�t>��ݫ�E�ïl�`�k�j=^�-��6��*Uz�sPK����ٓr3�`A�h���_Ch���ƨ�U�P*�i#y�#n�pc,��:y���)�r��ƫ�1���`�r���|����w�Ҫ�4!2�,s���QV|q�fŀ(���o��?^��r}��5�᧓��ҩi9V�O�[����-�uj�#��S8R^}��*��{a�����.���)j]�j@��lWKq]���C�Y�d�s��d��F�Ǿ~	�d��W�#}Ga���]0&z؅p{�;Ds�[ �Q��E�R�,,����'��g���lT%��kCuo���E���5�O��������|Y�㟏	���5�lѷ;���zS�"���?� �7p�,��Q�Ӵ���#�xRtQ���4ڸ$Ý�	�e3/=7�HiD��ɛ���N?���hf��/(��S�	���p>����J�H6gxk�H��O<_�e��ǆ�gZf��Fr=����xElE6ֲ�vޭ�
�rY��[%I`k�nݧ5vq�i����X�)�1�0B�@�qs@��t�$�����?�6b��LUx�r¤��o5~��8U��r��"�*�����I��v�RE��Z<�v���dO�!�HvG"5=��n�M�(�MQ�E�l�l\��ƛ�������X���y�� 4n&�s�`��k�R/�3����%�%������okMġ���b1�%���������@*��}�!���{6bۢ<�-��"!E��mI�a�E�NJ6+�b�����$���Y��L��A�u�CM�eC�������7��׃�w!��;��;j��
j-U,ć[T=�):QBv��y���!ݳ�n�ϝHb��uN �i�n����d�拜�� �j�XV��&�����U�0��[��ތ=pCP�R.�$��u@�G����}���n�
2���4��R�|�����a�We[��U��^�XO�Yº<=�c��)�Q��,)x!ѻ��
LIz��o�sG�������`T�4=��j[x�P�Y�֮,�N撬2Y�1���f���DL� ��z_��]����W�?>�X���1����2o�be�^�,�֫�=��16�%���rP�?VC�J��z�h�kj������a�M��g�m��Q.A��&x���J�'	dn��^%����1d��a�`�}��U+��?�2�vݑ}�<��υ ���,"�ˌJ{�5�����/�HK'�%9 �<��6 �5l%��C7�:��UjR�*�&�$d^q3Z��"�,s de �P�m�bں댫���*�ɏ� y�Wd�i��m<��y��°L�y�́|�nċ<e)�J�S��@��/|S�v�vJ�Ā�'
��`��o��@(�Ub�a��:����U���~D�6މpJrZü��J&[D��G**�<����+r��G^:T(Un��\إ(?���V�~JG�yH7Tl�n"�}J�Lawz�w���VM�J� �X�����������d[}l����7�Ύ!�����≳0|�E�T��6 h��������:�9�l�9��G�X�S��L�A���ݕ����IC��{�J�#��7lH�����P!��{�
�L�Ui�ר%1��f�V�df��N�5�g�9��z�9)�Y�W0�u5��I�Qj%c��o��1�����ƨ�n�DY֪4��ʹ� Oq�!��?J���O�?
��\^��^	mhLU�x{��%b1���0n�x@��ѵyx޽܄A�v������+h]�B�
��'�H�ȣ;�;1[�l�9�~�tq$�Q��Va�܌Зs��E �"�yI��B��>> �P��G�b�����ʔ~y𾏪q <���<�bA����%ָZ�&Pį��յ���G�Y��u�o���rn�ڞ�`����k�aߋc{M�*:�O�_bDe�L�������k�`Գ;sG�~[�h��T4[�
��Ô�ަ�6�з,���
�/l�W�(qw��5�pg~��:�	���ܖ�r�_؋R���QLg���m<|u�|�3¶z1��H�/�Ri+/�#4��05��+����C>^
�AP� ��5�}��J�Z��g��CQp�pw�VFp�ܵf���pg�MJL���%olV�uMɮ��(�7�ҁkhȒ��Z2�Sb�`H�6�`͔+f��_��+��H�,iS���Cq�\Cd�G	�lI�� {âz�v������w&�y�շ|Vy���o^w��7�36R>��3�J0�٪��Gd���.��+���y��"�����h�d��_ۡ;.!�]�@T��sѮ>�.�u"P�G*j��x_��,]=����i���0���:e�pLB	pՇ�����EM��9��Dv�9p�}.�7c�	|t�p�D����@�X�6fJ$he� /�S����B�5m�����;�
���r�P����n��7��E�N�x|�L����<TA
���=)±���'chy�;�|�Thǯ���
lZ�k������S��bXc]�����%��"�i!�7Ӛy�J�`�e�j��EB�/�6�щ��&f�?�������q�+j�鸝����-sr��i|�]�}y�:w�C�Qq>i��nJ�c���BP��a�qO���F���Q,���}�+h�4�Aó�2�V�9�{�����o�?:���Q�
g_�(�?��2MH���K1�e�!���s�Z�ؘ���6�}��(���*/����7Ji����x ���f`#.ܻ�E��<u��[[��a&�#���m�<\y�s��UE/Mۃ� *- =&)�|Ol���͐��ŵ��������b����T4�!߻�7P��YyM��ƟsZ�(�
�� nrz��7����.�������z�/R�����w���(��>8u;Xd��(���37�q�n�C��p�]��X|�6aCbY�i���G��I4���hM� �B��'Y��K	�;���ԇ��p�������dN:My�o*�`T��W"ms(by�á�f�L���Pu�#���P?�R�3�u\T��I�W[؋k켮�|)%�:∤$͑Z�V��*B��-���2	"�=݇Px�`"�Z�W�.�J�S^<e�49K2�phw¨^���v�3�[��*R�*��U� �9��Ha	�F��CH�ٓ
�ay�lĭ�n7��P�\f5Y�U������bA��4�(i��E*�7-�MJ��aW�C4��ܱ�+�K���o��]ؠ-�*�q��'���1�_-����\�)\Q<�|`͊��	z}׈�|.��Ի��`���F>`�M ���S�G�5�XF��������B-o>�~NCUaR�|s.��	�/�6��X��wܔS1��d}�'zЀEO#A�9�dRY��.6*�:!xs�I��Z5@���v�V�X�Ֆ^��l��(	��Ab]g8������8�|f�����n�]�lWB���8ΉͪJ�~4��/�b!����<GO���?D��#��Ԯ�R�������t��s� �Hq�`r����z��q� Ϭ=G=��F�乯ݛJf�S�Р�>�BZ3j`��d`�ö�'PM��d	�����ʴ�"��V�YXE�fc61�;|�*�Ru��骇q}�B�����܇?a�(�"=�,��3�-�r�z�f��O�O��%��׬����Z��I���_�U�����.f{!�d`P�ȟ���Q���\&j��GX�P�e7��52Ɨz��{�)��\�D(P�ס!�ۡ�s�p
"^��8���C"����#�Lt�4�&c9�!d��k:��3��*3G7�����R:fهh{�>c]��w)�t`�x���y����2�੷��Tt��x�� �qx���B��J��\p�@�O����0��L��@!7�UZ(~�-	(}=>!I��QCN�L5k�*Ȑms5z<��CZ��9ro�����6=�{wԗ����~�eR YYB��G�B4�����cV%)s�V��B]j
Xi��1$�@`��le~��i����˞�����pE�(�*��4��?C�v&��ޟ_�h��/e�d.��dQٱ�}�2� �'��E��Fu���0�j*����xCv��5���l����#�.���I���J~fY�Ǌ7���a�l�.r@ť�*=y��nb��� �s�y{5��(�Cn�.H�q�]�=4�"��9̆um�T�U-~�9��U���{��Ը
k�V_-p/n��B������ﲄ�i�O5�R����`�o���]ZFZ�l�Vu�U���(��C��Qb\vMT�6�
L�W��ad��n�$�Ō*�글�\#�t@j!��K��� )����\-�=\��s����9�?/2��h?�	t<�
z����D��Ƹ�P%G4O�X�eX�r߫�������vKlUwT�й&y�c_���R.���:<�4���Մ���WՔi��Y�}�NHu�Z���m�ª�6%ܪ���=~����do�=�p@���mo�� I?1�;%��Q�}��b��/�����uюJ�66s�L�(�I��R��[}�G�O�#R8�z����g
f�f�aQ}D�&�N��o�+��}g��y���zvS�������6Z;C4��:E��x]`��, �]�S�y.�S_�a���^뺄¿��Z.��K�!J���|9���&�癓E�7�^���K&9��r%��wiVj���DE~'_��O���G%@:z)d�z��L�1:�U�		zf3��`N���{�צkMl���������������
hݡ��v�GT��k]��y�I}RG�nRf�-8d �А ����P�/�$����戲�efT_�m�����qv0��:���5�8A��|$�R��Ѷ�P>�'���bmc`gV���Y�"&n��'�)b�⦎�H������1�H�6�>�q��+��Gu��^����_ī��s
3T���ʱ�`2{a�*�[�T�(��bU���K�i/wW��s1m\i��2B)�'�A�{��F'��`\1��s��� ެ55���o���(O�,067����o��DW:a��{�y` V�eK�R������$$�Qͥ��7l�^\N����K5��Ҟ �MݩF����ti�F���<6�ۛ޾�P�-�f�W��e�]�_)n���
��趾���*0�}�qTke�_pJ�U�&��G3r��Ka��v��N���s���0�X��_)�f4i�����aDt!���^����cz�^��`�u_�ʈ�I���[L\�~��xN{.�i\�C�D�ڑ�t�L���+���D��&R��t���ۨ
^�=�R���x�,�9
vb�dF����\GPp�^.\lj��Q��.��R~R���**��[�/�Q�T�׍�o�h&OI1����񒗷R%���^�9gD~Cm��2�|��^�(���l
��G����P�/6q�<�p�p����׃P0��{(���W��������k>	�G��lU����o�9�붯���Y�H	��OW�I��q��L2��=�4Φ�Z�)LD�%�~�Dg�s�$
�,�A>�I�؛`>}��ŅN���A��YkN��r��t1�9�����;��x�vr7h=/��?�@����>�¤jJ�F���J�Z�`��pQ:qD�~DI��n�p�䘈�Sp�Jv��=��8>���6�+/�zq�y����/�����<.����g�ltsm�W����hy�O���z�Z��su��S`�K�a���ጎge�d{a�����5^A�&6I�Ş�M��3���f��	a/�H[<�8)io�)��>'�i�&+���[=��ڦ\�Nf��;�x�
 J��:5����z�0Cy�F��~���2���n�9�S���"iO��q����H�5`~�;@)�B��Ǝ���u �E�/��J>�f(�,��A��̙�TN�p������B#o��S��pw�5��+W}��*��g�u��r�� ��������o���>�ݨG!�)>�c<�5�y�s韮��ǽ]�(�������s�|v��8C�e�(CQ��	q!u �wmF=��`\>]�2��v���O%[�
6�,�`�4��qV��&��Gn�Z�1l�����?\FC����hL���v]���!��d�kA����]:$uM:?����l�_����w!����_��䗫E��̋\���e�Hmh�.6�.d��Te�H�Tmc�N�S�u�����g!�#N��!^7Z��<���љ
EbB9�V�?�b��N������.�͉�L(��������k���if�B�>�o�0͹u������d�IP����p��Y��@U��ֱ�?^��94 $VزI�`��,`bN�)@Q�O���(�3 ��ʫ��ѷټ�,�^&��ӄ_X}���B�O�sK�]�2�fW�k�^�ȅK�r�H�t��j���vv�ˋ��ۊ�$K�ũjj�kn�U0 ��IT���a���տ9�Dȧ]�;�o���&�h�,9ݝT�_;��c���7=��ͷg��!�ŋ���p�vTyLD���.ݵd7"��M���oi�v:�%,�}��!�_��"���uS�[�����B���`�L�Ã)*B*���
t�x|������o@�������$�$�8����Dz4[!�}ؚ�6`�|����4dM�	NIO�V��x�H����&-���҃ț���)�ꀵ=�-�Ġ�H�����ϱ`�̜~=L��%��Fa{	э�Č�ir�YUJ���;�]{b�ڒ�|� :�Լ���`�c�E���&_sg	/e8C|��Mte��H	��^dXW�ǈϿS��(h�61�Cn���W�	��0`5>��N���#~:��BD���ꉌ����[�\3㪺��@�G}�F�E`LV�>�*��-Su=��A�[>%��\+n���,����:?�=%���vI.��-�0� \��{��<�-��]ŏ��)��r�TrLx�/{�|U����<�_�� h�P�ocQ~�Ǳ!�.�*���#d�k�j��t�={��)1e��"�x�Jfʮ���Y���x��;h~�LA���|1%�U /f��9��Xl�`�q!^O#f�T �#��5�a��L�`%ObtO0�"E������j�Zs�D��(�Î��J��@��s$�����[�}}?���+���r��%UI��uͿ��o��E����ƭM���̅H!k�D�},ȓ�*�b������;����8����i11���RIR+��Yp�q�wH0�U2}͇OӁ D�$>�sl1�'}�֬��@(]g���"����r�q�!�6�^o$)2�D�*�C�C���L:�s�e?1��Wmg�{�F@�	�㰼~�K"h�rJC�Ӊ�����0����s 1-,�^�s�īn�B�.k�}G�}r�Sh/^���聉�a� �+{�E�./�B�2ޅ��"�0#@����-jZTDL���1bA�������9[����^-.Ă�5����2rKW$7��s���e:���C�5����Ŵj%��K�������e�G�m{}�J߮�m�j$�wo����~��ii�����5�9��kH!k��
m����7;�T&����W
�c��xO���\e~DsXu�|EZ�X��x�f� �� n5�"����ԮQ�Z1�[��$ޭ�^0����������20L�Em}�Qc�t[x�3�����<��x�����d���v���|�ǐ1��`y	{ٯ���yC�)�,M�̺� ��N
60e'�����t����j0L�tK�/����PMR�&Uc��L�V=g�oa�6�o<Z6���V-� ��6���IL��\+�v�tX����R�UEʜ����^�^;/q��g��Nu���
��}2�`$�cf�����ц�<d�*��e��i���O���[.ŵ�{e���w)g�%^� .�m����~��@�>Ӈ��ϳՅ8�\�|�BSR�
>U�Bfä����K�n�q+[���(�A��K�j���m���8���a/q����HE�m�������	�,��
5��_�^-��G���h���5Ymz��j�>���6�)�\�RC���E!$��ɓ�?q��1m@�����w*��fйY��1Qؗ���#�,q,`(�}�2Vl��7ww�R@���i��QL��Ҏ��ߖ��H�I�E^'e�99��8��z*��\��T^�n���Ӄ�i����DE���yt?5B��rv�<e�-�N^}���*�I�S"HK_��a�$=S]���YC���3��i���O��d���w;א�����Y��r��5 o�����gq��,b�C.b�ej�%����f�ƍ6Έ��Fa��x��r�[݇��V��Vy�hwK�{��z�:���mN��@�2�ږ�����jްSuP�56F�����6^�K���c]@YR�a }��a�",�̮Ss�vG+�.�]�x�J�M��pU0���Հ-��/����d�|���'*\��5�����*���@���q���Ξ%*w����[�6��c��
ވ�{���
3d�V`&�!��AB6�L�8y$����+\���)Eڧ�C�Vo�a߆z��v��7ҵ⏟�*�m�7�$������Q���n�MB1�X䑕\�7����K��ea���S�1X\��oq	��N���r]����m��y��d˒��W�/��g#z����0���LΞ'?�h�;�;�k\<�X�y"�0��B%{��&EI�c�:�� ���Gq�,�$R����0Mm�R_���E������B��&K�_I<�;��� q�40�}I������r{���w�*��*4�3	k�R=l{�og���
��=w�#$<ԢB�>�����z��h	����2�Xʧ����-k�m6��jn0��'��y�q��L�;F� �
.�=�5AB�7& .��{����rr~y�"�D�gpW��`U�5��˷l��b>q@�����S5H�z�Da�X��-ϑ���^�m�3Q�1uXlt����#?G3�8��ʖ��[hL����9@�Xr�G�a���B4�ʻ�<��b���-��r���2���Z�"l����Ǿ°�����o�x�\�_}�Q���w��w!v"������b���U}�f���|�~�Q?:c;���*CG%!$h��B�D!�p�H����w�L���'˵Q>�x�Q(��g� }�	v�_}�M3qO:��,3��[q+�3����9mSU�%kf�5zf���MU�S� zj����;��\��v��4�t兕ذG��ʍ���=w*60h��f�;'���7�t9��(q�9�Fʨ0�ޅ%<�*�}o��(k�tQI�t�L�
&cPk���i��P�~�V}z��I��&/�2yR`H��IV:%���X4��m�|r�mj���B�<�^��΃�7NZ{_�dֈt�$�'���ز���W����%;��W������_!x�� Ŭ��_�:�Bڧ O��}��nގJ1�J��g�Ր�4��?�����0����p����a)��|�M��ͫ�R�*�K~�+���3B֔�pʜ��9l�0�А5���qxMU��	��i��.�hj�fb� ��)a1���'P�xv���RW��Rq��%�@�N��dGjLv�OK�
�e:��#~'��{]�>4���:�2��ve�/xW�ye�x�Q=P�W �~`������*��c	(�I[���\�;c=ntgd�¨{�.��M�;�It���E&>w�p����u��/��A쩰�<Vs�FtL�3�l7���E�J�{Dm�q����� ���K�z���nZ'�B���ЌB) �t�@����k��E�7q�zxQ
$
Z(�糙�(�������o��"4�E,�M1e�1������tS��k�d"Ug�NvFU�]��I@�Dф$Oq��i�mw�	��9�G�c��k��D�	��&�)<Ȝ*� rh��Q}{w'���"ߡ�{�L��$>К�Q@ޤ/�G�����Pb|�U) v�L�9u�G�~6�ܶ���"�"b����مE���TV�a�N�[������J�8��D�L�,ڌI�d��n191��7.SE���}�)��	&�A��	0���Q|KF�с0���B^�r �?����.��%���l�*u\,��}wz�Hg�Q<�c� �in����"��?��{@�c��[��XGz��a�0UY��_�Ōig�*���Ć�A��Q��^!MR�Y�ϓ�Ԯ!�C��}�����#�c��f�k�uʈa��KU����;��j�i���k��ْ1Cw���ef�y���n��X����I���"�Br����ّ����iַa��*��ɪw��R_�����x�K�%����D9�㨖�"V�F���ma*���Rt�V�z�z��$MmY��Z ��
�Y��޺oG͹>�&@	2ԁ{�@��������=j���~a�#�\����&��C1��Lb��s�n�%M�.����eƻ�rL�pei/�-�����
���o��eO�����2IǤg-��pE[Jnm?૯+���I�NF�&3���L��V^W}�B\&zt�%č�V�q�#�8���qt 3e��<Z�$��3<���P�B��DRs%C�C�������ي}�k�3$��27�'W�����A��;�|�.��y�2����E��؝#h���~&=���v+z�
6��跭�+��JJs;(!x�˰�
���2�N���~�C��z39���"�x[�4�#ԫ��[���h�r���p���y�rPvr����7�'q���#C���AYs���-7����lv��~Q>jO�h~2�
�C6r��Y���U �uBmgf�ų�B�7�<�����}Z�I)*,����Ō[v��ʩy��8�{Qv�/�(c$a/Ec�z.3c�ʵ3r�+NP~�A���G[����C��?]�j͘���Ip0\vTIJǼہ�(9�}0���,���e,��H\�KF��\��h������ˡ~��ꀴ����c���	�������Dol{�n��N_$a�I�������S��m����5+"���Ŋ��I�"I���	{�Q���X@G㭷����礳���_���q�d�ˎ-�3�w�(g+�tjt#�Y��}DXoa*�jH�#[
���0��ku�k
��|6�ɤs�
{���g#����*y>)��k��L+�������UA�7,u�v<Jᅌ���X5j�E�n��%��譡^����~4��I�A"r���F�����f��H�D�Ij�wrC��Op��H'�O��u�y0�5�VI����qϷ����I�,�����S�m�+��ͤ��z��BI�C��`��)�9��%���U�񹢗����Qɪ�ix�'��̀��G���~�^�ȹ��S�ӮkA<t�,v���[#�<�� nǄF���M�����ǣf��#W���e�N2cb6�h횈Y�>Ӝ2X,��Up�	z���#�!�-���+0���?0�6�$�����YӴ��+P+��'G��A����L٪,�Rs~	~�����"q=7��~3*h���(~�����A(�b_��.�9��D�t1:�:R�M��FFv���b�h/<ȱ�Zu%�7[)����f��ݛ�(��Tg�{�/~�=�������+�E�*Q�����_J��*�=;!��(|�;�0��Sg]��&\�る��5���a��;�_�	Զ�v,��m��l�z��^M��I҄��������y�Jz��(p�-�myY�`m�x��w�D3v+A�����<���!�+�g�"��hT qXd>b�ySv�r���c.�DPb��S������q�[z�d~���q�$y�{�@t| ��k̰ 1��d�_�qɣ�O�w	)"�p���lX��ʳl�}Ÿ"muI�
���i�L��5�o�l�B��t�On��]8�GD��s���d��!f?7%n������0��Au�E��QWKT3�x�b�K��Yy��-&C^Z�J�R�<�x��Ut��)������P`pB�������wى!�e1t�
�� >��,�E���\���(�Jw��� �ۥ|D(O<��RM�+��݊��'���;#c,�0�Ė*�M�iT�{����_�C��ϙAN:$�j���EE�H��Vx̶«l��{]R�dUb(W��F��-���"�O2�zi��Ev"��{.9����]���2x���PGP�'�GG2F!#�OQa�|���/�y�3d���2/1�*i!0ΐu{Xp}��9� ���}�th���>�We< 4z��Y�4�ke-���/�޵��*�gS �6��l���ռ���Ez�E�L����đ����4�%�=�_��Q�F�˷4'G9��V-Ǭo��D�)$ߦnTmd]���o��Ѝ�"a���l�L�Ie������됶���`d�-�K#�kbux�~�,�:���������l�Jp���� ��� 7_i�L(�Oƙ�v��H=�QX� �}��gM]�ɂ=V�S29�$��Q��u��nF��f$>�,@�a�E���M2�OW�Mo3���DsH3�	�M�9�ْ�GәB���3H]%�e�i�۽�F��CC��"��]*S��a�/��y�X��DW�xL������g��׷�#�h��yY����>1$廑�ϭkT�w�������Q�qc�����(7���!��<�EWC�s�$XJL�ZYwT�3B3H�����a� �J��?�u"9�؄�M�n뱅V7�+~�C.������K���:2�����ov
F��c]��1n����5�^n�@t�p�~�L�
V!�*k�^b�[�y0�n{��d�c9Z��.���|� 8M/<$��+�=)S� �W9��kQ�W��� ������t�0�[��G��6�<��%Q��E�GېO�r��we<2@ӽ��H�����<�
/ű=أ:.�_<��N�I�>��:�''�3_���4Z-�{�\ bwG�ܕ��|�����^��޾���^d�.3z��4>T�H��e�,
�"r3�Hd�8|�k�Q��m�[��D�:IW�n���軩�ϸO&�|�"+�u�*;uw)^َ����v'� ��G¯g$p{^*W�II/q�G�f�V$@�f�G�4͚gQ�X�`�G3D���`�dEo��AFP�WQ_9�jp:��r�]u���|ѫg�q��-�Ķ��b}��6e����?*�R6��l>Aw�%b����ժ~���19&$k�s�._�E$��+�|8��0��R%a���磣m9��L�2;�oY݊R���u~^RT��'3��+�<=�IHQ�=�M���}�f�6�I�n��&�<��`Jʌ̮T�P��8[/D���p9��pW��a*0��.+ P!>N��S�Ѓ�ڡ?�;	$�ƨŖAu���{�9u�q����&����;3:�&[�D��;F>-1�v��+��&Rԛg���:6����M��%W�,�hrL�U�|��ugf���-���p�D��:􉭟�"^���B�9]�6ʸ�=�����sI��i�8Ԣo������(a,�q;������m�߿b������,`��ykx��y��d�İq�D1�z![-��A��76��E��\��H�m3��n%��If�7�D���!���pR¤������Vɵ���p������Q�@���<]+7��>�x�C�	"+t'�͸�Ш/C'69>�^)~ȦL�����R�3��U��{��P��I�R��{��f�����Uԉ�y���O�V����y��*﮴����qQp)�h�He���/��s���F�"F��&�%�d�+�K8��ǩ3��q?���Mz��KC��~�aa3�15)�]��|8�P�~��Q�}��a���ͭ�%�G�b�Gq�t������Za2�O��}}
��/�L/j�i�]V��k:+�Zԉ��xe��Y_<����S<N_��߱6%_+�����h���"���-K�f���=�Hm���f�Th�<���
�k�gmF���kYb|�Wo3�S̥2��01�p�õ7ڗN�^�#��M ^]<{��.��A#҂ǯ�š�������!y|�w�:ضV7�V��뽕~��������|)ܘ����6�qܚ�_SUR�3�1|��tk�D���N!��2@r"9��c��b���J}�aW���b�:�-N+�[���k��ː�w~1V>�oʣ���/Av�ȸ�}�	A�"����8�6/���n���/|��(�ؑ>��=3�کF�L�x�p������6�cy@�� ���T=i��'��	���Q3�`Y���)���"�1�.6�vCf�M=[���"	7L�,��𿖦�-kQ�r��>D��H���b:�n�� 'ÿ��`.��bQ�H���ӫ�����b�������O�'L��1�����{�ő*\F�`Y��	̐i�p�-�qĈ�"�>��~�>v�پ�����6����3?���4��M���I��?�yV1�REGO>q���_��wbac�t2 ���٩��0�D�X>��6���}��a�$����|K꿍�`�ӄ�e��ۊV�Z,{�O�@*�%Y��U�4m,���=�U �$�]beӉ��eMqH�
c	t����x��wǅ��"v�خ�n��p�> ��#�Os*�e�B�8��=k�*�u������@i�s��d�8���jF�D�pJ��I*�4d�o��⵮��hx,��!���Zfs\��<"���f2,Fi�j �#`���c������ѨS2���杇'�R|B�-L�+�}�#Q�,>=ءs����K]���J��@;QJ��MT�w׏<�T
giQ��ELM�"�����k����٦�ȟ��O�$Ҫn�#��L��X���±�(6�B�פ?E<2��a�%
9ibo���2��+'V3��^Nxز"N͈2p�$�*���{K�\ܘ�)lfe`�m3�[�E�&�ާ]���"g�ʉ�b�ud��%���ocV��z�W~�c���Z���K��EHujL�q::T�dz1F"��H/��4[_����GH�Z+f��&"����a����fun(�0p�]dX<�[�7������4M����:i��2!�Z	9$ې:G-�M�T�8��eE�C��`L��� �J̼/�SB��!D�Q��B8��r!Ѣ�'�r/���L��*��mkj���M~'����8)�X֥��8O��)�<�Եu�C���O��������>O�3�B��Ѫ��u6�s|︫(�B0<�I�uR�S��!�ؖӱ�"�W����ﰪt��<��Ѫ/���o��5�����e*		"=���)S����*�$������3-偰?���N!}�N��+��w�n�PH}���s52�@�@���I��͗�0t��6_��C]�L\�w������ �8����{�(���g�C햀��+�	��y�ԌVw�"1�#�T�h�v��28k�e"��@�_�~zX8o^L
��)����<>0�O���dV��V�)EUR�v�$T�/t���
�_�T�.E����b��p�#���D�ű�����/ɖػ���K�&n�3K��QŪ'1���'/�[d�[�唴\,Iuy�EPMy��8�qHYxfx1�<�Un1�='���ɺ�pOQ�.zE�S.09 	�8لJ2�#w���+ʴ���,cg�痓���-b��(�Od���V���'<���w(y����G�ޞ��&�����W�vx9�ԐujM(L����wb�.�EL*4m���^(p�k	j'�Ы�-3���I	�v�Y��E��
t��q�����������x���%c�w�!�F����
��hq�ڌ�X���記
v#|2����Q"3��r=�_Ҭ��M�꫿��n��9�ϣ�c�6��J>�/G��Dg�;0�g0��|a����v�e ~�3/�ln/�+�#�	(��p��:���.d�')�,c�>��R�DTK*S�U�C��I]u �n-�<?I-�`ZFqD��R̋�$��Du��e�!����v$����^�U
��)�,��)e>�(�/n2y�`�WO�����|�ޤ�b��'�y'�ĕ���ig��n�l�M�+} NL�X�?�T���� ʁ7�������~A������N�\�<��a�ѹ�sa���}��o���t�~"94�v
.�^?��B�2<űO����!xH����v�6-8Ʒ9dq�{�j*�rТ�*5���e~g>�H�3o�{%L��Go%�^��	$-��0���/�{(()c��\(����Pg���9�5�sB��^��7�����,�ȅ\�Z��T��ƹ�����v�;z��	wO�Z2�8�>�_)�=�(4���I�7f���8飠�[ꛥ�K�U�mZM�I�Ϫ��ܒ�,jCV��aK��U�7�;;��~+�Gst�N�{� n"�W���������;��/����PyP����|R9G3��u��7$`Ɔ�k�v_;5w_���˲*��2�K�L�c��q��X�k8ch�K9��P�IB� 61$����,f�V	�,G4O2/y�\��S�N��������oW�x�� ��x@�b'[A)����_O��y*:0��E�T	�D����g��)�E����k���� <��31����@��`�Q�i{���2�PVZ��IO#�i3�O��!�M#,�c;�h��x��^��9���oil�,�z�-*�r�P��S�*��g8C�'�Y��P��sK���.1�E`�|��'�OR2	���v�8���d7&��g�r��&>=c��.�zG����s�"��v�>��1�{7C�p��Ѹg�`\3�v��W��^��$Қʟ�����U��F�<	�_#�+;������B�q3jќ#��Q��^�+܁�Fծ�x3��G��nP� �U�~E��K�'#����yt�m�t;���W'Xz�� G��rH "ֆ5Ѧ�	��G/���~d��Cf�`��������a�&$���̤ۣ�on��Qi������ �"��ip���kR��PL��V�o#J�W�V�p��{ϣI]�McQ�yE�'�=��9�av�l�VT'��_���|�
��ul|*)�a�#�Y�߭Qu<e@�_�l|Aq'GH�dH�\��J����� �V&�@�(cj��C�!�W�v��	�ì���O��FH��4{�A{���W���w;Miy�Vئr�:&��ILT-�����"�J����Rדּ�~Ho��Ê��/Ҽ��\	6�Z���.u��������6'���.R;|77M� ���L��i�*{sxT�y�o�a�T�D�hfht\��>���2�2��Z:�j����;�߳������5�z���Vqfl�=c�W�Ղ�rk*�rI�zXª�s�U����p��(�F�}�̎m'FX�����%�Li�5j�y�W�`*�A{��qs�-�Ai�gqgI}Y�7/N ��j�*3�.`{����ޚƒpP#F�1�6��/]�?ۿh�>����d�?����)ZY�"�M)h��E�c,v�<���
���,�p�=�"`��m��LT�G���:��Σ��Q�]-���{$+
O���8^��+��`���ۃ0���F�kj�2g�nx4�M1��xV�����Z�!���r�my���R!~�r��3�=�!��6���Wp��d���$���>r��sdj�o=���e�Mc�*W�_v�M������G�&��C�h�6�iU}�0"�`���Q�!����V�#����S����MQ:���禮����QZfd��l�����ݕ������xQ�z�x��\�,�1��C&�=#�R�m{���ʅ1��_by�N@�b��}�6c�hm�X�:��@��C�|�����7s��fY�_��[�x˶T,�z��b:A�%'o/���l)�;q�"!��,���b���m�%���mE`��h��.wM���TNx3��Z��u�y2|���1h��BdL�����82t��ҟ�~��k"�.��T ˘�28�V��Pƶ�ͷ:�~�v�ĨH�
���"��I��� [�`"_��1ĥߔ�]���/�z'`�����<I�� � ���ӵ�ӗø�Mد�}�D�g�F%��;�+@�e[.�B � h��bE��Wӏ�%y����B����x�e����=:[�$C�g��}G�դΑ-ŚщUgJ�i�6��4B�o�6k���A��"��Z\��D�hwd:��n͜V7����-,�K<�,f�Po �b��ѿK�Շ�r�@čW�2���p,OM�9��L�񋔔�ysm['`w���2�d���8?*��p��1r����d�[�Wn_���QR��m�:�TU<Q��%�K���y�����T���^%��咙]~�A���x��8k�N3Y���y�e,���}��#kq�Z��w�&��yF�CGmipĽ1���qe�~[��rIݡ3+�BE���6�lG�̀o�@�[��n~H�օ�Ih���.bA��V�~��^HA�(�f�������?��3�� 8@�˄I�Q�p1����ԉ��c 6����l���������G�e�<�ŕ�r�&��U&\+�)�0I��i����� ��v_�I2�>�J�����6a��t��vؾeY[���C��E�R��f�9ݛ���Qy����x�P%d��΢�bX_��J~f6��ZԥBz�c	�y��.%_�H��f����i~���Ұ p�RX̺��B�=x�Hg����q�{H1P���G#Ǽ�?���2sJ��Ao�N�n h�t��#\�8�[mע�*:4gvA��ߐ�����Wo���1̯�AL��P�I1�����hk�CS��ث��5�b��ʿ~�-.�6�܇�+:X��w�Г8�L�-�/H�22)��^=�6т��7A���t'�I�XO��U�V?�p -�f���
i%�Q�AD}|&�7�Җ	�ȗ�Q/�?1��,[�������X}��K��ҵ"��F-ޛ{�}��X���~$$���z��D�W������E\���/>�PT!jK�����R���qZ�� �U7�t�n2��n�s��c���(��=��#�������y{	�^\�K��kx������Ĝط5��?������P��~┘!6���ɺ?M��Eo��~+�ۣڳ������'������5���G��D���_긷f��ȁ��IP�Z�{�����u�s�|�/�XlxW;h,���pj��^殡M�x.|3�%S 9�:)
f>K�O��V��s�@ � y���\|���)�����f��;�he������O����]��Wq��Qsn���;h�	8	7���N���?x�q�MA����b7%]���lb�T-VY����Y��6�� >�>���E���V,F�'�cM˽
�+��O����1y�^;iU'0W�x�~ڨ\~�!8wX;�Ļ��Uy��������(�r����M��@�kGf ��*��4[�TK<�O	7���đu�`5v#W�T��g��FEf�5�{� �7�VYz�$����gX�`2A��B�
j��~y����8���C�᳥6�?���Sgb�0�o:�g�ư����� [kt"�ژ��J���>�f�\^"�@yw�y}7FX&�6h��2.���<K���Q����P�����v�\�ZX+�r�݆��MhŹ��P��l�5cWI0M�r�K�i.����=V�۷@�_�s���U]�plpP7���$�������Ǻ`{�B�Z�uliLu;=��🭧�VKNM�m�KIK~��7�;|���Z>|1� I���9'����Zt���j6O4�昱Ń����Y�[x�	�Q��&�G����O�@`F�׎ZЎ��B�h�Bp�+�A?�[z������b��Ozb�pO����XR~ :]D�SD�\U���gcZl�u�-���5���i(}�����cW/L�:���I	�����b6�:�d�I�樫C��-2���O�_����:7�~e����1�L���u�̢V+�
&"���__�:���׎#�STG��/H!�ѝ��3��r�Q������u�����%��?�N��W@�l�)�����a_�p?V!��@�x�&� �
�w�>N��&a��*����`�t���3޶2q�n�w�M�Ed6�Z�gLZ�J�g���y�.ԶM3���v=R{�m�f� ��~�3�� �G����n��3CPV:/�NR�h�T.��8�J��R#�I$!>��v�x�}������_xJ��ne�e��帠Ȇ�m˦��x�+��N�"���x�#+��QW-�=j������t��{����rk/�-�z���2|P��\8N.�w�� ��*��̎S�����wac>?2�moH�,J�)ɗI�0LN.�~3WK?0�u�����>�Cl�2S��~a��ܯo��OZE��|-��ď罄
@�OR��<)3E��y����~d�^�˻�Q~���Φ,���/2O�WF���vwSbn[��� l޽,�Ssv��l�0�&�� y�����q�y����% =�7��]X��/*;��0p��3o�#��(���n+w�l�m_~l:T�T����sgC!����=������U��jxoL�lBtl�9�줙5�Ӆp��C���l�),��$�F��R���0oa<Hn�@��`�v��~��d��sYE��)���آ�����Q�J0��;m\k���Z8N��������h�;T�CU_ՈD5�.N�}�y;���4���V��͡�Fy�<�
f��)P�/�b���c�B�
�p�W����u���wU�x��U���%�6���-��0ۿY"c�N`%� ۝_���Cn�[��xp��z��F��7�r`��v���(�9(�N�I�pCͣ'|ı�3Ɔ�
���X�:%��5�*����V�u! �s�X6ojg1�ä  .�\pͩ!E�Mq��m4��@�@F*��I�jx	�rvդ/�z��M�8����F5���Au�C�O��������W���
dҏ�'|I���-w�ߍ���U�T�#PEU�[�ܓ��c����m��5��3��(w6omIS;�t�q2�-[ K?cܢ⟄�i� ��_��S�恜��=�-��}���9����BuK�T*�Qpj�QM�]�;X�b������|�o�����u��ţ·���7q��pZx��E�@,�Ad�XK�Ԝ��|�`�#�-7�T]��qս��\"	T�v&�=9Y��/x�[:� ����\\��#l�6�	��w�rR��3�"��'��O�7qi�j|b�K2[8��( �=����DtO��#�q��C8�U���G)�&���/i^MN:��Jq��veU���aG�)�p��<Qd=�N��O�y7�$!�e�a�w7u���ƵN ��{�do*�>3d��-��.���=gCz ����OM����*����^+�x����})+�r���D�;P&#@k�E��3j�t�t$IӻE�̛|��ʃ�5�eS<=���"��Hp��r6�z�Y;�(h̐`�Z�ѕk��E-��_�Х�~�c��ʪ��r�����W��b{xQ]\�ľ�'����`��$<�`����bY��)���)����N<�@{�]�/%VŅ�6RlN�;K��(FF�;Oۚ1u�Y c�r:�򓴢�1���O��h��ʧ���z�+��ƿ*�[�b�j	�ɸ� �b}%�\Z�C�ٴq�ıă
�� Fn�B/��[ݞ���٧~&�έ��?|�%G����0>{�C�miLg��
�i�&��ґ:jP-΁���_�Uf75���2�'�-&��M�,�7�Of����B��@�m�_V�A�I�;�U�_"�l��_W��%���� Cc�V�-�2:^7Y]���P6�u���]M����j�5\���l��3v}�g�Ւ�c>�ÐL]��7�I�?o��w��Q�5�J�u6�;��(��^�Q��� �Q�S�.�t��Ф�lإ��M�#�Ȭ)r��k
z\�F��&B�_��1���&���:�JA��o�j~[#��iI�>���5�����Y�-�a��<T����}�t~��f<���A�w�e_�G�?P���bS�������Z��Iv�[)Zp����]�u�ꨜ)X�z9=�8� Y!~޼�Е�:�v�'EC�`��]=
�|	�\٦��j��}�.q ��ǚ� ��O����s_�UJ)=wv����72���4���PޘI�_]HT͏�V)�/W���z���n<�����*�U����<���|l��5����<�	W<X�^?�h���G����U�,D��}y�ke�o1�|�p���+T4�5�[�A�j�X�-"�{��fa_]'��.�%U��#g`�5?O����^\�Q������nOC��-�x)%Ƴ���ѶWĺNh���<T"sh��ж@�"(�1�?B����;a~��|�k��=U0�Uy���f'��}T
{�?QUxP�+zR�Uu�Ɇ�sN�݂x�h�8P#�GDC�d���D[2�������U�>k�+��gt?�������n�&[���ƲL(]�I�`r"=�*G�=����5[j�$(��l��� �]�I_��U�Nm�[��"�4�gg�M�pdS������`2U��5db��(0�6�H>r#D���˛� C����I_�,�A<Aeu���a��ȻF#�ʱ�dO�8�$�6tQ��e8�r��[߬�zɚ�v�����0���\��%��ĆsT��g�[�藡c��V~E����m+|�b���L��Y.�]Z'�a���ǴM��e�zu�O���}�.ǚf��7��&1���a����i����[��M[���i�!�r�vUp^�9��<��CY�K��������ʭ�����+q1%�������c�B֢3��8_&!�;l#yzG�b���)��ԅs�N\����]���)��pTM�����^�$_�b
HI��Vzf˩"��av𒍂PNYL�������q<$j:Nl��U�u?1#pG�YچO\�I��P�2\�}àD2gy�>���k�+5�/~4r淈��S鰟�����X��[��=V�~�(MSu;C5�T����*����ٟj!aøg���s��}]���%JV��v�t�<K^o�X��3wuG�i�Xˠ���j� �Ή����=M���:����V��4�Y)fTHD��W�^Z��@�]׺T���o�B!?B�Z�O��8��x�
��th��+�O�����D�ɜ�|*g�=�g��hn���р�!�	�on?&�������Q�ò�6��w,��L�3��܊j�rN��b�q	�7�$SJ�e,��n�l�9�v�ۼqa���-�͡Gl���{�G�Z`/��vF.�%Jӏ��V�*�j݂���	��bמ�o�
U��+�#�{ B��z�{�����k"|��NBf���4��*YJk��:l�F�ε)A��(k �B�͚WA��|�2?E8֣��ZLe�+� �/	&�qI�5ː���o���F�n/8�]7�`�@� �s/��q��K�M�aH0��E��a��:��$ǌю�������9���V�YH(`�!�š�=�\Ra��J(=��s�.5ǍF^�&SH�]up���N�we��s;q��u�ϑ�� ?�.�8��b�Rb�#q�|{Ȋ�i��ϻl����l��LEo���0Q�,o)�u��0�`V��2���BܠF96�#Q��n1�CY��N>n�.:��`�:Rx���DB�*="~�k��2�t̢%�I�,��bg��H���D�Ȕ/�?��n�8�l�{����쑕� 
Vv?�a�!�ڮL�~H��ɉ�a�1���]�+gR�`��Z����հ�Xs2FF��Cs^�u<�����N��	6���k$AaQ��h<�s�����w�DB����Y�ܞ�W�hm�L��� �'	J՚�FB=)�߅�y�Q�/ߖF?���؉��S&\�W:Ʊ��zd��*���Q��%��{�� �5u*T_�O{����ɼ��R�uQ���>�LZ��&Ÿ}�����J����	���ܕ��`!ҟn��ճ--�"�� (�5��p����O��)4�'��f�ky����4w2%.w"�"Ia�-H�Ѷ@� @��H�v��KP�	��"�r#�����\�8���@�"�L�� O�����M�����1�Q� �+���B�X~�ػi�4/TN��^$����^���B}"$uk��oHR�1��l5-B���y����B����]�����::�V�`p~��C�������C7p���>A�w�q�}�c�)�j"�d7.��B��Xx��AS38c@O
v��ҩv�F�mEc ~}��}�
�S�P?N���=GvZag��(�D	>�L��S@Y<���/E��������m ��m��]�6��U-�nd�|�}��Jb�;�2����^�d�+G�)�����ʽ�/�G/t��1��r|̑���P<ؖ��5db���3���?7�� _G�]j�\P���J�Ш��+I���^2�ȳV�]��M����c�����۞���wk�r~QI�P�J��Чf_G~c�� :]�{F�-��Po�e��M�!��$���;$h����E�|h��Du�QRG&|�1�t첗,!5�<�C�@�:�����/X]Rt��߫-mL�<f��:�@Z�,2��3���U\�.׼���9xܕ�|�*�z1t}��#�R�wI��"�N0�,ע�㾗c���v�eb�˦��QMr�s���K��|4jԝd[���i����f�ƂL:��	B���l��75#E�e_��7��{}1g0Tz����F��3�PW����r�ɱ9�Ai�3�q)��� �I���]�Ғm��~J�����^�e8j��N�L-K��{2tn�����9�[ tv�ٽ%\z��\{jg7Y�č��S�JW�r��q��SN*�e��ĳ�A#��0��T��r�ʴ~Fd� �H�b2��hL͋;A{ɧ�B�9��c��^�o$!i���^y�ŜT$����U\���c%=g�W���ݓ$�ۄ�!���/V__0�k��d�aPH@��e�X;�*)|��~d����P����+F�L@i5�[R�V�T4l�΀W�	�|��x�����`����K-β�lq�7Lh�Y��%�Eذ���fǽh8	�� �#��uh��nx{�wS�� ��5�wN�ch�pi�K"��e�N�#&�'X�HU��ٷ�eā���,����y�$�@G7��8��Jk�s��e�3��3%�	#2\
����f�_�����^uG�bn�H�SSI�â�Α�l"j��i��%�F�^g\19��أ��NQ�Ϧ���}�=�T��M�Z�u ������;�:dy��ٯ�~Ye;��D|>�耖����B�5r�&[s�m�ɪ�M��Ej���m�"�$�Lb����:��5�5$����xpXF��P��΃ՈRv�Y�rړ�pI_�y�1K V�\JZYv��J������%�b6��W�� �J�pڷ�z�¯�?s��XpEx3D�D#�ǸK�0aX<�ny�̷���о�9�a���~��pK���5�����8�vį�ۜ�~L��5A���D� �Pd+�����3TBL3��0���A�ѧ�Vp�,��h0|���5"��[��i�Pݠ�+�9�8�J�J4�b{�]}�5�]s7��[����?��J=[اE>h�^^���;LT����v5��7 ���Mƚ��
H���^���@�,�wR����c\�|'�%h{�� ՌѾF��u6 ��&�ڢJ�!ȼ*#k�3(T��F7a(Q��_<��'��R�HJ].����t�*�S����j%��Rp��7�j�_l|tj+��VӢ��uc�QCP^íL��*�N�����o(߷����r:'0%;���O�b��b�����>���TXr<�ψ�cc��
���=�3�yq!jr��毈�,+���Ӕ�y���oȃ�r�ȉ)l�x-�sY���1�/��u�ޞ��e��$p��C:��5ρ���O/"�_f��]7
��p���g���\�\&2:����@���Z�l��G�&�]p����@�b��A��<fR�B�(�y�]�}�[��T�Dtt-�#���t�:�9!��ٶA�>9�x�Ch��h3��";%��e|>-LEs�s �l��M"z�h����#�D�.Ը���?e���"a��Y��]퇡�T�� �`�ʺ�[��]���Z`9B�*x�T0;�(�1��~v��g"G�}�1�QU���%����3�$x�*�?�W�Y	�����l��$��B��o�2�G�y��'Q,�k��!-'iOjHCbk���'�T���`�j�������dw���a|oE���
���a�{5`4�����h.�|r��ѫ�F��	�WIJ��g͗�]к�]ob�C���\w�z�dl�vZ?��%J��V%��ʩ�
�x�>DY��;9���/Ҵu��z,�~u!������\�k��n���ቘ���1��-���Gһ��z��j�O39v8�4�;}����@���\~�e��S
�=~��GrK����/ |���b��7�D����P�����dR��a_$�n`�;G�)E�4�Ml�ʠ��Qoʋ<\<�VD��d�~2�&/f��IV�}#'Q��;E���w���2��ݿ���sz���r�j2b�Ӵ|�#�ep�\�6�e:J�,!T�clg�Oπ&y^7�P��h3?(=�Xd�?�
+�h�R��,�3�Zw=�-���g��
��n����@�Լ~�A���21"7�p0�����`����<�h�ʅ��1W����z�̩�����{��N�����I�������!��f���M�U�L��E������I��)ȥx���X*���X��B�	�gƯ�p��%k��zo�g[�Jr�'���3qƇ�Pv[���c�Vn���-�5���2Ν���(��۬�����~)�(3��n*aι�������'�R�y�W�~��e�L$e%��ye�P�ױ�<��� �ii`K=�N���K�M����y������6�d@���c}]ܫ���$mlV��
L����LOuU��+B0w��(%h���y?�U���r��L
"�^��#+� 5� ^CĖ1���x3T�nP�/=���=�"C�T�u+�^��z@��ra�^#%���Il���Y(�u�a��`����'�R��8qX�x������SQէ#}=��*���b�/�����fC�ZOI|��(J�G_�i�����E�I������)?�r%�=�]M�p�F:~_K1�ecw/^B���/��m����ⴋ����~i7 �q�i���L��o�hҮ�CM�����2�������E��^Unt��l]Ñ�2Қ�	]~)�خ�z�~���B[T%�>=��X�ԮԆ�&��\�����O�%�yߺ׳�]� �<��o�C+���]vJ�v�)>���{A]/��.� ����`*����7�N���藳/̿]��P�(��g��;O��פf"j�Hc:�(��7X4��-��vq�%gho	�,�)�"Q	�.��0�9���9�B�-�lv����6�e���{��C���sY|��*�I��n���ih���/3|�[^���K�ӈ�N� ��T�4��Q|�J5�
�-*'�W�@������{���Q'jX��?�Zl��ݹ�[k�JD�,�0'c�	����[\֥-b��o��m� Wv^���QZP4/>&(���\	�P�_�,��x�>_&|'���.ܭo1�.������3�o���|w{�r@h�*��MV3֘��+��i�k_�f���6�VT):)���M�on�%�a^�{�Gٗ���,�0�����8T©��mQ����3.53�� ���3m�~��$r `�=�݇h�Fg�!�4���W�I���=b7vo�_��rAt")����.�,�_�{�jRZ~��3��2��"�m��y�pd�@�M��<��� �M�E�+D6Pe�P�%���H/�jN����	����02JҰ�����<�9"�}�����Xd�W������	�ik�^h�n��2.�S��Ь�(�e����.9��{P�ˢ1�H�ʌm�;�©����p�x����+d<쯷K�]u�S6��j����^���	����Z����E}�����V�m��	�P?f��<D���y��)��$���
�Y�2S��%M�{�KХ�qO�*窢��YaQse�TT������]ק	��)8e��kf䘷��fc-h3Gz���ư�Ǘ9G�\1�W����e��O]!S�s5�[o�l���%dM��럻ZbD�9&�
E��<����@�Ot[a���OQx�(&:��zp�`��/���	L;�r7@�� 8�{��k�?�>��H�S}t�zD</�vy��'��=�P���ӿ��G��{�����M��Sm���y%
Mj(OI�b�l�P�a�"H��P�lJ?5�K�`�)} Ә�o����&
��b��{��U@3�	Y��V�<�m64x^��^�hZ��N�K@�˪���nG?  �uPZb�.풣/��Juk/ǚI<f�z"㚎��B_�u�}D&C����cwy�L�*�Q=����� Ȉ"�j�e�)l`�>���z����& {F��Jq������,�|�=��Јz��tǴ:w�>�Fw��-= tm$9�C�q�������_֐������|ЀSe��W���}�2��ޡ	q��x�L<<U��mh��1"������ �j��`U���-���v������p.�Ƭ0���,2����)����Rtir��1:.ϒqVD���)�� ��=�Y��~�~��D��i����dt�d��R��Ͳ��3U7��|w�"v<k��UI׈��v��ʭ�����FA[�x'UN4��=�D��@IeI4J��� ?\&l\Nm�해k������Qx]��h����l)+&������|��q�ް&�g�?���_+&�f������b�v>�Z�76��M��C;Ubhç�z��w��D:1�RM����G����(��B�Ƶ���$%�%m�C*
W��1�]>9����2��ϙu��������So$'�F�@B9�E��^�M<q�93U���P��s�:��L�Gg�cq+��k�(N'I�td��[Ft�E�� ��/m�����XW�������u�B�����?��x�FLd9�e 8�ȝ�����,�fO��b^,��O���<ޙ��8y���ƅc�A$�X��<㫁R2��`����4�b���8���Ah��ߦ��!��!2�u\'n�G護��wg��]��Q��;4�sz�ű�-�A���t��u�He����l��
�A��pY�����$_
�����yM�x<�uT����4v�MCJN��X*��	����1���<Q*7�4���ם69��>߬J�E�
C\6�G�G��#b}���[7n�(�d������Um3�CwL�-h�5(���gF�-6��%�_1p�r���Ѽ����61��ֆ��g��w���B��?y@��X�e���Q��ۿ"KZ
;�":̅.���X�U0ʕ���lǔ�/���B4�z�����Ly�O�����~�J	{ ��^;ш�)ϱ�}^���m�E:f���eV��aflk[K�f���t|i}�
&�t�R�����1�c�*{!rP6��,X�^�k>���~8ZW�.�m��  �	$S����sć�Sp��N^�PK}����A�Z��!9��E�:q��Uj�$>A��}p�P=�Ǧ�O�h�d��͂oŞhk�`}+ļ�,�%ǝD=�g�3m�����,n5�)�*�o++�	]�ǵ���	�V�pc �ݹ����>5.l����� �]0�37c��jCET^-O����}������F�h�p��ޡ��ˮ}���\N� &���m<��0&�S�k����8��e&փꠉ��H��p3���%*�<_�L��6����m��d�.<��9����ULp��t��C��63��s��F���s�O�y�xE� Ձ���7R��N�V�{$N�+��^�n�^�l�:���E�Jr�Yg�U!x)�(qTP�U�F۞^�.�n�K�ʃ�����B<��ȿ/�$��[�QT]/a��9;WGg��	P�s�� �)58ն�ߓ���WcP����cq�
�	a�Dn�j�����i�w
��W�"Ӆv>��cG����:D��A��툃f�}�F�`�s�xp���P��S����O��~e ���\kyB�_H�.�!��z���_.��y?1����ŷ��a�j�ܼ�$�m��X=�Q3\!��K1��O�x ��Mot��8u�OpR��8뚾F�s �H���>���}.{�|��pz�(<�_k�E���tάo��x揯�xe��uɢ�Ga"�ȱ ��j�];m��(�A�B�	@׏������9������˲+�x��@n��������B���刔(���{6��Aa�[�h�>k��I�G�0��<T��]�a������VW�Ƨe��]��k��p���h_�ǘ+-�0����OΔ6ۋ=���tG��}�$��Yt�I��iQ��K�ep}��貶�Q�r�	O�G�z��#�[��n�?�������j�Uh����K	T�Ț�SK�#;ܺ7��#D]=��v���|Q��	��\�}�}Ch�U��"�i�L��{��x�dF�dli���t�.�B�JP�6{�|�1I�	< � ��X�J��B?~`��n{�v��[͓��Y�cl�3�]/������9�� ����ƒ���O�n���.�b&�����nJ��7�O�MY����3�s����>L�%�E�A~����}R�6�����,�Ɗ*��~Åv�����nzE�Qs�P"e[ek���v�z���of�{
��6�A1Y��2,%B�~ު8����G���w�Z��qb{z}-5������O��f�I\<�a'H�.Kl8�)�~�Z4�\�Ё�d!��SJ��Tuw�cJ��j8�yfh'n�#�=�eS3��_�����e�\��)�n��Ӊ���H�2"%�O���5K�%-F��f� Ԇ��M�I�2������W�v�sHƐ
�QZ�#>��DK�S�!���P[�h�϶q,��=����š_���]�Ip��V�P���v.�[B�vvY���9��$����3�դ��Ie�4p���A��A�df����Y�ѵ����P�gjD[09�&���a5r��|�+��	W�9{b'G�W�j}�ؗ�2��<�^�$�����$γ����x0<��i牪� 2�~��3�͡1�6@�k0��p�2����"�SEm̝�(@��6�����Շ1��y�
*}
��lN�����;�Y�
-@Ȩ��\5%O����^"!�x��O���Y�����rU�.]E�v��_��Bg,O��B��P�=�5�>���&˘�7Z)�B����g�R��R<��D�b�>f׮��U6m�\`�K^�+��U��[����np��vAYU�0UӬ�r
�b�M�bc%�/���s��pL�5T�5=�' ���7�"���%m�q&˗L�rk�J��"	�oW�芛r�r?R����m�f>N�����`w�z����<�&�'�ٱ��8�]�@-T&g~�����NWJ���%4��-W](�S��t`B�Q ��t�A���8/�M#("n��bj)���"=���#�kXV��c��p�=���c�Q��:p"ي���Ox�84؇�[5��F�l-(��`%�~�����
��#˨-�����w~HA'G[A���%�`V٥k��|�m��Ep�<XH�(�Yr�Z1k516�V�>TFΰ�xh�}�aWHZk�\��G��R>���r�*�" 9�>6x�k�����d�4Dѕ܈N�����|�]�ZhT�ߏ>@Q�c���6S���#;3d���pBEGU���TN�ecR�,WFv���<�vj���>]���[R"��x�����'o��(�^aA*�&L'�8�x1yj.�pKv
,���9�Q�ĉFK,%׹�:9�fZ��o��km@��8�Ԉ��2���_J6O~;|HO��a$>Yk#h0������-��&t����@��?�V<�Χ�_йn���������M�R�^�z޳ZC���и_NH���|�Ğk?����u$�Jj	lZ�����a<�(U#��Ϛi0����p�������ǌ'{�'oG��=�mr X�8q����/'xze}$��4�������&�~Z��E�@H�뎚.f��R5�3(T��6�o2A�K�>�,��k9a�!%y�=����ns�u��}<�����R��S$���
�4p��"r��ʞ�Þ�k低��{��*��QV�D� hI�-�	�*)������H�M��P��l-�l�p�8���ZnW0�\��oӇ���H_rhe�B�������j�[A�A�2\Bs	:����Ï�?]`ڸ=�@-�8z��U�@�:��Z̞�j���^�"�I(Z���%��4���~�"���o�|kL��B�����䆐`6����4�=�m�/�D��@��(�E�"�Hc��<��z��S1�ݸ�����8�(n2�FU.��XU�E	�Q�uė򢺐6>���j���؏s�� �}.�Յ��iN�z��H��/��-���0�G:��Қ����� ��Iϊ���Ԍ���Q��x�r��b�d�h�#j��T1��c��Æ���~���m�I�X����~�>|p��K�d��H�[)����6�K�d׾ϕ�|�@�M�~4ϡ�qF�����z�@	�d�t\�+e\&2
���Y�?T�U'[��J2�̻�fve[� �F��:�aۺ�VX�-�7m@�#"9�T0��/�:=����/[w5;��OI�41�s��F�� 2�u���K3ДI�HZ����vF;��D{gy��xM}�B�R�Y��,Ss�H!|�����dK�� s(�肓��HHc���y`o�K�Ţ(k��OiT�s\��CkEG�/ظ���6Ia����-�$�N���@y���HH][��d[��Jȓ�Mc�o��ςx�����B���1�u�4���޵��Qe \�E6�Ďʵd����j8_�f&/ŀ3?1����`�{1���@>��L�����SH��-�%��}���c�Q-QL�7[`�:V�_L��(��U֬g�"��P�a����3�g�L�-ۃ��	�X;�dJ �Mg�����B�Zǵ�$��ǭ����Ze�{`�j��� ��� ��rM�jH&j��L�U,ۋ�m8����I[x��x鯓Vg�
��&r��]�[��V�`ZS��S��^̦A����1�,��x't�臞��uV��)S+���Y R��	���Mh?W�R=��6�e!��@׊�Q괚qN��@�!bq��p�O&f�r�5���`�dт�גs�5V8�O�Ja�7�u�V5G�iN	��'�-�
��42\���@���	���r����q}��r�}��]C� k��qݱ0.q	��D*��T�d�Ej�p�����ӊⲐE1���=���2�� �)��,�|S�Q���N��3�ߞ��iD���o�T=�`+u����� <N
�j��H���C���4�9o�������!D�̗�-T��E��p��=��b�"�D���0�[��0sr�3�K��ぶ%��5!����VՄ]�3� ����q�"�N>�&�����w#O֛�k	�x}|�|�oR	�P�Á2����n����	93��������[C�.m��je���ϴ�ϴ,�[G)��3��h�`�Q��{=Ӊ��(��Z����B$�#��ٯ�e��OU��foǄWS�1�n���K� � ��#��Fi��|�r�n�6��vT���c;�6܄!- r2A��گ�ՂR�Zo4;�[���g�����O��,��������n�����۟w�(���s���K���ԓ��5�wA!��4��R%K�+`k�1!Tr3��I[�n�1	�*"�yS��_���MV�b��}�m1�7ϒ4W�#ޠX��Q���y���+�m��d�
��D9^jR0̋��+n�.���+����N\ad��u��b�����L�j8�Ⱦ!IO b�#��\"����Ѵ�["�0�i��!��gcUB��U��9���[i
�o���ZR�R��T���?ۇ�rGB3��W�/���	��"[�n�����}/��c��G��I��
1��{�B>�8����0C��02tԑ���9fe�hea����-������X�=���Kèn����MC���8��)a-�KW� n�
�����I/ ��Ss>�����x[�����+��?J ��(+]�@�R'�������C��D�7�Х�uA�� pͱ�����Ҍ
��,�E�ʟZEMy�@!�gAe��1���ܝ!CH\�h>��IE�J�#�^�ľ�i�`�hz=MVQ�@i�Ă��ӕ�
��<�K�-Ĥ%f�7N)��]�г+x�֪��Y9� ~;�P�i���b��,�,U3�0�8/�#��	Z�Z���r�F��)`�J��̶u��U'�᫭�S�HE]���@��z������s1��
�82���Na�a�������w'}6`�" �CMF����G5gH�ZuN�?l�3�C�Wim-�5�T���ɋf-�^�7O����FQ��@q[���A��A�ȁ��4�i��^����.�A��t=�yPw�[�J��<�Ն�o����V� &��x��\X�k�J�~t�L?���+nt�P#�-�+��������L���q��i��@���l`�`0�q:�0>t����/�	���k7�-�<��x�vW;1�	�d��ۉ=}����O�I�VEwQ��+�RS��(_��]�~j��Q�����h;����.W�~��ї�]W[�*��`[�msSF$E-�hj��]y4L������b%M�tZ�D?؝�i��V�׳o���OגE0�%�8-`��A�$V���J�L�v b�{�j��%���)����������w���a��Su#�mÊ����s��J�"�h֍J���7󕃼�{(���L��A0�t����-�;�5W����;�R�g)��4<��q�0�L`D钉Q0�y\�PO���71�qǱ��/�E{oI��^H$1���3��=t��!��ZJF7��/ ug免�B��Um��!Df�ǌ�I҅x�[5��i(����=�$��p��֐��j�`�kmŉ�ae  e�θ��
��b�I!}$5(���$�1,̔鿧�U�6��U�i:զ��C7u�o��d���xM{Ա��g}���j�+H-z?��d�Mb���#)q�7kP���x����1z�Mp�P(�}-� �a�]��唠ԏ����V2�@G�_�aR�*�\�hx�Պ�7+n1�q0O�X)��u}��#_۹R���ϥ�,�g�v=V����jl+�[cr&3L ��My�.eh?�y�b�''�|G[<a.��k"�A��Y�B�����YRp�,XIZ_M�Ou;�:fX�	 &���6��]�~��oŠ�PG.儬������ٴ�6ZWЂ�a"d����=S�r���!���Fv��_#����۽Z�u���6b=�y�l �E
bBy	�ܔ��@����p�ώ�&d��J��Q�	�oM~3S�N+���i��x�K�>yq*��������ͽJ۸8����bZHo<�� ���^�]�&�p/<��2O��ο��kq�-���|���b6Q�z�����Iٔ�����Y #�0����2�(�:�#X8*�wǂ���*��X��g�\=6<2r���%k�����^T��$��a����� �B�:}j>����V4����},�4���P�ISP�x���p����Hl7z��uQLdn��v�����*�z��P�&�p/5��|6���5��p�;�	�T����6��g���J��Cd�2�T>�.*��N(�A'��He {��"ۊ�b�϶	h{K4��]���γf�u��"!{w�k6��m^���I�Yl8��ǋ�/ൌa;��3x(����eEj����@fzH�:��ѡ�L��mh8��|� ��1�Ap�%�t�eƂ��r��Sm�O�VP�w�{���TLi�}�E��A�$7ܽ�qs���5Vb0v��l5m�l��.N�	G�8Ny����� Jz1�`�O/a��u@Sd>�g� ^[�9�wf�[��f���"	�He�*xRs��{U�;R#��|�����5vN�a'����8E����im��c�ju#�o�?�C�P,�������j���N_��x衁��܎@�BA��+�$�A�����ۍW�_���d@Pr�ty�:wbāV����M�)ڹ08b���vjgݾ�=�'��E��7=�gX��Xͨ��(7��x_pƙ4�b3[�
֗�<���Vc��3����kK��7��[r0��7�� 6��=5���u�%؊�B�zL�F�̄�Y����ɘ�D�]��2������7�&�O/B�J����]��c]Dc�2�LT�;+���f� 0&{r�"}9[!�U�=��:�������I��ޡ`��<�&�6Lr��^�s�<���I<�|���^��@�~���.����y ^����Y���R��T��=��Qp�n!&[��5��9C�u�"S��"r���p��i�Z�bkt���DgR�0�%|H�@h󰣠*]&�i��@�f��8�*i�E7'�,'��}	��pn|�Jr���Ӓ��@��#8�NIW�.�e]R�����b-�l���;#G��7�,�G�)���;=1q�欟�����Fs�4c�>ˣno �`��rd��.<p�H�5~����埈�Ό���@K&���[�����̈N���3ASɉ6R�6���Lr ��� �{��˜�r��O�_��uV"����3����kO������n�wJ"E���<c�c��J2�9h y�"�$P؃,���_�T����?�%%8n�)�.Vפ�hFy�4|���J�h���9�H'���?��B���ӢӜQk�e���jQ�u�~"�o���<n�)�
��l��͂Ű8�٭j+K�e�:�m�� �	1vT�5_��d5�2?=I� ��g;��-���pޏ��82���p�}���+����5z��5+�����e�G<ZE��_=	hc��M$���Z��H=uS�,0�=�β��	a>O~0�H��?�:O�"�] �T�(�[TcV�o���0����7��ԐH���S\�&x{Z�qc:��d�,���Ɠ�J�5C�É�q~0h̀=��4's�h�||^�~���~�����7�}��-��7�$�Y�u�# &bS-�m����Q�V[dEZ��<
�k�=u� ��w^�@�j�~pY����,Xt]q�V,�RqA����u��1X����m�8�!�1L��C�` E{��A-�*/�RWdDܺ�良��yp{j41��P�{PI�n^���縦.�wv���`�`�̱�{��ї:�K�k"���;T�?"�DL�G,�e���ݜd��P����lX�)��m��_.X�`=��Sd�:���������y��J�_���`�P���(Ho}�	P6M�N���Mt�>�7x~�Q��os�V����+-�_7JC�}��ɀ'D��� ?�KI��o�Җ*_��͸�$��Z9p�M	R�B�jge��Zت_�Ui<߻pM���MK������S��9L�}n8|\�c�#U���G�Tc�}�f�b<��o���W���Np�	�6�1���6���L��t�(ۉk�Zrڴ��ȶ"��Ǟ�v��o�\y���09�F8������HOA�]��la�r�^�bHMg5�% d'�������GZ��;�h��=���"K*T�!����X��'g�$V��<�q�I����_�٘�\�C��a�$��n$��ş��IE&]�����@������
a�C�Pe�ͼ�i���� �~�*�m�x�U�]ݩ?}ί�h%[�7]��@}���υ��nc�|y[����ж#�'�1]'D�*�S�4Z�~�J:78��ο��DX���8�R�5b;��[��D��;o��z袅�+�+�Ԗ��3i:A>{�^7��p����8t\��OH��Ŧ~��s���=h�Q��LV����-;F��ή��Z6i�K��¼���<xC /Ř���x}�p��"蠑ز�WH�w�v��;��̺�d�7!��2�g���A@0�H�g�(@��R�	ǌ~�:�O!���`F�~�4(ohW�S�(�����%��d�j�m�C&s��?Gc��+8�X�A�����$��xlY�[	 )!�@Ҳ:�[;kX�����n�3wÇ��D$�E��%&Y�z�6ypK�ꠑ, dʁ�J�=�H]���ޑ���n׏"�\�X�vS��p�J�9�۶�7������f�|0g��+m��O��=�3G�G�0-����B�HEf	'�N]�Ю�	-���'xg�E��SjR6�m��%=N�c ���5��r����o�X�s��w�z��.F��H���b��K��Vv� �11�:�(~p7[T����b&������W���*���MU#�@}������
+;��"��huY�M5Y��[3<��hڸrA����*
��l���I��w���-���� W$�I����(��� ���|����v��)�>=_�vy,����X�%]�&:��%�NQs��Rm��B�h��)�p�qi�z(~��:a>��2i�~�>]�iq�Q}|���'��銏� �
(c�]RZ�3�����j���������֔"����/C�;�!SLĈ'�!_�۬tҷ3^I>�m9|�2	��1� $! 
����#�����x[�)�قN�v����w��~y��	5�S�cL�F}ִ�H�́��%Q)>�����- �J<���#�M�F���2���Cʆ�I��#`�7D�5:����^Z �}c������H�0^�ۅy�z8{�>��j�����amՆ9���O{�l�b5����n8#3���S���L��Z��|��Z�9�"D��T��~�Kx�(�����6Q�Y�ʶ�3�m5 ��w�4':�2���hl��&�	>���,Pl�n 4�dc�����" �>f.��.�_�-?�_'
d#X��&���s�i���?R�f./� @f�����O��%��BҲ�aj���~���Pˤ�C�Y��؆�-�E��:�&t��a	��~�&2&��~6�B���iϼ�Z�+�Ky]o�R��i1q������j��;�a58��y�d��k���A�kZ���;W���l4�lsn�"R�B&��!Pa�GQ[G�ڥ��<�c*wA�S�V���f��7�p�G���BA"ڟ���������40�Z?O`�b�w�##�h��2�/������dƼ���hi�w��F�o����ސ _�3��N���yP��s�a�wdPt�G��L��p��C����_���_?�q%v�';R�B��]x.���_ݡ�6�X��&��K6���%-˾/�>h	΢����p�j����7��yy��$���Adk���`\dm�&���vNLk�V���2���ÐkbX���M��]�nbvH��.\�e���q^�c.:@���ƏGL�Q :�01�w��m���o}K�*�U�r� *��P h���� 3A� 0|&�x���H{D"}�
>R'�ITr~�|�D%#K�S�� ��؅nx��)E�Ρ��O��߁+���(tǮ!jS���ŉ���D�Zv_�!O������<��QI�]�E���-vj�7�q�ۉd�6���ʄ.f�J��f����O��͞�K��u1˴��~j.�?�c�x?��DF�B#ㄻ9�<��,0;���_�b.���\�d���Yd�B�� ���Xɢ�`if�e%���-w���I�����U#ǠG�Y	>Ԯ6c~ɍ{U���Sg��i�V����3k�U��6�C�is	aX1�ݔ��ȚYR�ٚ޽�wF�P��ܨ}��!�$�e+iwl��3�>H�"�8S��W��7J=�`�w��� ���/%P�I�5�c��.��{	�[*�����}�B�*�N�zX��q�UL?6�(���Ѧ�yp�p�Ĥ����>�T�sTDB	;~i0�����ra"�h.�)Z(��q1��
���qp}�9�l|}I�A6[渉;����Y(����)&��+H �OU�#H�o�/��`�R�H�U%��1}�SZ�nC+��!UG{i����
Fď���_��q�i+Ql鍸��)������PI�=fw��G'��m,����Tfn`nyWit��c�cz�?�� �-JZ}7e�8mڰA �f���h{����՘��7y1��Q�����'݊\���A2,WZ:P�Q�Ͱ6�E�Э�GIE��Q��}pms������`P�E4��vW�H��RF�v���sމ�I�sY��Y��٬�1��	�Yۛ�+�)�yĊ���ݑ�f��|���v�$ڗ	vW��b�L^˅lԵ������W��99׃d�O}~)�'Q⚹��c�7�3^P�ʘ�#��oV��r@�<B�;F��ؑK�������(�G
�Z׾��s��1®����W�k������^y/u��TL�򢖸�[t���*�ϸ+�] %md�~�˫=��-�+�˵�����Kg�x��!���	�b}��r�\,�~�P3-���P��$����C�lI�_)���bT��3������~b��&��֢mg	���y=.�ˣHW9~��M�[6�9��4���U<�a_�պ8.�f<سq��!E�*ʍ+��^b�Oq��y���dn=��͢�`�tE9M�⤀?�_�j��OR		�q����߉F)�<�y��2��W�-��t^@ ��T���a=�xr͹�R��od:���+N���2ֈk<դ񽾮-f:�*[�p�r�,��Q�@r��o���v�\'�mct��#�W6�y��&��q-G؞;F�|- �7��"�$��r�޷�z"�K�z[�Q�l5��(�񨁌�h*i��b�����?쀵}�!�����
�P�;��r��I�\;q=s��O����D���~E��s�|,��5���8�"�X	��@t����'���!���� \��1$����1���V�ٽL�4�D�;B 6�d��=�'�B��g��+�h��dv���l��T�ϔ�b��ʿ�2�
�/�t���|��j�9��}iʱ����.~R�~��7[Ip�s�8�$:�#W]�NK�;����P_��1��F	�o���+O�t�+�^��̖˺<������/[�t���������S_n#!�i!Fk�?��"#�5zKDM��IZ��}3ҴC�a~�[�ZPg�G�=�����ڷ\0�j;�����]�ܡ!u���%���|�Z:q�*UId���E<�F����+a&Y����5Q��י����	\�&@*#�:��*�j!�מ�Ql������l�žEZQ����l����Flw=�t��4v���Q%�����r���C.�a�=�`S��T�H�;��f�b���@�j�lE���Mf+���|�L�v�7�0$����P��|�D�>ԙ��3�JX�鏄�G֩Ԗ��V�R�?��5�TD~�hH�*e^��O^�x�t�������G@JW#��w�!��������L�{U-�
)sk���)�(M���mMt���U{C|�����A� )�p����F�%&N$��Ʃ"їW��tCU��w�YڦB�?�����f\��4���?�&ֻ	r���Hí�5x]�b��&���Ϙ��Z`U�]h���.���K.���̑l1�\�h�?���ⅽ1���Z��Қ�L���C^}��4��2�<�n���}�_1�Pӏ2�_"����&��VSN�g���`���WW��';ܯ=P��1%}�����1$bb.k�+?�����n�SO{!Ӡ��ת�<I*B��m�*נ|���A�6�\�A]��?��������G����+��<q �%�UD$
VFl����W��r����R���Ex�*����c���#~�c��Ɍ5��-�Q��o�jɔ�F�GˁaUfK�N"����}�/[]��4ں� ��G�!`��C���ǉ?|�i�O}�?P�Ճ�l�R�'�-���x�C��E������`��sK���~���B�B'����iP �p�pU�"�2 q�f^��7����>��mw�H�>C����?�r�v�g�$�f3�H�^��Ҧ�@2�T0����@��oY[%���5�P��G�4�����	@d�#%eѮ�SiG�ܿ���Ժ�1�y�h�f,�mg2#a���T�A������n��7��b�o�%JP�k�bj�Y��r
*w�Ou6��+Z������TH��@3	�(�1.�9y^����<�"�v�g�<�
k�x4D�
5��D��lG�:�F��k���ܵ�x$*r�>tl�+�̋m�b��Z-h� F>&��i��N�I����+��㠃p�]G2�dzm2���-�Pܘ��GB5��x�rw��D#?��M�v���i�H<C7�̨����lC/�GJy������bO",bÕ��t����J;�#ڏ ��v�!ۧ,�-x�j��kb8gA�ee#������ >� `:O��N�3�]ݝ_5r���53�2
7��F|��=k��j��P��� ����n0� ��-&�[�Щ�y.:/��7�q|hZ����7ks�P*���z2(�X��_L�e�m̍5E�����{*�	�LԚ��J*Oy�p �:�"2p��D`гPW!�{z�Z���`���9�� $}��먶�l��X��E(���Ⱦz�&P�0jֲx.�>b���Qf��δ*�U����L_oa��Ml_���_�Υ�q:���_Q�}*���Aױ�S���A��B� d0��0a���h�RI����B|g�,@���X~,���=5I2��u4�%Y�e:k���իc��}��K� �H2Vb@B3�k�H�������3a�ṓ�ȘUp�9����h�� CyW&��^�r`��s���h/�� �>��&�8�U�֎+s�.?_#�~�{X$Jg�J����F�Y��=mfh#�*�˶�/��f�o"�E�J�
z��p W���ҟi�.־��'�3��tb��W�K�"��Ѩ&*~w�*��@J�������WB��G�X����ӷ��Kx�p��.�|���O�B� &D��F�;Ͱ�� ���&��=�oX3��g��9^Wb�3;h�
�]��I=���=���v����kma�����a�2��ٽ+��Q�舟�A��i S�pC���ɘ�vh{�@>��
{�%�$�W�*��wH`^3mj��Q\ �7�lʻ�SS`��(�MV<������u��Qd�|k�$@����LZ=��s�{eN �d���M���ж	�EE=�Gl��;j�MD�^.uv,��$�HX��=�o�-2x\�*��� ����i�[�2{j��C�U�!݊
���n2{��Ґ�6�.7�뒤>fQ%�M�8���1v��aO��̻�Ĕ߽&��R*��fzsW����6�ʳ��ӵ�pA�q2�	S� �ڊ%v��,Τ3�����5B��	I�B��^uG��5��\!h�9���T�gFm͝9i�L�|�O���Gm~Lуn �1��X��G��$�p�Y#N�RW�+KB����Ut�}�s���V�黜|�f�d��`}�''�(���5Ly6%-�&-|1g����{҆����:_�$ n��U�%�`h�,~k� �"o�zy����%"�f7T5Ed�c2�3�9���%9 xg����;-	q�s�;r��X�yY��9��(�HR�L�q�<xD5���;�� �Dt	�*�mЎ�Sud�\�9-Ԯ�����AP��{I�A"c,�Q��j�g�p��R�J/��ؙ]��7aL+\c�%1����ގ���E�^�S�J�(J*O-�s��9�+o*Y �X�<_���k����5Y�6�����J�M���?L��@�Yu�A�5���*�E%�(X�):�i��c�B��y�ר ��ݬV��Kyܾ��<T3�1���'�G��`��Tph���L�A��~��k���,N`퍤�N���>�M�����9�GrkW���e�04PV�b�m�O�K�m��\�O��	g�թ`���eXo�C�#���0Gƍ��P����07����͙���C�95�ri&a��`��x���Jޡ����r�F����D5E��g�<&���['�T6�:����a_�@�Ű�.�S�a�8^U]�b��bN7L����ͧ7�B-��Q�~ǁ�_=�j�X�l@%5���)�f�IX_W�j��h%�;�5��O�ݙ��3`�+d��9��q�?�?������d\f5��&���*(K�ٶ)�*o�a���ӿĘ��uj�`��1Ґ�W���hߔ���\�	�go�	Gͥ#�g��*z��"I�e�y1V�t@���}/�!W�Ѯ��2�e����̇O�]�mR�����~Iб�
/k���-ۚ�����'��*7��䵺��i�����]4��$AITZ�ҋ�`y$k���e��"��M^��
����"�k�`%���;�Q��V�hX2T�K?��\>��E0iiiMPg$��r�Mfd0'���;RtH6�_�z<���L�Y�N@�Zpn���]�c'P�jDn��,�U���ێ��5�%F��>����k4���M��*p�G������W<V��a��g��zL�T>�]�S��u�S�{��6�ƪN���?4�Q�Eo�>�Ҡt��6�����QD
��Ն̔�Q�G�������[cɯ`�:a�Ψ�J� E1[�>\�i�%Βb�kZ�\����Y�1�z�2:_��ab��|O3L�f��4�P����UT��e����`myS��X�6�v<u�Z������Ć��}ڪ����n�U�����Z��s�%Q%T�|����mއ����DZ��~��TZ�\�oF�C]S̔|ˌ�^ct_{$!N=Q�O�耎���v�D���\/��f��tn>�6�����Z^{��| ���z�(0m%6����Ϟso[M�?�ߝ�n��B�:�T��3��D@XV՟�&$��Se?H��s�H|>�&Z^��G�w�,��$*�[n�G�>�5P��nD''rX�f����%��<�����Agm'V#r��g2p�ʽ�i�x���?M����gW��핍��R�	�be�;o���jN��Qd@��d�^�f��e��ylO���(F9R�
�m	�Ȣ�T�zPb
8�<�x�����ژ�	;A�$��G�?Π?�pb�e�G�n�D&Y��:_�#��4-]�	�ǅ��<�+�E��|���t
eÁ����Ē2�.�pLSl��*^�Tβ����,�U�l1����I�OL^Syz9��j5�n��fą DYg�O�|�O���K/i��c��8��N�!���Z���EQ��듍���/:�x�ndgC���a"�r��#�r�iS���Jz�h�~����0�#��[�����إ��BV��@����/����wCp ��T�A�qrڸ3K%,�6MEw>y���~��$k�����&�DJa����D�g��V�*�[ҡ��P��f�`����8��cz�'�)� >�_Z�U�Lb?��Yf(��[����jub7>*���/cR�n�f��n�6�ks2Jo�����9Y�
��K	����e�ʼi�S �չ:p
�;��u�s͙��lQ�M�u�	`1;l�U'�ob��7��I6�,�޸d	>E�D��:�񅖓Y3�^d�JĔ��`M�q|.�֮��+Z#gv���i̟�g��J��	f����i+� �Q�C�i���ch��+N)0��.��DR!�`�Æ�=�FE9F,i���!���3RP
�F��^�^(T����P���2C����+35����|(n�L֕���V�~fq��T8��P�E�	��Gȓ3,5-�5��t�~0��l�0ڊ�7�Jj��I���yC�/��0˽���}v
V�n$����F�;�t�!����� �OX�Ԩ��P|Va~+`����&�?��"�1��&�Yf�^?��\�4�D��ķ@j}�GN�v����9z�,���A���Id���T��r� ����:4�M[̎V�a���H?��&����s������4K��KB��9�]���Bt[��R��N���S�$4���*�~�B�[p�"[�u"�>�Nce�����Z�,�I�u �ߛc Ƀ�QV%ӿ�R(�y���v��i��G���ޡ�3|��Jw@�$�,�/+@�_�AJ.�xi�DE%Rd��T���K�r��\����4�F��Pm��.��#���4�����-X�7}48��eR�,�g�`g��7)����h:�9&j�_���cfe��g�b��9�x��#�c0��lO����3I���)�+�ݭ���k1�A�ѣ�������|P�~�E����4���9� �������E�e4u���b���K���CA����B�Z�Kz��LA�݅�������p�����Xʺ�=��BqN/�v��l�,wH�4�-N�#�
8Q(��vh[@�Y"����@*c� �����P(MO60ʟ5�h@�j�u'��6Aăx|�(]�Z,���Q�-�����a:�]ω�p3�&2�'���Uf��ݺ���.Y��3���6 U;��Oip�����ou�������!}�DKJ�h��^��S/h�;�|Ny��LL�"�C��U{[���O���nA�F
� �.�\�J�#�"�/�2�?^m��,
�����p���ؓ�'�dpl ����>�l�	��b��"���*�՞B��R�Y���U��)$m�5;	L�)u�*
�T����U�կ�Շ����%0w�W���	d#�T��l������z��\<h�s\�eɫf_�;��8y�>x�ι\̽G����:7�s���i
lq��e����)iƃϒtiM���*��/�۴A�õ�.�$�ª�}��#������#�+��Z�V7��>$$G��4��j�Ȅ���ޤYT�������dj�Avp2'H�.�������I��K
�c��̇��]��2��q.΅�i�N�S�25
@�~KgЋ I�N{�{Dc��o`'\ʢ��.�>#��4����ݱ�N2�������[�F��2Nձ��=vǧ����8�������:��/�el�e�����3pn��=���0�=����9��ё�����Q��D�[�i<�ϸ�9	����������&>sɘ	�τ���	Z������(�PW/��G��s|�*=%��P���fBV�V�[��,C2Rd��u���U��Ȼ��К{P�y�ԏ%P�Ĕ����j ��A�h�0k���3�١��ش�5�p�b��!��&�8�
��#��|3a5'P���u�a6���$��y��)J�!�~� �d��(�Vk����N.BN
�t�9N�q���Tģ�;�E
�N�2�~���
��h?����g�y�~�Qm���	c/>]��e���H�O:p�5ƹ����^��©\Gy(Z�"�����1ᡦ n����ꀋ��X�E�����.m�\_�����}�	�ױ bFk2{��+D� _�c�*h�joe���_�L'Ч�4~�e�����i+��I�?�4����[4��FpeTf"<���X�������<k{�)��#k[�J�G*|ېΫ�Mq�h�\x����,�WdC�L,�dR��曊�/8c�*e|E��r5O7�@�����̓��A���B�8��4;�����m�hW�qC��&�&�5��`�7"����b�j����#"�!�z!�\)�|yj����)ď�x\/n��ml/68��ؚ����Z�;i���R���FX�׸.Ӕ�y��y�JL�N��N�vƣ�a��mЃ𵐘��8t�h9�&?A_�uMX��'��.بw��c��Y	qjJ���X���h�ŵh���<d.�6��g��!'N���ib�QP�O?����K;��NL�n�]2�j�)���7դV̰���[/��qʔ��g�>'��si�==L!��S�%PqIv�O��j����DD�2�̚F_���ܓ���t T��NFO#����騱sؘmFl,u�|Hv����JL����}�x�����e3-�8:�nЋ�|J�ӈ,j�k-�I�1�ľ�㛟Gk<,�١�dڂ;A�z�����,���'�sS,ZgOhZ��$�
������Cq}�]bwu��ˈ]�ğk��TE��ݣ��@D�Q
�H�F�a@��/r)��.Ц��V���6���D�a���G��	����b�)�uծY}�-�t����L&�s���X�@����	l�$�.�WeT]�s��)�'ڍ��Yکt;���b�q���5Bh݀n�ؑ=�|�J�C��i��ZJ��U#@`ef���T!�-%�w��7��^��*��z�b/������^(�ی��������XU���l�"�`#x�A+9���P����< ��2K��N�֠��>��	���v��y�;���i�T�t�j���+6$5Q�]�6��
�)�z��>N�[c~�������6�W�w�8�R���d4�>I�cX6(.�Ɇ��8�Ϣ�sé�ڍ
EB���+�Ђ�Y}��a�]���~�s��=I�v6q�؄�f+�ߐ�e�/0CW��p������m>����|��6�(+��!��t����)����I$GD�ۮ!սY'�z�К����|��'�f��{`��	u;r���HwȾP]��T�v���/�٣�L��&�,����h[9e��-��v��l� O|\� !t �j�g�O�[*;���Ļ"q*e��@��;H+Z�q(P�8��wDD�qB�}F�y��4a��A��8��.f�+)�f�&��ɂc�I���@P�q��બo����|��3|�8��3~LQ4�x7p_�8Z��P?L�G��k��@FU�(�! gI$�N��mާ�o�ȹ�ID�vO�xj���C�9z}'�n��6`ې���!��Ƅ1�P/�LmFL�~��!���l��!4�+|��m�LF���-6u�a�����\�K�ΠuĸR���}s�и��I�F���bmŨɦ����*2T��I��#�	�?+ы@n.)U!vՆ4M��CF�^��5���e��@i��)5qV��|����A<�#�K�x�qq�JC��
���bC��;�7�����(�4߰�*�MkH
w�kp��� ڛ��3[�-^� �o#<��ӷ*�݉�����`;�ebB}	��r�X|�3��'����?����lu�u;|bٕM��߃���l(�h󥳓MB�ΐ�䈆bZ�����@O��/�Y֭V��U��D�E����s<#ж�4.��X���$�ޤ,_M��Dw}��ʨ�����.�<��s?}�bh�/qX	7�Xk��W@U>�"���Ԗn���H ���]wAG}�J�ska�n�"C1�������oю0�
�M-)�zlհk�i�D����̂�0$x�~~BҸn���jnZM2�rj��|2^{LkV:Ur� �S�c	f{vU	�i�0p/ �"����=R�I�D#�Ԥ���|k��J2:�}G�Mt��sDNN�Q�5��Eq0�o*GP��p��\ "6�`��b�v��>reN�#!��t5������仴��[x������	�D?��Z���y�A�[��d��|maW'�-��S���O'���3Y\��k�e�}9i)ƕI�wO�5��Re^SW�9[����·ʒY��hí���:���e�}�V�2�K�M�ÖΌK����Ij�Gn���7Rf�gUP�!�������n9���c5�4��8���sc�� RB!΄z#*�T�5��	�5@0��(�l�S�)�âo��3�H	��	�n��2�Ħ/_P:ꈂ,��x����+�vPo�f��٠oG�m�]-���pnzJ�B��S�bIw��/ 	��4�42��\&{�ݙHAѥZd�v�)\1X��`~�����,�	��F�Dz�{ ��+\�r�z%7 a�M�N<�_�4�]a(�sNa<��@���m_|k��ח��9L��>j������6�a�G������}��@������k]D�]h'�(rҐ+�e}&��%��?R������� 
MB�N���s̥�c�,�S޿^�<	��%���9� Z�"�����i�Ӌg��o�ѯq��ז�j��7�c1��n(��Pk"|-l����R.�~�' k/��yض:Ra$��Idu8��j'F�` �4A�vI��%��C�C|w��``��s���z�*��:rPGb�f�ʄ�k��M^�I��2{�Do��wuS�xyaCA��I�O��(�����V�f�*��1/��Ū��.�=�)s��=�^��%(}�X# ��.o�w.j�K��ew\f"+��z���/=��YGcKY��@�_®й�9A���t�I��~�#�T��B{b�hGJ(�lٷ����j�z7p��������t�\U"[غ�tR���8=c��2�T��.1��zY͞��sn���@���]��Mc'?��W��	��s�>�E_�R���������qܙ��%s/��K.�+����ߦ~ﻑ�=�[�����`��{!Tr��1�$~����t�,��ף��V1�'�oU2��oYXy�9��XN�m���h�&���72~J����E�%N�MRo�̀�(�e3��_�L�)�� �����گ�V���{>zhu@�v`1�&����_E�,N����M¡ �7�v����*ﺰx���a-�����)���,�8��X�u�Zp�e����[�	�a���$�;Er��S�M�M�$�k��7�F���0��R�6d+�%N�ݖR��a�|;(a���$��X�*�¯�q}�w���T��� %�Q_�yT0�G?\�
�w]J��{�2�FNz3��[��sʾ�Ʈܰ�,�hȵ\�3�u)'�+ODs�;��E6��~��>�0�<��[���	Vb�I�/�Il�#0-uU��ƻ��/J����7��>�1,[��Nu��[�S��^�2 vD1=m:��m�ڒeDb�-�5�78H��vޚ�Ai"���h�/Y�,���ν�o� m�>x#HV��6�Y�,X��kp�7f�����`A҉9�#�����������!gV�����Ֆ���*%�zCݘtF�7�+fW�Xy���հ��̝�d�J�I��D�
f�<����p��v�+XK� u�p+5w���&š�hj%���c3No� ���0��)[P�kfw�B&�~��1�J�O&���id��f�p�p] �	������pH��椣f���*��q�-���@x����{`B���M���eN���K	��K�v����Ty����\p�Yj�$�t��Fto���g�U�}�4\�v��ᷢ��,��<���E�h�)TL�w�"���b\S�n݅�LN���M�@��r�de�X��B��;Z`p�ʐ\^��zP�,���V����+��l�RK/�AE�mJ� ��oܦ�b<�|(z�ނ��d�^,�.���MP�V��NKR�͊�SvDaA�ls"�ދp#&>��I��B��5A�4e:@�(Ɖ-��Ż�J�~�(��賥Os�rZɟ��<�.����o]��˸�B?��x�^xZ������5u'A�d����,Rm�\��b4�^0.p���ܧ�.�>I����o�ׯ��3�%�š�Ңl���32}�%�꬘�VPVj��7D,Z>��$i#�L�A�;L�d�۽�	�y�ܘR�b�'z>���h=W
:��!y�I�o�mL�x�$`��ǧ�9ql���9 #D�]k�ǒ=I������M�cm��M3v vU4L?�\슄0�c%�B��ѵZ�%����|�����e%>eB��K���b�@�_�r�C�1�b�����QtR?Q�x_��eb�L�qkNL�me��.������-'�Cp�� s6�����SWz2�O��4��6Q��¦�S�o�Q	(�[��3Á?���|�$ɻsLz����B�nȈ�kZ��:���Ք?�|y2򎈱�Lb&ZE�5�t�ӽY���b��SU�m�=��DZ'�|�ik�K��Q%�^�t2�$Ԇ P��ڃ��r�9>Tz�U�Oln�����2E���YV��chgu�����j9�R����	$Z�{mu�e�W�1��>T#X�c)����<r�K� �Z�������y)>��Ń.nZ����MbMו�&3كW�Sj[�6����W��E��-�"��8�_���W�w�e���bv#\r��!H���
�-�>+-�AG�s�V!�cQ��0�;k@2�{�����a��)�iX�}���)j/ ��:m0! 
�I��A��-�Q7Sl?��W4�y*�͑a�C�@m �C^�$��Nٞ]ϧ�I�d�)U\�(S�M�뛖ߧ^_ȒS�'טo�����fm�/u���	K�2�L P?J�X �ލ�L:���c�P�� O�����b ��R(b�NF�.�D�1����T�X5O��տ��C�sQ\�:8f4�1R:�c�7�6= GcT��E�L3�O�E3�
��}�l	#X�
mm��8� K��6�>N����4�:��t4��%��� ���B}-��,|	�.s��ҩ�z8!`t˞��m܁�ÐH�x�2ڔLM⁸���>){(�P�^�"�U��O��-	w(��19��_Z,1���K���4�w&��AӾ��͈����$��%�WԳDW$S]*��x\ #�K��R�l��Z���}?�i$;^9����Eެ[�+���9Q���^�JEG�|'ϖ�$X�Ӓa���j���j,w��Baə}B !=zv��>O^f

_9*��^t�P����;mmA� ���CB�E â��àG�@2R�h�Ģ�DU��	����Zp�Vŕ\V6T�x�\�;�|&R�H�B�w�ۊ��n��2��/$�n�X#!O/�ॴ�a24dg�e��9�t��^iI>8as�=wd4@2v����t���?�w�ɂ30/k����db\� ����ӗy�VZم����Nv�<�i����X Hq)�=av.��-��?s�)'�Xn����8���B�~�Ϥ��X�d�ٷ��i�y��5j��U�kj�]�ԗ�s]�Q9�? N�����v#�g�	طW�a�_qP7��6�,�8c�+�Z���ӈ�9J�s��M��<"lw&
'��t�J��O��^�rYn:���TP�u��@��h�yZ��?��̕gs�=�8��(���-s�q��w�$���ʅ݌���+,"�L��Hm��, Z֣V����!��*���w2ǿo�=�S��yJ�!�����_�8AwAʝ�����zm<X��[���]����ã[�k�DCH5��`��?2��b�7��q�U&LP��W����p��{W��x��_ڰ�f��X�{"�����t�������]r�;���WC�o�@�	�^�G��SE�MR���0㾤�3@�0Gb�LU��N�q����-�9�j���M�]{ ��]���#GjdE��v�[[�p4Dq�i�����P��}\d'�9���aQ�u����1�V,f�����j�~It�=��i�#;�t��W|���t�Qwm�ؕ�o��O�i��34)��()�UC�n�yh���l����YM��T�o/�[T�Qb�Z�.FZ�\�w���3Σ�.�C ��.�H�+J���鯩����S�ia,|�*����N���m0#S���4�e��[Mj!b���Ra�g�bm�sY2i-�.qJ��__eM}��4t��1"g3Y3I��ƙ""��]k�;X�'�5�A@ycG����W�6�ń4밑m���	��l��K�I፽�� ��\_(�M;%o�m��4�W�I�jo�r��G���Ȥ!#|t�P�y{�q�)Q�1�1�b��и;ҳ��Qm�)'�����e��c�5��=G4����������<)_�1�k�x�
Cm}��G���Q�'`��(Dc�SĬ���Ez�SV����|�\O�$�~�
G�����wcy��wlK|��a��]���m��<��fK9@sΡ�q�0���O�m	D�>���Dh��6:fE4./Κ���0���p��0�b�Ycw.��-Z�-/<�9,�t����0��&\ �SN�C6�%�'٦�=�?	���<R��W��J�N*1� ;1YL����5$&g���5ˣS�6D�́ځ���z�I�,&�e�\~O�Rν�e���U#<�����5�n̔�	��|ܤ�kr�	�"��.y��椅�]��Ϡk/*�����yv���y�nɚ ��5�i.��@��ӡ��/����@V�",%�lt/�r�F�� 96xa��'_���݌���l*\��onԠ9�����0�k�����~��F]Ӳ1^t@�T��D����̴d�j�\EWF���e�#����A���T_zPfF�l���i���t��I�,?������$����G�SS�ѡ�|p�����w��#�NG�?��c��$"���R�ɦ2� (�}!r���ۡ��>`�bge�a1�k��a�-X�p��ғAV���9�|(k�pFZ@S��-p��7�<�EC�Blգ�i��sԫHK��e7"��Ae9�!����X��y�<�B�$�Eֿ�{�nh�?t��3桧��f�~H*F� �COsˈ7�IO���S}��%��q٥m�U���oZ�5�MF�t��|GO��F�N �JÕ�������$"� �A��"3U�� ��n�PY6��b�i���(0R���I������({�ɸ��;;��f�������-�foz�M�ϪoT:��L�3�K��u�5)��rִ�[d?���ҥ�n�f����Z:���� �ݒ[Gf}\�ٿR��%ܘ}`�5%��Cj@� <=-!�{��W���A&j�I�0�?�o�! 	�=�~��
4y�&1q����?62���@���7���Lv�d�H�1�4��u����l�����(��-l�:�H|	yzi�D#:��	U}�ָ���	��Y�n~2ɪ5�p�P+̥��̙[[A���~~nG��~�&��]ݡ�VB�5J��Ek��� �d�JƊ�?N�y��J<��?����z�`�T��J�R�h��`��1�lħ49�ɴy�/&Y�^ꃢ{����I��C]\�Xu=��H����q�B�0PE8���2�ǔ��W�m\YЅ!ȃ�a���.��Ʌ��"{i�<T�h����Ŭp�y�4�O&��z��2 �/�X�����"Ͼk�G���v�2���R���R��tn�@���ma&z��]ߥ�X�L~�����PF�>�$�DÒ�ޓ�6��p����v`4�~H��d��V����to��s|g�ߔ��Қ�/q��%��\���ٹ�g�4WQ�Q���4�dH��ĝ�qL�l|���~7�Tڈ~#�Xga�z��չm�ni�:ơÕ:��p}zi��m��]|^X]��a�,F��H;9b�6�*S ���,��s�TA"���gqs�N��f�-`G�`p�E���@"�=­�u��:=0���9��;�ޫ頿�K	��2[�n�}�2��p���S�Q�c�9���Hs��0����F��0�?����f���S9D}�;����|�E��̲�f� .1ؐx�Q�����v���������tdi- ����7�������8נ���|]^S�B�9~�7���j���
��1�%l/��~)p{:�hi�dbk���Տ��D���L*�/�K�t��[u	����Ef�!k��s��;�fuK-uW@���F��<EObM����P���H%�j�A:'#nm���Q��W�=0c�h��^u�!��^D�F��2^UmwN';(Tv���<{\f�����"o�W�g�x��4N��-g.����ξ�wp�D�aP���·z楅Kj��������DO&��];���W^.�k�,a�-><I��V���X��x;M�2g(��k�_��������qK��h-�T���zY�g3E)@jъb4�y�����HLQ������
��}�K�GՉc@�3QK��{�Ϻ���L^|��������(u�7�3X8d!��(@F�H�� �4ɱ;��>�/���Hh����z���½JQ�>��Q����g	1�R���*�%�pȝT<I�g�=��&�~�z 26 �/y��b��������r���4?G��y�d���y��se%�L$$�ë)���i�kb�A"���7�V7:�T�ơ�c;~k��.���5A�hH;�y)��n�*B�j�2���b����J�����-c|�����^�f��+N�;k�I�(!���S!�����]�F�﷋D|:(�v8{W�Y%B2:��o�i�*{ؤkm���j��Y:	4�˳b�)����]����D�K����� yB1��zC�_>I�`���X�=u4�FQĲ���t�0�L�6��6ReګO�-$'q%q��?�ݦK
ݡx]&s���E��K=�����<�ɱ�6���czm��f��?,���<M�%pB�`J�ʷ1D�&���(\%bҮ��R�˜�֏AK�'����������J��^�X`�T�4��}Jn��H���2�)G�yMO5bmD�ѽ=~�֘q6{��~�m��q-+��0�``풇��n$J'27f�s�^�$ ����/ �0��S�ī�[��>�?�[ g����;�h�"�"�M�KЖ-��E.�F��+���Ҳ�3-�����^���=LY���N���ڻ�
�!s�SׂH�� ����e�ޚg@��(>���PX���v����ͼo�$���N��N�p:E�T^4�{�=�?�r.�3з�M[Hb�O;읳\�O��"�I�����N�=I�F�m.<ə� �
���ך��u�X��������Fk�.�>��;A �B7Wj.E_w�����u�9�_���r�u��(j���3�L2Џ��U6��Z��mo���Wqm`�SDd��#��nJ�oE�[�L�j<��S�'v�����2�(��1�!n߄>�کF��UJ噖�כ��M���\��l����CE���zKu��.""�Tl�[��~����Z��ԙ�;��er�(�*\-���k��o���<�J��0A�NLw��'S!NO��(�U�N'�`E��v1���=���0�CiA�l{0�s�+���}wq�q�<1A!�FXv�D��}[q�������Ė����f�l*�C˚�+3=�=�¿�xa�+�|����uc�@JMu�P�N$2,?$>���F�NX���P۴ᥝ��<��Ds���,���rj����GM?GkJ���Mm�}�.�)D��-V��vG�#�W�B�u����U�Y?KKu�o�l�9�y���m+��Lp�̇ŮD��
v|��B���)oY�P�M�~m�_ޝ��Zy�[Xɻ��J�r�>��DFh��$�@�,�'�_i�(��~K��~"�X`��Lҩ�y�s+E�����.#�B���h�����֔I�F�x�E�L�5{-�zp�ugp����H)i�ǉ;�	�c�B|
�+�ݥh'՗���4>�z�d��|K��jL`H[I��B��\y�3�k[�S�ј�]X����z�e�5�`�ɭ�EfD�Q�])7Z���f����.����I�&�%>w�J/�ۜ�dM7_<?�֯.eR%�$Z���8�/�~� VPT�����ꁻS�����;�i�Q�y�:m�K�:,Om����/�v��;ʐ2Y��	� M�nj��q��̩j�[8������2�����85E�So�XY�h��^D��ܱ������^�{v�.ӧ-�XI��s�\ȉ��[ď:�qh���㸏����h	�x�.�|,g]����
��Æ�_|����7�zmIؚ�ٝ�Jc��ϻ P���c�,pӧ�MYw���f�Ƥ��!���\@`\|\{
�5ԋ���)ir�-\��|����$�e�� iC��h*��TـB^u�m��5���X��@m:a�����rŜ];f�(�$<�2|��F�,f��v˪,F��������:*�����~�K֮Ҽ1j��k�s�h�V�v�մGPy#.:~W�;eú}ٮ�l�T��۟�/�����K�e��x��|�z��$���^v�Ye�q5k��fQ"��#�����C�~E�8y062F{����|!M�sN�p >W��XuW�"~���L��K�M�d�d�pZ��ʉ�P"S1d�bR(z+���k��<��k��Q>��N�b�s�li���P��9 De�.]�&�K�����Ef��4;�.(8-�#X�1��F�[��Q�\���"��r��5z�
���$�ôN�ed�l�j���0^,�y@OB�G8� �J�	4���A�j�Q�����@
��2@}�WR��5��;��ӽ��~�O&fŽ�cl��9"UTJ�I�j� m��-^�����IpܣE��z'+$�C2��-�����ӆ��%f�;��)�?U�#&i䱭#n�g�}��CVK.ntQ�]���Phؠ��(��3U�����f׼G!���>��㼖��1<Z�ta�3�}rG�������zM�w%w�Ni`�^�9c�
��b9u�/;�Q���T^�&r���B�:h
b����*�������ibYޡ����>5��0��e)�DW�XoNA���&;�}�̰ 쉜|0����$��d�P�.�U�PF��H�A��k9a��Dn߼2S�i�p�x��p,`����a�u�̎�Dk�e*q�V+��z�0T fH�K����\����#r�������
�L��-���.���
,�y6�E1 ��Ȥ!�c���w���.�x�{��`nA7C&3��:��oe��1>jo!�Ɯ^D^C�g�'��[>��U���JQ�|eCb���r`����f8q��0�?ҹTN"o���%AuV�="��I�V�������B�#
�|��K#k���� V�`Oi�����'�Q䃖�Ӧ�6���x��`8J- �3֘K���W�z/<�+D� �^ӻ!˖����;��%6Q\�O��� ܡ�}����%�WoG@v��/�w��ǳ�=�Ӯo��k$2E<v�}h�u�w�1��%ҁZ�x���*�\z���l%�v�SӞ7��Ίݭ)xe�0�[iL�А�8sb\�c��Bo�&��Ŝ�Lw��~9���Ƹe�\�dL���tO�i�? >�,h���E�E�U9C�e_{}r�����d9��c�F �߄�#��1�^��o����o:H�]�~�v�d}�$�G,������$U,�{��¨�^�9j���fJ�J�K�^1{6ǓΓ�*�o���l�j��.�~�6�M-�X�]����ܽn@�4�/_��*���d�t�qt�\o���mm�?�{Ζ���<\v�qZ���������KJ`�}���pVmd s�I�d+�)�Q݃�Ĳ��}Q��Խ���9��p�[)����I�F]ۗ�.}�>�Ԍ�L:�LyܞN�I�dA�0�(N��kl��G֎<��>O�}��G,�������&>����g�7
8'�r�]&���(5*�?�p�t�ڧ妧��O;�����YԷ|ޕ �T�)��,���)}:���]����X��Z�׺^JZF��a������\�d-[���3�%��R'6y+��$���|�e/ |8؈��6����5=^;UD&�xh�.B�y��W�\�H�]��̱����Oc�H+� Ѻm�H�;Fz=�x@'�y�o���>�`ZX��	k����z��"����t��|P9b���!1b�</��\�tm�0�F�S<=�
��g-#I�Q��H���z�������M�q��Γ�>a\��A�D�[b0]VX���/(�i~�͞�?�=��{�u��&�$��4i���=V��eʮj��vb�z\Yr�U���Q��˂�(t���qf�5Tn��:a��ߌ�����K��}[��!P�?ab���ג���
$��E~$�
����&�-+rq�B�6���mxYx��H�����{Oz�CWTӅ_f��G����﨨�JZ�5��ү�+ǂ��*��Xbd�&���3T�ka��9t�(���2S�ιV�e�#����)N������T�"�STN�M���a�&����V�MӴ�إ��h񬄤�r��Gݘ�� b���j�w$�b���<rqBWDI`�?$�!bj�٭���>�X�F7�uw/16])Q���G���A����<��jQ����;����R.�C��!OL������h_�_��o���7E���r�Ft�_K���˓�C���!���:�|b+����
JtM/yFM/���y����k	�{�5F�w�4'�!�y��w��{���sE�,������2N��M��o���܀�+�I�C��]��Ge�}��q�̓�`�
�g<��P)ă����������Ar�|�Y����N��Vp��I��\�_��^C��f��|Wpg:#��5K��UJ� �=+R��I��ѳ��$"P}��D�X�j,�,7kc��-�3=q��%yF��0�e��2�I~�'h��:���Ʊ���(f-T���9��܍F!Έwz�VQ�-k�zh<e�� ���پy(�pW�֓��_Qª��#�o�tyy�i�%�����I�D�8(|�=������p�_}7�7���,�TO9Ƨ��ouwC���JW�߱益H���F)sC����;(�Cu|��n�xo�Pֻ�h�,���#�:k��u3��UQ�9��=���rK/07�)b�D�+������H�t�i~����*^?�r���T��֫̚r�ֳ�z�,|�[-�\@���$��W�=��'���L�%�Gc�wb�$����֏�G辳�Øe��"�Y��lK���)��-�#+`0g�@�����q�rO��%�����;b�:	��Eo���Y�e9\v�őpd\{..���P�U'lG'��i�'u����+�q��}����|>��)��R癫���U&����c#��Z�y�hzުV���;�w�Llt�R'�}�k��=��E��:��ͩx��5���՘����n��c�ޞb��=&'�І2�����F�\o7�,�Ý)WkU6 �Vр��B�)�����qZ������Z�>��\�k;�9�@i�K�$>i��z�� t�N�Hx��U���@�mjeH�=`ʥ~��r�ə�"q$g�d�����p 0�(��m�P���E����l��l[�=��ASə!��&�r%�d�K���V���j�	4A6h�s!B$Rj`a������q��îb��d]1��W�kU��<�S/+�-Oq^z��9��<M1�w�5 ?W\�t)�Ǜ�1�My���>Ԙ�����ޤ�����A3�5*��c ��6��b� R�*H�c�ߤ�����k�q",%50��ɅuA��E'�Q����6KF�(2�6*���H���p�<I;��p¢?X(��ϖ�OL�FSr��=��ɯ�ľx�}��;ӅC��!w���Y�"%5�0�WZk�T�qlp����7Ere� xʘ1`��ڦ2�=I�e�s����/�H��Q�o�Y�����yig�sL��m>�pB* n��H Q�f�I�h�"���F�����fb]\#4"lYq$ka^%K^{�t����:�~lEJ�n�Z�ss��j�ߓ _��~�պ�쐦��tZ���,��<�˥o;̴����Bg�J����5�m2�t<o��O˥�	�;`o�B!U�� �Ɲ<
���w�}�$�=�RU��	������{�x(Kj��t��Η�Q���1�ݥTo����ں�n��o�Q2�g�>$M��ri�=/t���)���S�p=��Fu�L}��fG�;*+�>ц�lS�ے_�,�ya~@��g&��y�s��L(��9��C<��^��6�c9Q�q6��E�8.�D���,����Дǿ��Q�<����`u���X���[���	��ɫh\mMk���T�D�&��.m�K�E6�jئ��S��ܢ�a�T!�4m3|�G�_�t�F�3L�LraZw�7��62�rˀ3�U�D�O��Gd�z9��W���$�����g��c������%�"����,:GdG�/i"ʯHa��У6~!R�D6�l�_"�������دC�PL���=0��5������<���Q]���X��yOk	)惕~LH/���p˜��艕��lL��M��!�3�j�^�TF�����ف�r�p7!�V6#�a�<�9�� N-z�����XB�Z;]�;����h��r��̡��j;��ʏ�|�x4����C��Y穸�k�
�3p�" c�}Y|\m�������i:S����
�=��-�M\��>����cE���)����e��fΝ�1�>�ѥQ�n�V�9�x$x1�B�\3(���c�#��C��!����-�)�n�?�E
�||�Y�1�ā�<�"?�l�I�NFn��"�i���q9ts���k�hc�{4۴�P+����!�F'>���Ͳ�^9*��g%`�t�f��%�+����i�ma*�A�����o�gTjA,N��<��:�C�v���2��'N5�EߋEP�ޚ��Ҕł
�%���j&2�J�e����cJ0�~$U�d��(��<@�7;�I�/�׵��N��+���7�#��}�)��)��j��^�Z4Z�g$ ��4Y�b��:~�z���e��v%yjwⱣ�I�#�>IZe�Z�w���{cz2�R~�PZ��n�5�@�˪G�[�`��3H��L[ig��ρdgˠʛ��N��)n��+��Ƭ���%I�L������T� �{ȩ�T���`���:oJ]�W���XQz	�U[ ם�F�]3r��xoS9\���{x�i０�~��-Z]y6{|cAp�S{̖���l�ƚ�sF�w��{	��v�oc�UZ#<�>���R���~}����n�8f�����K^D_�Ս��慒���8� fB�1�1���f��*�!f�p1���O��_��Ӥv��d�b��'����G{�g;�����/ԯB'���+u~��m��{.�q���P�pTڟ6���q�s�1�?"�2��1�ɯ2�n�
[��L��7�X&�6N�ҩ\�̓)��3�(���H��5�ǚQ�2V�ɜ�:<�˝��u���]z�SN,�Ն`۷�Qz�@��h����V��(���.�V��a��]jt
 ���#Յ���bsG�$����勾�K������[�}ꭶuW��Fy�ӛ�TL�r�4*�B��+���x�d2�VHE��&j��F���ׁ3���S�N�j�O���ƫ���)��c ?ⷯ�)]Z(�3fʐ�N5JB����_�qV���n	��#b�4��v��!���l��	G��9t��_8�f� �	�s���~d_��c��M;Ԗ��XB심R�Iٺi)���-i4�e7�9��[�ݒ�dt=ʇ�+�5�`!+^�eE��F��>ڙ�����_�����#�0�*���?id@�OW�q�E�į�PoR!)��,b7��7$P���7�,j[�����2�Ws"aN��{���d�0�ב���6�+m}�2 G�ǘ�����L)�A2E"���]�{���U��p��^�ъ�KH6{a�N��h����{��Z,6|>zI7�Xm}Vq�9��U��d��=�A�W'q�&R8����D5����&�w�#n����.��b"�:ĳ��2Hm�X.h �5/�O��K]k����/�~�K�mr�(!�c��p�&��� �C��}M��f�n_��G�h?�|x�E��mD�֘��m3W1���Ѻ��������F��H�2�q�@e�LF��lr���U���akf���FL�߳�R��0&%3p���P�T��^�(t�-�G�ċqt�)<s����~��/ р�W�B�P&ت@��5��)�꠫��؏��in�ZI��2z�������8��h�C�T����2�"�䦨�f�,%�d�u>,[o8c���ٖ*D��v��eK@�i'u�i�$1�K&�R�}>אG&�V�L4�]mwgm����3�{�)��� 
q}�̠��<�U��Β3Z��c�r:v�Y����l�]��`� ����aH#�����������J�f�D[�ٞ-3�ׁ�!;`��u�G/�<_�­֊�U�Q�]0ߢ�����J;��x�z`�W�+"�m}yEk��.�-D��)��T�&Ev��rꎉb�T�/rO�RP�S0����E��=4���)[�Ȅ#�Z䦺�����^p�2�MC��v�5ɋ���߬��@�&�$-�/k�:;$��u|�+�X�tӦ�I}(70�5�6����g�����-.(�, �*R�l/�߀ߨh%{�5s������b�$�qJ�s�]QG�0����!�&��r�=��q^N.E����޲m�^��<�Y��;���r���!��۟�����E�ɘ���#���\|�׏�1�y
�|�Id�d�K�k�v�������:��G�62��v�&D'�W�>iS���r�_n��+�lR���ڶ�0�O��DU]�ʋ}�k���M�]L�/qA
�9ҿg���Je~I'C��ƹ�ߙ�̂�rB�g��w&7F~;S`7ᵶ�� ^"���b��@H���2e
��m�iɾ�3���K���:��	��/�,5�Mlo��G�s>+��/B_?��}Zf��2�ko�5� t.ه��bEM�X�?&��g�E�}��xS1�2�6�\��K�Q�܍��x�b:y}��*�Lay�֟����S)����߃o=E�O[�mjtv���'���b԰i��Kx[���*�.,��@	��� >��rNf�=�a���2���I��~�,qS����kZ@�0݊&,Gz��>�g01&�c~콺���#�0�������af'��K�ֱԽ�|_�i��zu�hh���[�����V�ݓ�}�Qۤ���a�9
�wǓ��Y�:Y�t��e�8gI����na_���"���h+��}�2oSx�3�� � �9 v���S^�6�����Z��b�4��M]�Q�L���LrO�})W�x a{��5�,��<��9D���ZLH��ȀdlK�:*a�$�MM�߅��� m,�/ͧK��RBqƈ�5T6�]%$���
+��	Rn]�I��vy�)�n~�bذk��:��F�Z�,�"�-�#�w�Ǵ/��4�v��qW>�/Uli¤�o�=�1":R4ƨ�Gd|YO��޵�_3�jP��aK�ي����0�g����� ��4��l�Ҙ�w��0ߺ�7I8�����g�c�4�|���`���5=z��ȴr�L�����O�`G��qE%嬘�8�U����0.[�����W��B`{���O��)i���P�qH(6�a�����B�a"�TN�J�8�R���p���P퐤NH�9�� j��(����}sP(0�q>�K�ˮ��(��#���Y&]F|�/`�.����=�Rl������ۑ�?.p��Q�HS�@*��Z��X��uuFd��BJ'G��D}=+������s��S![��[�ږ�7���xP����ev�q'|�/�9R��J�ğ�<��'�s,v�屺�jEss���`
q{�<������?!F铀�ۂ�2�
�u���{�ه}.�^4n=K���bI��t�=vm)�N;�=8�%���<�#�2Y:��ۜ{���]ԍ]�����CY�I�Ł;*���y�#ҭޟ���p�9���T��A�أa�)���&)�0�8�*#�.0�<E�׸��K���}fX}�\O-��f Oc����=��$�c���J�O�	��!2���B/H�&���,D��$LN;��_Mq�R���/���]P;� ��D0��p�����]:V�r��	����߹+��d}�3	+p.�q�ٛ�*--;���l=��c��q��:u�
���Ǣ�\�p�'Wv;�;�{��3��J۔���I+�L��{���	|[�	Zb���V��s0>�O�IH��N�=6� �B�%��(ƥY���f�1)�IEא���/����SQ�����(!��i�JQ~�S��$Tb��^����U�g�e<�D��\%���jS��>��A�-�2�\�؂Wκ���=���A��y��ԍw'MH����C�4���	���	��+�ujuk�z��A<��|=���U�iHi�����������#(��dc}�D_�k�"�V�Y�?�nE�.�(����n��aǩ�Ix`C*O/�a���W�3q�&�������4��S��t?�0��S�R�7�xy {�P�8h7xR���ؔ1b�1g	�\{n�� [+bn�C����[��������.�+I�Qm��?!�������J@kv��R��;!nxT��ce�ت�E7���Q�ㇶ��K�r;����b��bH\?�o��Scοa�i���m���?U<�V��������Z5*.a4}�%b�|�r�U��6Z�,U�m=����-t<<J�K�ٹt:�m�Ɲ�v�h]�`l;qm�o��y-0�=�rE}��_TNb�)̄��Ok�ċ���1-P��ވ�+4��%��u�u+\��0���XFӌ�]~J��C����n���=M�4-`��Ifbf�Us�㫣>P�;��j�����V�|3��Bǔ(W�������R]��!�"���F�7_@AK���~�8�c�U�����'.��C:SZ�a��li{��{���T'(���%&�Q�M�4e&
����l�ƾ.(�7���8�5�J;�YP�����ԺeX�sf�F����,=9K!������	Z]d���uJ�Ҋ!<�VIS���*���g!��*������Iɿ$3+��m��\-��*SK�g��Z~����ie<��	�u��*]����ۂM���=u�}��on1�lK����k/U�Z�^7���=� �'#��W�H*�ڎ`���P���,��Oո-��[��U�V`ȭ�S�"]'���ȕ��a��[&dLo�P7����zi�H��0���������Օ�H��]��XE>S��g@NIDs�J)h�W|�94p8�f�5��HE��d�1����=|+���ѭ���/윟Og���֦Y�\>�g69����U3O�bN�&DW0��Y�Ee�b�Fhb���=ܡ v`��Kn���꫁�tG3��O�3t�K��iK|r0�p�s����w�U�|��ь����b0`�v�v0F���?so[k�6�aUMU1�(�4���e6����L��}&]�D)� Jx���Sh�ٽ�Ș���Ⱦ�l)�ّ%��Ny>�L"�'������?yc�	Imo���6E��¾���Ms6��6^Mq`�:}�P(���j��J���eh8z�Un�l�#��Ƿ��ptA�w��� l���Q`S��m嶗��1X4k>4�½L?�K�!�hZ�ȫ�����>�)�pG�x!������ӳ��3ΰ�O+pY��@�7P����wG�)�p|E����bzπW.�a�d�w��u1銈'S~��γ���J�;Z�
A��#��� �Vٿ}�cb�z<.q�z�|Y-i��m���Bt��"����9�F��'�K8a{ ����}�ڞ��S�ר�P����p(Ǘ�v~m쮔�xLOI}�u���7L��W^��zQbsߥ��5UP1�M�twcUJ���N9w��6��{L�f�X+D\��&�q #:3�������c@�hys����-�<G0/���?8O�]]��f?�eO�����٦���tY�c�f���7�xL�̓Q>9%1c�[��륮;5ڍG�%,�~d������[M�Qzc���� �O�M	�ޟ�9^f���GNk���C��(?W��1����n'.[\�"����]WW��K:�)K�ۻ�J�HA؝�9�-.�ʨ�����ϊU��GA-O����ˆ�v{���o�r�K,����%�Q�z��K��%��R
E �wЛM�g�6:�>qP�����+��
�!%���h��B1�]r �h�4��%��fza���X(3P��Y�e����â�3h���]7����Uf�&���P�Mҩ'E�L8�J@H(E�D���83|pf�������"���(s�}��J7�C�׼���[��^0S��c��7:���_@�|v����e07��L���S��ndjPg8u�$=�GֳIH�a>�k�^���  <������]��[�rX0�_�W���A�����9��r`~J��&���dw�5�V+��ZG|�	_䂺�7r�d��w��M�L��AA�7`:�6b`uc�ҡ@#Q�� t�:aZ����+T��?����mӉ����W�0J�d��;2�'���n�[�zy��O�Γ�b���P�m�%A�}������!@�)��)�ŋ���]��q��k��A��Qk�еvz쫅xS��9_9z���~����}��`{|��p��l�K޺�_��چ��D�WY�eX(͛����	B`�F��ֽ�I�в -B�^�q$���N��?�[HD������23vm�����]]�BfGg�`��l��Ԏ�m��H�1��
E������8�������ͶZ~�j�75�������*�:����E�`
�9ݖfj��rYe�j�%E�k��q�$ow�����Ddu_3H���[�q`K��*Pi[m���KlgFh{�}5��x2�P����娉�Jss�s(�^����%�m�`���0o��$�&őV�xV�>!6�31Wx�H��5��o7<
b.yh8Z���~�Wy=�J�1�Q����@[o����
gxC�}�5��R
{ ��}��� ��YڔlO��;<뮤��`��<l;���Ҋ9�~88�ƪ\e;��PB ��M�+?@}�B۹5�u&2�f�^J�r%����n���0D��
�p	Z��7�v�����`�}%򴘐�Y0���7cWxe�3 i���F���QrE,n8?�JBP+c�=o��֫#�"9��_���9����Ņ�q�˃G�7���� �M������-\��� s���Z";��lc�]����%�)�X�,��6.a DQ]������X�ܩA#r;SǙ螲�V��k�����󇁧����)�v�2~^��!ѥ/�,rK�+�c��1��q�7��\�0�E�!�<>���&�i�� ��h�Ok�0������T{�U����Z��u���7coƛ^�7�P��VΝЦ!�Q�6�ȝZ5��]wa�z�!ṭ�j{x���S]3@���M�������Ciz�J���7|)�$�N{��X�+_��S�U>R�R�*��L.�Fs6�Gd�Z"s�G�����}�|�/�Ŋ	xa�<P�GS��h��"�q�+g�,����Wt��Z���"�d��cZc��y���8r(!�?�|j�ê�d��b:#~��,Zַ��D���[���P�PiKC�� �M[/�͞���"ie8m�=�˳�(���!�5���	�׈�qmf\��Pά�TA|Q��	����&:!.h"��V`I���>��1�P<�	+d�>ހ����_����F��>ݙJ�`��Rb�@"3ٛ�Q5F!<�SaY$Z�P�?����celj@ܜ�C�w�-µA?7�D%���1��jT�B�>����+����7Χb��3u�>Vu<�sQ!|ۣ��jW�"��R�;v���l�-���F��.�7�k�Vϔ�Q�.<ف���+
/��V�PV��	=�K���d	hI����[���=b 7X��l�m�vx�J$�2{_��b���}n+Rz��#m�;��Uн�/R�V����v��ĭ�� </�f�%�PM�V�'���~x�a�ͺ�j��Y�>�Uc�sx�	}Z�~�s�it'쟚���Z ���<��ܲ��[z�\�|�2�8��Je*;�cPJOsZr��:ւ^���2�1)�m�L��k�-�X׀y��[�l���PD���&��~�ԋ��s:��0G�f�<#��3x5���4�d�1_1�ݲ��9v���Eg.Bh�� Y�}��o&�Ǻ���0�|S#��V�:�� �{�D Y7�'R�E���U_�hj_��$����#Iݣ�W�=�M���v\���E;���v�2��Ц�M��P����bo��>D}���� :�ieզ�#�Ǹ-�̏QF����YL(�%|���	�oKu	��	��((#[sv�zK���m����j�;�U��G?w��*��g
l�ct_k�Z��k:��.9A�λ�TD���'7��\�y� �c��֓iZ�M۽)ZI���I�{"=�ӲGd��=���_����H*c�hs^�u^\ȩ{VS�<��\�eI���F�$7d��*��� {!;ҫr��qڀodZ0#ȉp�sp����L��������#�"���\\�q�b�܎4�6�"��w�:���I�P��߷��� ����+�D����~H�����X;&��#�6�	���>��d��S��,S�/��`܀+<���+�L�p
�R��t	"J���7�;b���I഑���=B#�u�S���)w�&�%���S�皪���؄4H�%���kW�A6i"4�E�G����6/�w�șpa�\�ʽE�V�c{�t�"!�&_Ϩs�����R�J��)��'��%���Ҡ�wY��	�+���WU�*�n/TD�ߠ8�'�E��P��*�h.�61�+`ݺe���?�R�?�y���c (�~�3��ӹ��Y�Uϳ ���\k�I��x
)w�,\,�799��dڄ��k��C���\Zyh���qKW� >�h UN�%bP6�f7X^��E��㺿H���R��m��#ibH{LPr<��aXk0z��RM���4;2�@����Zh�z�H�~��4h<�f����fJ����&|�OS�
D��s��RA�`>d_ ��@�d]��K�SPʬ�i�y����<$Sl�Z��ks���s)ASm<��Q�4M.����H��Pa�[I�"2?��vJ�����Q�`!�sq�3۝��4��rt�kO�N@Q�����Z�m�k�����x�N����j1��M�˩���
��78�F�#r�[6��8%��VG�ZG�zk_%�Z�,�=�Э}�0�[ x3-���V�X�z��:�����U���&�0��������~߱1�Sԭ�R�ЌzXe&`�r���Z4e�YfA��"'�!�A����m�8��	���V�k�f��茀.��D�[1"S7�7�Z7<��Nt�����j�|� ޓ c!����kp���X:Q6ꖡ�Vh�)$Uݏ�Raȿ6��#}�
G��c���[�(���9\h�+c�;p>X�����ZH���qxK�9��{.T�����+o�&:��R.L]5dG��}�{��hqTu(Z���42�7�1^�I��*�&��_�/o�3LUG���q��%�g���d2�7�J3Y���>���O���A�سpI���_G_5�&~����L�y4M�g�5kE��(>Ů
�۞���Z��F:[���%1e���Տ"CS��}6�����S_V��Ή�P+��{�9�� S��5t2�;b�@��8�D�I��*-@9�F[=�)�N�$�X�HT����+ �"'&�|�����|tg��H���i�Ϝ�Mc׭�=����>/��cg?�*��~�U4�m��O�ZV|���=��JV����&��̙�����i���}E�m��L�K����r�,���!�Jb���-Fp��7d�f³�8F���i����P�.�HXɊ���Wbl�/ 1���wU��%�����G�Ɵ�܆ϵ�h�OeFw�z[��� �ϛŕ�y"~3X��,Ӊk����p
#��z���,�lqt�i�Z���ݕ`�]Y�u�nI��!N�̼�#_��޴pZ���4��a3�0�	�⍩�#�C`!>��Q	��9�؟U,n#L�PǳG�bAf-
�PﲨK|��iN�1.%���27���d?�����o����L�=�|5�߾�q��a�����޺�Rv�wҫ��N�2l�J/���"���� ��4,��!{�����p�]�T���J�}�V�,bf���q�0c,�[o�;s<j~�V'��5m��2j�ٰ�j�9X4l��|�s����;1�z��e�2.�T��n`S�H8W��@����z_@8.��~=��Ҳ�`�2���]%�?i����)j>��u��L��AkΏ,m��-I�M�QOԺ�7��Y��e�甎�wm���)���i)�U��H'�� +�$��s����$�d}��gsI@C��ǭ�.��6��8��bQ1-{-rk9�"�N8qЂNf��Ē˓4�2۹&3o�Y��Ҫ�����X�}�x�&�\ �ĬF9�ZW$G��=8�=Q�+�A�O�電���I��$��A��D���̲��3ܪ�� p��{,'A�+Y��+��7�=_�w̧�38)Ў�,g����{�����j|�5��ں���aG�َTpu>i�1��/w�!{��1�`?)qg��A�_�P�f"x��nmj���zW�oC>Q! �A��gXF|��ra��͖�����ˡ(6��I*�@�7�H��h���y�}�jt�v8j����i�2�uC쿁����x���9�����зᦷ��o]�%�-
:��(�TBFu��u�X��h�����bew��j��Tј(�Fﺩ߈�p rv͕Z/�ֺ��*�zR	b�q�,�6���_��0��vBf�:bp��=s�(�HQq��L,�u��oEk�t����(wH�K(�%���R�i=/�s���|��t�� ��l�~�@E�5^��wcP	E/� ��}��>�>m��ԟ=�X��I��J��C���}Ϭ�o{�C�Q�����/R����W��{˲�mwŰ�GP���u��U�k���^@�<�����6���,!\	��������ǃcg��갉��z���_Ȅ�+Ѫ�''آd����-�L}T��@>�&�'�^R�R;��~�y~X��aJ�k ������8�2b���(� 5��;���$+���*��5���t�!��{9wi]����|#_I/WF����x�����l;��2/ަ��r�$��{�6t�V�?�bZ��NV���`�
A`��X0�aᙔ>�"G>d��և�((��bV�	���B�`R���2�7��{�a����p��BGf�Z�CΜ�TԬ��k9!�4|y�+�9ꌥ��?�6o��;�:�"(̊��U�_ߒ0/���Lk�[�/��mFW�&�Ύ��NO��\Y���'3'��4;� 	>�����D�˙�ĉ0��Mh�Z�l�!���H��T�e��24��]�|��1�Ɯ��?�����Ӏ����]���*�|��G�N��0�qT��dò�پ��U>*�����B��%��{"��hy�8��.�!��4���	�MMOnv�Ԉ�J;
��9���w���W��t�5�s��;��,j���`�i���i�E�Ń�<h�2��zv�tyF��Ki�p����AI���ynn�� �(l���1��m�9�Ɇ��t?�>TE��tK�X,�f�^`���a~Px�O��w3Κ���G��ܯ�![!���Kع^لNkC�O0Xg�}�5����癬e���[xGbD ]�f꧂��������<8�ͥ�eQ�Ui���P��E��i�m	f��^�ZY� ��w��LV
�\�F'F��T�=~�I!@3��O��&mx�8�`ZP����t��4��e8<Ihۓ�߭V�;O	h��u�}\���Gnƪ�����@�������N��rT�M�)#G�SU��>�$�U�:�;���~�l�a֥X�PѢ~��f��W�&�o�@U��u�ەY\�R>'����<�	j��)R���r��yt��7���5;��	V]�r�_z�$�&�IO�t.���jv&A�����c0�f����ş�F��eTj��ʨ)b-KJK�qpQ��޻b��}���K"梠���h�&Ty�J�I�n���DdJN��q��^��E��1qd��������<�I��6�L���j'��s�z��o{������"��:�+��$���1/$( FN�-¿�v�ZN�p�e�]�"[��'�hh�����ܠ�����0�C��li��?t��D%O���LEm8��@�(��/KX/� ��(���;׽�͡e�Ṙ�Ҋ@�PŪ��VIO������|�K���Q���4&3?A'�DP�{���˟1z�/ʬ��_H�� ۸���U��
�(N\�ԩN�} Hr��I7�h���M9�����Q=���tVjw#5��P���ڧ��u�9/��5/�@5Jث�E'2Ѹ�30���N4_�=��Ɓ���k��p�`�V��@�Zy%s�6��p D&^����i6�ݩ�3{�We6�&O�ǋ_#���L�Р�D��)v��USǵp��k�g�S��A������Y�9�wZH�2�.���F����#E�3�D9�a �i�g�/�;��8wr�n�G�e�7���/?<j��k�	S�/��
Hk��U}�ǟ�ձ3ں��Df?���A3xO�'�9m-ޏj�9�ҁ�]�|������M����W���}7'|�zG�`�M� ����5K��c�B#8:y����r��ށ^���u��y,�la��t�~?�V(�~�ZY�Θ��2/���ӊY�GzT���jՙr�m�#ڃ9{�x��UnN�M�[��gq-�Pծ������Ģ��_�Zn<p�u!�����"�vʭ��+2��'m�(��)R���cAwq4�t�	Y����}io1f�������a�)By�4\Ei��_<�)_2;��^�<eߨn$I���;n�+��MIgs���bo�!���1���8W��
���BQ�i�O����8F��u�'�:�(+@�`ܹ�84���!��Kn��!F�c�w�:�E5��t��iۉ���׼��C|U;l�4]��s{�������0��Lӫf�6W���b�D~���,��3:`	B�����ִ����]��;����GA5�c��~g��Lz"�	l }[��~�\?�����MEچ~BY��IX'6{���`�˘�c9j!}z�*^�U�N�uƘz���豀�:��=�ztz\4�9��	z����eɂ '���>���:�ݚp�g���ZА{L"0|��y�'��YI�a��7q>�&��
�aG�̕�{��m�7����Vo�� Z!-ä7w��Ҏ��fkUI�ǌ��� ��m�;����#�q��aV�=�����o�ؽ  �90���4F�b�h%20���Kh���*���Kq��Ǜ��_ܜ��<�q�Jͧ	�It�5�o��y>�I��5aD�k�a�#>���N^4�����v�7��LN6޵�׼uҔ�����p�Sa���2@J?6�����p����������X��v=dx21�;f��_}r�yC߰+�|�k�~�C���t#:#B�om�K!��fw�����.�Ș) ����s:5��ھd5w��I��J*��Ɓ�w�E�w����UCF)�%����n��	}�bu`F�B�R6����7`�n-���r�by
wH��ډB���Y�\"���yd�J��6:ז�o�����gi9̍i1�+t��:�@G	�&`��:� L�D�(&h��'�kf[fQ�-<,��0��!�����S����.������*��g��6�2�m����CۂP#q��U��Ԛ�[�����d%l�LX�͝�����js����x� �| ���1�����Z�B:%Ok�W�۳˴pt{!f�a��O�8� O�
P?O�����,�T�6Ab�&��R@<V��$R��Q�<o����
n-��z�R��22}����@����@�7&0��W\��Sy7,����@=��+���.�LF8m3��&Z�%�19k>E����W��5S��W���|ǎ [��s1'���L�¼<5����l_���$�����ũ9�7�g)dP���k�
�ͩ�_"�y@�/e��T5���l��5������&��&)u�M�|�R�,x�K��7��lټű�ԉ<q�$Ԥ(�2�$�jf�/0�����r�:���gsW|�#�����ש�0����x[$Û�KI4��48��d��q7�\}7��8���B���!��P�������^!�1c� ҹ��xX�pNPG��Z����ÉoQ��zi��d� x�ml/� K\��\/}h/)��ؠ�,3V�9y�aS������� �P�sٷB�g\��4?�{�#z��Tb���~�~�$��]��t/�=� ���^�="@����&��sTɴL��: ��<p�)�$�ċ�2�(R��2��8奮�F�H�Ky;wV��M;$}�K8}���1j��=���y,Ԕ56����[QQ!ND��m�^��%�p����3���߲���[X)Ĳt�Joԍ���{��0�vOK�+�p)ZI��8#�ئ�V�1B�d;=��R4�t[6y�L�@��I���K�h�-�f>�R��Dd�"Zpc�>����xh�%�/i�|�.cC���Q;�>�'J����8mk� ����o�dQ� k�PA�����h�������C�r��N��tT��4�5�/�p� V%i-v9p�$�(��U���(إ�q�8�:��O)�.�&�9��j�Q�.Y�>��M���
��8��C�Ϙ�Q�����@��Ԯ�����{������������%& v���s��0����L��v)��U��7��3�/��R��K��Ӫ Y���aRw�o4�Wq�a<�]�v�l�9HĘ�L��!���9�|���|'��N �^eW�/~`O�ĥ��Ϻ�By�HP�h�����
{����vs0��y5ҟf�B��h�YH��mm�X�rrL� �b�j5+����Jk��³��R4R���ć��X�5��}�5�~�avL�6�u@�8��ټ�fA���H�
 5�������TG�D�=�L:�*ءثoR�b
h y�m}ORz��V�
?C�aΎ8qc�,��tv`oi>�%B ��8��,�2Dد̅�"�N�#�����2��^{���,v��flꑚu[5t�况���O���e�� ()^QG�<l��5��wZ�Z�:cLJr�S�rqX�f� Os.w����:�#89�.'ަ{���� �aaB��vYV�`#��SAM��
��JI	9�(+Z��1��I�g)�C�K��;�Ciw~��X���C��:׿�������#c�㬦���#�oF���^��el���6����Mu�#����gp�=˺���g�ſ�C:^��~���"����+N�\r����Ɨ���2��N��2e�Ť���~B8�㧭�~�2�/��qI�[zA|�v��[H���[�?��g�+(b��n=��X�J�L;	m;G�Q� ���eW��K�A�f�~lc�)���0�������u5É�<�l��������uvE��u)�^k����&��QsЂ�������7���̤.R�F��i�e�2Bf��bH.ƻL�W13$Q��'�����=�/��)m���v���f�,Y�L5*�d,0}����9�3��%�D�Wݎ7ꆁ>�:L�Wn����tH�X92g	T@~_��T#�AY�,�gW��H�
��q�e�D�9�A��<��j��|,��ğ��GE?P`QAq�\��hF;מ�f��b	�*Ԅ���45���:]�N���_˳�g�x,a���	��ݟފ
<#f�]�tJݏ��W�Tl�=�i;��cH�� ��9�o��Nhd�M�p���+��;���2�������o�(j�%�!Y3�v�]��r��`�j���� �t�Sp$�Cx7j�E���.��B�m�(g|�nW*�0q=�}�~��k3o�Y�,�{����L���#����ngZ�V��N�����fj�T�}ϊG� �z�5 �޽߶c|d��2�g��m-\�{ز�4g�&3Q_���Am>3���C%�89p��fް�Ɇ��ϛ��V�v�Z��:0+�'� ���r�"� ��k�uZ���?g*c��+)]�b
�z�����Kp\��:�G����
�Ѷ[p�G�~�K��׬=�Q��u�2� �@�d�j1�GD�/ ����L�"�DV��hm�K�O��]q"�@x�v��?�*B���v�W0\Ab��D���T�|=U6	.����:c�F�}��C ����HL���"\H.��^HMg�ރ*�Մ�����X��Qe�Yġ�(F�.fnk��ռJ�������R��]år$p[��[�(����\D|��=4ԃ���;4!����u��T�%XX|ϋ���7Ȭc��׃�I����:�{��{���F��	ڥ�S�MϮ��u�P��Lx�_&׉�րʪ�q��<mڋC�Y5�n9|�S�sY��[�DS^�����ÜyUj�
���[H��"3��<ۈs��eʤ�}%P��X��8�����&F|�-��S>1�H�ͱ��V6v����v%S��)���g���zZ��|�u��r`Ϻ��o�-)ћ��^~K�O?J�	fs)^���8�{F:���",�ܢ�򰞃�̃K�>���)�ܐ�� ����g��n{໫
��=���Mv�&�#1�C��t��c�� Ҝ�:���N��'֠^\�X��"-�Bf�_��ƀVh�8]��+��]��6���!Һ�f��J�g�ʭ1Z;�@3ش�BבּB:�W:m+�%�]n�G�v��i�I���l~a�]�,2C�\��1(�d����{ɕx`��Ď4��Nˎ���.W�,��N�D���I�nsY�mկ>�擥��$��a���`�����mV���H�>~��r#�M�Q��C��za��~Us_utr�n�0�R��d�I�80��`XE���hS	�!/\�r7��tC­ߌ������x��(���M�����K_�?n���f�G��Ew��(���@��L�k�_KPC���������#wyM��oY-��eU˥շ�r�pT8�G����d��n�tv���Yf�a\�H�� ���ᅯW7���B&� F@p@0w�*�l���w�s�}R���&Ǻ�S/<�aט�K�-C��g�~��0�� q:o�lU	�.kk���7��>;,+۪�{E��K��f�3�O�����i�omS(y$ F����]�
����P�����֕����#�Fvs� 	(s�Ra0�ĎK��%��X���� uO]�l��i��z	�sG6$ȁqB��RJ�8��S�� �c0�E�Q�WN��wx��pܔs����d��;�B��X�#@u�9�����������a̭ꜗ-/��#�;�|f_1
�2!�m6i�a��\B�YT7�/]�8~!���#F t��H�ګ�c�,Z�b��l;�(��R�38ډ�YZ��9#D�9��@rF��Igc(���s��&�+���E��G���V�	��vr��Z'�� 7�8�� i�W(\�.��gK�� ]���\�O���I����B���u��#��|��F�����z���`"�~��$�G��,D!��$δp�\i�^r]�6�X�v�E}q!�`���$>��<�C�C��,�4F��n���Pfmo������-�vNG%�E�s�9~.h%A��7s,
���n�%WrnJ��K�#����٤F����sU� �q��怶'��'��
?6V��!�Ko(�	��]0=�C}���g��_𛉰:YW���&-8�������XJ{r�F��q����v�Ώ� �b j�:X�-�;�H�J������}���|C�É]$}(A�a5���/�8����f�ǃd6�@q����NϬ��([iHE��<�9��6=���������|�5r<43d��5e�o�rU��Bi`}���q0ߌ��8�]cCiY��I]��:r��u_/@��SB���}�K�#��D����BH��w1  %ʵ�*6�M��v:	�-��˫���l�^ȫή�^TR[����ƒpAS�	��°����j��ᷭ�B�h�QA��/��;/M��55�CX�h��.�e��z ČFt�]N�Ĝ���\�m$���)��F q��W�G���c��4*+�d�#�n����Gbl�C��4r���t���h�Zf�9YL��VH�w���;�^;|hhe�&G�X0B����c�<ȹ&�w:�e�1���T�D$(*�p�c��M���;�zC���Le ��� �,<��ɒ����zӉ�P���ű�
B��M~_İvQ�Sh��Ԉ=z6�I�u����8]ke܌O�#�P�js�5�Z����֏�M�:�!�Zp�����Av�5�My�[��@)[VI�5ʾu�]p� %�ǝ`��������}�q;����b6ȿm��;[NӲ �)���&� �᮰�D><��������5\_��zU��x����_����UD�';��PG�9w둛QV��ē3Ui��s/b�E�<��2�;� �Tq'&Ͳk�`$FV"V��g,�f�]I�Z��;�E(��JS�Z<��+�50~+�����q����YY��ڑ	��,2?H���E[*§��ۮsb?����C�L���hń,���1� '��(��IW~��H).��%,I�)�)�~bb��`��F���g������7����b���~ft{�Q�[(}�ÌQM��OY��Yʠ���FA��vh��C�)�J�fS� 8��t��6��!!x���ih�Pj�W���NAIwt_�3�2�6�Ϳ��:�U	�������@;[��a$�N [��B�� ��v汌�Dq�:�V�]�l@0����ᔦ��l%�;>6W,�g(�ޤ��(&���}:�I�$��7F?�d���|�;���vB�����.F������[��8�p�i(g�ۃ�T���N�"!�u���d(��*��6񘠜1��{D���j�,O��с}G���$.x�{�,;YL|��M:��S���>��:������`4�iP��-6�r�y��󔷣1役@�[%e�_��[S�}5u���J��f.���.����4a��R����&C�����?������%����K^n�S���Q�)��j
t{������R����l7a���g0�Q����Q,�o5����P"�R�� PXot�H�&��Sai+��,M7��B}p6͊�\t��5��ҵl2Ɠ�'���niC�_�������'���sм{X ˣ3��yP�|�Z�Bwoi`An�+5�	�]S��yЩ�xq]�I0������/������uY'�S=�,y�W�"R���<�Sx}�ׯ�e���/�<���5��v1�?hN��;��$Ӵ��,e'�AI!���Hf�]!hF��a����7��rٍ� ���¿��}������fq"�����iH(x=L���!͜�{�Ta��\���	�������Կ<������2F� }Ŋ�=�K,C5���aH����es�����c���0�l���o���fPE��Q$��5�K�Y���y�[6FU]������v���u��J��g#�rp]�0��q���H��#3D�?g�k�9�mn(2��_vx���)FD�ӊ��%:�ҧ"��EsJ�'$�!�^3Af���h8M�u]�͂N�8o6�����C�V��U\ �|��nh��A����.���-@?]�����bĻ_��S�9s�݁D��T��ԅX0"@��p1�]2k6/����>���t�ؤ^��H�S�E\M[a~9����bUYx�i��v���,�h��`3e�ʣ�%��l����j�c��C���س�Et]�N ��x
Wa����l�\�����HE^�O}
EqRĨ4�1�@���/�Ol�|	x2��R�qK��1�#(�		1��-�>\E��3JmE����ӊ�6�37�p �����z�(~GŦ�A��pu�ܡ�00S͵�B-���'2ec������k�s�Ӡ�ΡHN���+�bj\"���$���ׅe�7�l��^�	a�+�Q���+)�$���Q��D�<�k��)b�?:9�F�=��yek�+6���7Jł��J����$|9h�_X�4���ݿ;��� DI@ ��J�����d�a2s�+���_u¼���V������h�
��2q^;�z��-S��P* uP���ㅕ�xd�Mc={3�w�zi�+�2�W����Wt�M��`��I�PU-b�%^���9�c�@=� ]���I �����r���9��v���(��+���~����x��j��
�u�GK���6?���Y����^���Y����Ѧ�#<k�_O��(u>L�L��׳N������D�^rP]���dw�<���M4��D�5:E�j_�#� �9t�a.�%�	�7�>�9���k=U�N|P�":�u5��Z�P>���3vzIx&��x�piP5�Z�|ӗ8��Ds6�$6��ZS�tU��$qSH�hD{D��+b�dYa�l�+!�[����Co� ��@T�FܬII=L�]n�T������;�����?~����)C�����rD��(xE%������󷡐���x�Ƣ�s��x�����s��:�{�2��%)�$��Q����B"7kĸg�\�?�� �k���w>X�����IXr��!�uR9���fP5��f�Ľ���Qn�l��ڡ"�w�S����h�����8r5/,�VQÍ16���A�E�Dၓ� -�id�u�B>�~	��C�IyEt�-9N�xE/�2m��~[͂�o����f}h.3GG$fɋsgm�/��^�T��#ybf�����X�	���3Z��>�)Q�>�CHNr��x��]�0���e����u��d��R<�kD�u�<+'UL���"iH!�'x6�P�?��SU���=配�fg�

Nv-嚭��_i�4[w�`��3������B��ջ�L,+��_���F{'j�^��gsޖ����H����$�4�2�P�[M_�%r��Մr	�9[)F/�J�D��W#�es�;�c����Y�;�;'�c�����t�j��H��R���^wQ����"k&W��.���w�Yx{�{�0��Qc艦z���9T��]C�*W �N:��FJ��R��t%��:�5��L�cGl����$��*C�_H�t3�j7!��6iG�g^�j�X%<������R?�y����`�:�v�s�J�	���ݲ��߸໘��{����tt���^t�
�"�~t�3D)<f}4�+˶21�]��&��Z�rW������qx����Xʨ б�()��zV`��!���B�����iͫ������U��wlU��?����˴�ẗ́���nS�<�lO��!ؖ���<^-E[�_�Q�ų�ʆHW��ަ:3M��!l0λ$���$�N���0�hV,וn��B.�	������ϳ�ǆ����5���Q�m�e}�x��Dk�
�����' ��+J�  [U��tqB�)��>�݆�b/�p���R����F��������t�v_�^� Rt9��ۙӑ6�����6��&<�O):JUpb��K��H��n_��L��q�jﵗZ@�&+3h���x�/�W�d�	,B�kQ�:�C�ͱT�}�r�J�G`�h�'��]�@��b�����6-����J�b�.����C�z�%Gc��Ch^���r��Ԩ�
�˻��-oB]+I���dD����|F_�C�iO��AӃh�����:���h~0�k(	��gH)<��h�����b7 ���\��G�P��"�.�h����B��8��E(���1I���a��w5L�k��xP)Ըn�̣�{���R=��07h���2h5����90Mh~�\���]#f����cj�\�}�6`W���gQ���3d�/7�I�3F�FG<�b��E7���ȫ=v��,^�]��u^��P��b?�X�Țz��"['|QO�*ale_��o$z��=��WD��0��5�ogQY�i��')�I�&�©&m	!qs��f�mvﰈZ5�M���T���Y9� �Ne���N���:�U��l��`V9A���v?]�K)t췖���u��#�ݻ(_�Ð���y��R�ų��wa��ۛgf���_c�b�~�)*_x�O�nZ��C��s���������;B;��W�F^�Ӊ�ve9}S1���|�L�8?����m���-m��: /�s-||�}����}�>~м���:��^�2�s��!��|k=�0�G�:	�П��s��Bu�b�9�b��r���D-�U���qCG ���V�@��)>0n�?y\7�M���=d
�H���qp[3(m����S�����@q2��*f��;�is��
�=�][L
9�T�m�n��>d���Iʯ�G I�pil�G��ׯވ\���C�YC{�D����'���������h���w��E�����2$�T��.��<$5g����-E��/hhd�~�F9� Pf���-�(�(�i~��TG`������#W� ��_B�mH���:NOs�<�G� �ܥc��J����p�RBL_���Z��ڿ��w���0M����m촁���t	��!��z}�!�{�Sp�K�?ۡ y���"��G1����eK�<���m��c�����u-R�q5ė���vo͓�n�(ѭU2kq֢�82n4~
���[O��K^O�evA!\G��j�z#̲{n�A�2��[���q��E��4�����ei�Y̥ԘP�'�{B�ߧk���h��e�2�(��*��c�g[x�����^����C���۪n���1m[l�g�����`����1�V�6?r�������ͻ��I<��	}j߰7f�Y�tH���R��I�i(�P�1���)?.+�cl�4	�X��q��1���~����V��e*,nAZ1�UD���0��&�f��B�è�)��\
$`�֘��.�%�;׷�w���2>�����?���Z��\�m��wK�kmW11<p�61v��	��2q���_��c���a�O:�`��O �sS%Ay>)�%���,�*E�p���/�K��D�ձ�"V��x��o,�h��byRI�T���Y��w��H�/d&�V'��-+�	%(:|��}��ׅ��ҵ�<	�����+���:7x3���x�$���6��'��FN��B�[7!�=0Bw\��G|���L��߷�(�E�P~�`��sooɄ-q����̢�^�롥�y��2�{��}�����k�"�]Wj �W8|hj���Hv'6��Mf�/�mm����eo�ƐDg�$�3�X��A�OF�U�l��>,�3|��:��co>��a���6�4Y�S�@`��<4Y\"���������7�G=�����]�D�[M�5�r�wN\V�W~��8%ޕ�,Gk������)D�"����t?�z0���5ڷ=�։���hL�.S�H�4:i�`�t� ��s;.�x,�4v!5���<�'4��mn�v��n1
���En�Z�,�9��\��ϯ���{��PfĒa�q����g��$��*���|ΚG�M3R�����(*�ƙ���d��b���֌0��a
�('�>�x�P�1[�T=e=Jf�J�(�ct�ض+�.��p78��?����ԏ���pj;VP������)���H���EPl����6t�6����N*�Vq��-�魉����/[-0���;rr)�5@(��!|�� ���c������2��Zz:�䮹��Ǵ�~��M��,�7H��e���>����`]Q̙{nl��6�Eǃ=&�PF}�;�s
&��V�`�New��G�\��Z�"��U��jMdc���D��xq�(����	2[��|��w�	��m��7��Gz��ZC᤬�j�YfX���ZY��u��.�iQ����ѐ5����I��;%�� 6n8��R�1��"h�k	��MT4�i ��9� ��������`�������^�hM�4���<�e�L��&�L_��xU�r��@�Zv[K�h����_����@|*��޲Q���u�*�+��󕘍0í=�vX��r6t���1ʡ����﷚�z4ll?�pb����]e��'&�#C�'�ͻGhw�m1�:1�$KȬc#������n=�n��V��x�6?�1`�o"7�e�jV����**�ٵ��:���k���@�g��䮲G�''jA�e(`�ǛK�U��h�←��p���y�U1\� !1�r�o#Q_��eT�N�w#�;R��|Y"��I���Қ6�p�&Ir*o�Aܱ#4���L�
���'�L
a~e��D�ڡ���"i4W�A��n�j�S 6����O����}��Z��)��rR�����b��kE���;������|�O��X8JiO\�i����w�>��a�e���ɳ�&�b��KB����P��)��݃ OAę�3x��Ō~� w�����.�2����}��;i�~Y�״����s�j9^���ż�*�l�M4$D:���K0�!A�M�,M@S��u�Ӛ�-!N�.���ܪ�w��)�>b.�N;�ȒJ���,��T��y�O��}�w98����0�B�����[ݾ���]Ϯ0���z�:Ml���_̬��kk��@���}I�g�FC��՗�L��Ac,GQ7��6%	ܵo"Q�""�6��J	nQo��������L��o�s�U^^a�s� L�E'���eRQ ��2퇳����>N��i.6�c�_� v�drN������D,�N�OU6F��'�~�k������	�<l�a-(�����!�O� ������D���@A��>l�,����I���S�X�b���z�w�8��QR���m��{������O���[�YxNs:Ż�ZȞ���� ��~X��)|�6�
���=m���:.����J4�W��.���$�y���-3M�6[�㍕̹�K���"���b�ԗP�4��,؍H�֮�����I��ӥ�9�4�2����T#�n�[U�G�Qy	��ޯ���Y@bL��I "��"�y_�cf��y��o���������Y��Mq��y�h�8J���~]��\��ʒ�s�C���&70%+���4L�+�)-��;�i� ������(n�"�h督��.�F�Y���5�˵��Hu�6mK��x��ۼ8+�'�������_#���8�맺s�(P�{�ؠ��q��6`�M�
>��9��C�[%�g�#��S����|�: 261� _"+����@�v�A��~���x|[ ���r(��]�kQ"~9RNm�/�����z�g���s|��!�\}�<�^���{����Ĭ�J�a����Rʸ՛��fH/��zB��Jvz�� �D�$�~�1�T�M��hJ��{ԦO�ޞ��`�x����(��Z�e2�[XX �~�?���v��������g�N�&לcaۚ7�Zăp`(4��]gS`�� ������p���t�p'��z90Eѩ��p��IşM0<����_��yqg&�$cܽ��/���NЃ�����#D���W�Y�|��{\	�NS���l%m!Z1��e�@�oL��y���t@c�5׽/�pXjE�<�G�I ��Y�>핚���­��v	�$�Amz��Y�y=����4��M����"h��3�yMk̃�J�1Z:3�O�h@�XU�xI'콁��W�����|�z���O=<�*��	6��_K�<j�?Z\r��4{
~�;���{x���/���39|*��e��*��1���j�/�Id��[���7�x�g�Tly�A��k9���H~4�&f�̙zC,��/���%��K�Ed���J�,f�@Y����ª��]����Zy��r4W#^�_��7-��[�[��Y�\&��M��l�?�M�BErӮ��J73�ʛ�[Z#�7�o3"Tl� ʫ�u��c~�<+�9􎡛 �w�0�Э��b�\P�O��B�Y�ʟ			��g�MS�ԏuV�K12�� �誇	5½@�7���<횋��VM���4�h��'5��#C:Cƌ�4@$�I��1�s\4�Q����BةR��&�},\1��j	R�����ln_��xhUN��c���^�?µe�H�H��$B�M�#�_3�F����OR�w��
� lO�,���rN���]�d��U��~A��q����2�3Mnj�j�{��|��a�f}�*y+[�*�9#ٴ��c��������)��l�ڡ���I�HM�;Ӡn����Kw ��sI|�
(��;��_���9%��jƏ�������:�77����|�,8��ؔ��&m�,)��p������-Q�r����	�������sL�0��D���x�v�����BՄpYۼ,!���uNxo㐂S����F�cµo�m�Z�&���4Ԃ����:ķ\��<�˚��m]�Lئ,Y�'���}:������y��X��d?���D�c-��c^�&nv��C��X[���:Sp��q���O��
�n��� �lܓ�D�*�62��Fy� �:����i���r��^b�kOw���,�$�s�a��4K9a����A�?}A}��ƺq�1i�)�$Bp���ߋ�����\�MK0!ۥ>@).��5ϵ�N��XP'��Z�u�e�|�$��fI�^v$C���#��f�}oՅ���In{nw&ܻE�}W]�}Ȥ2��֭枫S�D���)������ٝ��wes���G�I A�7z���U\��U/e����y8r2i,��O��#-,�>\H]�(�	�����v�&?�D����[29�Y�� >6THԎ['�d;t$��ߟ�/E3�W�k�a�pI�;�`f�>@�����й�
����/�hUH����"�θү�q�SڴƚA�H�<	5��Ϭ,(��;{n>H�~y����R_A� ��n��T�I�e��2@�D�֙�M�A�����8yG��5`	th����∪�pTW�/F��q�f�@��I����l��τ�H^�UOo�ɨy��� �!8����s6�n� �e>�+��d���Y4������֠��d����}��N�=liA)��ض Y�t�|*IXp3�W��U��$��?͍P+�1R���2-C����~��c�[Ti(���i�iT�rڈ�(T��gS�����bR�ß��������o�����X�ƥ�`�+{EʑPQô��[��a��B�PiN� ?���c�e��$U(���1�iљ��:}{nv!D�V�+l��&4	i�C�	t2^��Q�%��G�SW�)�h}?u����T>"5;��v��3C:�Z�L��R���m�F� � Ӻ�s��q��ƿ��I���6R+�mK��R����:���&|�n�]��+�2$��$�' �'�'�������-��$�=)�G����j� �L�
����t��$���Q���=������B�=; �9��	,��Mw���MԨKT}���a�ڻ�r����EI񳪳��2��� �u���kzCu�m@!XNf=�����Q�dR������E`I�ЊB�.D��3�d��q7��4Rm5�)k!�[����íB�w�u'�Ͼ�>��G��y���AS���ߧ-H�9����8*� �n���T[�9߸#XO�Lŏ���U�{���7z��-*��&:y
g"Q���7�CgO07�?쉠��*�d�ߵ�c��e�L5���]�㟒��.>���m����Յ�
l�P��@*]<�V/��o����|���#BԄ[�ƎWK<y��械*�N�/�,2O���Ļ���:�͞6��4�I��\
0P\T�Y��{a��˴w[sV�2$&�N��[hn��v_��7¿�"���X:��C��H�FLΖ�J92�Î�Q��[�z��R�ʿ�,b5�M��FP,��9�v�}>�g�Y��r`e�t���!�y�v=�S��v�jXlτX p$��O��0N���������@~�A6H7Z�	���+$F�oq���&��X0z;�<t)r#� ��U��5��x�I����E1�`e	��{���[���l��<5�{�6o�İ�=&��������!;d&�W�D baގ��D�τ:Q��|	��{0�vsG� �]�"�#o.s�_$A̘o�������91-O���O=u���Q� �%���9���m�?��j��\Xs���Ȣ����s�}4�j�Lb6��܉-�0^�O:%�x�����5+$�aBܪg���S�^Q|H�Y���%v]�ȡr@�����]��B��S�Vd�YZ/�mӬ�+'��L]�m�������0�
պ:Y���I���a���<���x|<j�Mc}ab�4�k�e�����0�8�ZW�	�^���(xfˏ�O:g�6r���߃{��[��-{nzu����I���(�y��X�A�x�zF���PvmCG(�}���+|{EBy��'����$z�]�~	Be\Pm��}��*�dk�$&]
� ���+���9���p�P�cy���w�E\�I��:�"V�Wn�o���;�	]N0�� v����T���n�^a��L6���B��� n��)�i�U �d�2ph)W��d�l���ĐKo�ĺk��yU���X��T�s�R�~��9�  p�Y���~a��x����E�
�����J"r>��,m"���R)Q��z�;�2��B^�Qp=x/��&��������j�k�ʺ��#ʺ�2�����!_��� �{--Y�a�(��hx��0�F�@~����c��j��n[�t�a��W���J7�2!�$@�i��8|�{��,�Ȁ!jW��M�'���D\�4�B��ϫ�!i�K��3Zy���9=TF��|k����R���2k�uڥ��.�c�IUI��Z$)�o�5 F�#���e��Z\C�{Wo)Z0Y��K��#�� A?����U!�ΰ��&��y��4�@��}ތ��p5�x"\"DJ�����&}��nt޲23���$��6�_=�F�8~Y�6�q_-�j^��D�i���aG�IJ�&a�>ܪ%�#�=4�IT�^>ڲ���C]^�e�(�i�t�,�(�R��;3����f����ND��j;�%-*��`m{�W��{��~��F�5&�3��$V��*Jn���0�a$Ѐ�C����P~E��������p�:���a{��j;C���N�3��#�������R�`�a�� �����GT�[��]�^ U��J.�����s7j6q����S��!O�-��'ȧ �_%\��Ed�����`A-�V	����$y'�E���`�E�=1�6�2Ԩ:I��uA���#�ϱ�Xb��H,h*zsN9�K��@!��<���h�����-��YS�%�0��g1#^�����{;� ԗ�N���C���@N���9�k��%�X!-CPmô��d�sM@�����
.FԊ3N]�i�L�L�]4H��^uI�L��D�
zo�7����e�i��Z9���Zl�F~��u<�a+R��J#����GD�Z��y(�+�]�0�S�3�M�b�%`,`�*��k2�H #0�g��1 n!���	�.rX��I�V��k�Z���a�SԎG�-N���$O��L�\�֌����?���q/����Dy���%=�_��Æ��#�ǘ���O�ۇ��Y�eT��XM�l���ыH�2I�a`�A��(>��p���O�P����д1u�/� ��t��G1o��~���h�ߐ��$� i�:��L�'���Q\�W�9��[�_}��n�bF��N�Ǭ͋ &��}VKi}����Zc9uPg�Ny��M�PP�Q'�<�2ӓn�(��q����t9C=A1Rya�Q^�"Ui|�,x��o�)���>�Jh�ư}`��f�ٽ}4
��}�����s&wlK���)�%.�DpH��ÓuEzLYT@Ym�b� c$h*|[�ؼY� ��0���~>O���,)JKQzgP˩ү#��XP8�#8i4o[L?��=D_ԱT8�pC�q	�8��9{���T��$�l��T�؛d��Zf��
�����)C��1��W�D�{!<�8��t����y�T��4��]X<ZDu�a�#�)3x�Q��� ���KcėFR�\oO�X��%nP��ԽD��Y�KÌ+���8�|N�	��Z�8ן+Z���&aX�t���w/��v�	����������/e����hWH��}�Dp�xv�/�ƕ� : ��1w�҂�w?$2l�HY���ev����.LR�nTF��*�X������u��|˺{}�'�����M~�Dv�Ρ��4�ٰY��.�X��}��S����p�C
m�3�h%Z���R��m �I_!�kփ��N��G���a��r1k��]�����<�&व��2����tT ���zr_�[`��6 �kuW���{��;z�5�_K�>-���iK��8���hh�������Q`�Hr/gT�M7o�Z��_q:��J�f/��_z.z(#�7���+$y6Ww��y�@>WȠ�����Py�x�u�T�6k#u�o��nm�r��I��|w��⢩�cѧY�KA�4�	�EP�MK{Q}.����Ղ��+�,q &��۫Ĩ)�7�ˀ>���6�K��Jۄ�!|T��� �����[T��aゐ����fL��*p��}�XYV��=�,:>đ�S��.5� �*�.���c���̯�"3I6�ִ�C�� }+����'!d����bY���ŕz1��+����u�D�Y�B�B��B���pIɵu
�\4w�uQJ��2$�>}?��X�-�B���͵��C��ˁݢL�m�D�pmĘ�x�ǥ0�����ް;J���9MTh�GI��%!�MD��%`��T��������Y	�Moc>ʆ�0�唄���^�	���VL1��6���`pq
u匲�,�;��t�?��g� �f	Y�FR���6�i�0G(:+iZr���xu2V�*x�߹Ȕ��2(z���?]��}��,���6�����v�0��������� Y�����R�~�劭B������X����%7I	���tl	�����]]��Q�K�,���+�=�!���O�C��O�gh���!��tdozQ���U�� �Y�2���y0X�&IHL�*�|�@(DVc��Ì�U�p���O}���V���hj�%R��=�K�xry�~ja4���<�[s���Ö{Ep���<2\����c/���]i��E85$q֨z|�����o쨧3�/��	g▧���c����d^J�,���*��EM/F�o�PuM�C^�t��4���ն�$�'�O&��b�-�3Rpz7	d��.:T�Tɯϒ,5��L6�`)�?4'Q����0(�;i��`�|�Z�9P����z�q���ze'i�po1�\�ͬ�&�2Lw��6 �[�a�����_t���tK����S;L�i͐<C�f��#4����Q��Q~�o��Q7��&*[�I���*t[�������G�^+0VY������U7)9�:�DC��tWj�l]��u�	��� �XHF��)q���]���(a�c�� ag�
r&�����\��>���N���c�6e�r-#�1���d�ҏiE��^���V%JAPb�Y|ڥG4�?tш��K�`�p�:��-�HWeeh&<�y���>��c�R[���s\�k���X>�����*�-g#�|�n� �3x������j齖~a OA���wq)e�5��yX(&v�����V��
��)�ɒ�s����i}c���bYnK8�PHx�%d�������)�6�^�
n$��;&�Z�!1�?�d���g�>�<~�v�������I����Ӹ� �T��O2)3L��}�a[�Y%���X������]:�ʥ��&�G1x�c�w��K��k'e��%���K�y�cs�_]�a����FԚ�>6�+�Fg�]n��!�ni��ǎ��sb5���ߴ�8�����:����ά�JC�l�g��R\)�3k�w�,�K&w����1����x��n7���.�[V ���$1�����v��e 7JZ���csr�B�#��_B�C�
{8 aF!:���pг��� -��ݲt�ͥGQ`���~),�4�&�������Q�ơv���j�@w'��7^� ��c���=��4����](�(&%�>|���|�(�/T[I�w�d"�Zܟϩ��!�����w����z�7F_���N'b6EǏ,�i�,��nr�8��'-}�~��o�zĈ�q��w_ F42�Q����)4���X���=m0�?����3O�-Yu������hvo��j�KG�O./)��]���5i��~ ^����FZ��-|n�rz�FJ�����1o��Qq<��X\Hf��.�f>T�pb
�Z��iV�߹)��P�ʱl(10'�F.�Kk?��yD��u���&�Y���Iz�����9b�I<lx�����ON�}���arF-��!fn�W�c�U� ��u"3��[CB���z���0�S֐}��L�[�V�M�/��p'���:
s��R	�]ף	��Z�b%g�_�U�>V�RY�5�a:�r�O춡g��:���<yF�fq���q\��4�7$�U���7ci�y�]�!�Ó=��;�U���:�Ĝdm`	��IO*�������nK!�
#د��
#0#8L��U\R��}�����9�J��!�<�O�>^��r���#�  �.-U�]�Ђ���eVB�0�"�)�x⹶� ����t$�Ajse�tV7�T�O������i���i*�%#6k:��7�>֮�%�{+�o��"�1�F���z��z��t3+�m�F: `;�ۧG����5vY�9�R���ˠ��ՃN-�HD����s�� ����_���m¹�Wmk�=6&M�~\-��mDV9BqH��݈��c\�C�8�p+�pu?!��^ƔB����p~L�IfH���HC9��T&Z�40� ����k�h��U}h��92�G�����g(�)�����C-���R�׌�i�|S��#�DY�q�=؋@�`U� �8U�v���`0�r��B�L�(��-!l�_����+���-(��$ؙ�����O�^�}�BH��Z�� ht?%1R)�ڙ�4Qo7�8琞
x�������[�}ᆞB˽T��M1�M�O�E�I��j�(�,P�e~�d�s
 ���u`��݆�<��g�N`�6�|�u��}V�䳵����|q=�+J��?����IF�:�� ˄C��1��	y΅�f�ƻ>�|S4�τ����M��B��K�q)~���q�hE��y��}��na��i�#/�0���k��/�3�NKˉyI�6��:�%o�����='�R�k�{@`c����	|�c>����r[��8a�1Ul��>��V.�,E��F�~�&n`d�>���ǿ#o��S4<Ӄc 2�AWB�����Wz�"���r��4����X��w�khL���"aC�l�+t�I��n�t3�ۼ^T97&d�F{DѮ50� k���x��E�ǯYt��BJ&��e�H˭����'��9=�u�y#ʎ͔�{-M�Xא��*�)�=	���[�Ho�*owdu��	6 ��K��F �8��6��W��a�q�����[FIg�*�,��)5�FXb�E ������v�I���1j�����cy<J+�R��I
�d�0��[�d���=�M�#�������#�˜QZ��t����";��"�{�Ӗ�`�}H���X���M���m���m��(!x����i��s�`r��t�=�@j̳��#�����P%���bF�́����;�e�/)r�UFѸ���s��?VpO�I@��|(a�CF�����g�����A��H�``�� �y�w_D]��Q���ԡA$d��JTi�uk�N�˧p�G������C�]�� J	-]O�{�$���<��1D(���uc��:�}Ɗ"����j���)p�|#a7��.&�C��u����7���]��e��U�4A�G3�#7���O	��3*����Bm�Sߜ���P�E�[l*�Q��m�g~��a�2I������gAi��J��[4d3y�2��� ��U�ᖣ2|�Y���'�pz����2w(�t�5\����o�B���R��f_��,<��b�YO��"�!������$�~����~�V�_�����¥l�V�A �Z[�uz�-�[� &WVQy\[��)@Ͳ�1؂@�e#ʽ��e�_ވO3GE��dr����CtF�G�E��3m�knO�{=k0��<��	L��h��8�hE�|6S�����m�0���?�x�m���ߊq�SqՍ3��6�>D�K���Q��$�ҵ���xrt �PvNKj��6�*ژB���;Gz-ڼ�-�]�hY8C�XAkV0�-7�G�� M	�2�z0��K#�.0��i�f�6� �$��>��s����
�
�6�� ��ݟ��{�O�M\���6D�A2#x�7.�|�ɡ��*n���;�Iٛp��ҋ,2O�e~�J��J�����-H�=�<m�Jy���}D2�i�OB�\��X+M�'jU��
2�$J�H�q@�o�Z:��fMU�[��-�_lF-�o��kCSl~M������6ʋ�I�����?$�
6�2��&Ȗ*�Z��@��̋�������ZH$�u�����a���е!''l
�ɺ���ċk ���&#�(��{�R[��T�zyeVYrt����i�\i6���cte��9�D�Y�:���(2��T*Q&|�;!1�m;ܩ�:�`��"�zMˉ!\��48�6}}���m�M�d���(�!w�7�6F�����6�_㖫�dj��N��)���G)���j��)+.��-�����>P5q<C�g8� }se��i�Uj��7P��������w�m�L�[R��^h�0��4.W5oF���4�W��s$*������в��b�*�ϒ�(8��Yq=��3�?��_�މ���;�+�[#�����6���j�8zx��t�]�L7W~��ZDzq���"�uj��$*j��v?�w�_�`	6�Id����.�r���B�Oii�/0��*�>����!�Ϲ�S��4��jq�]��<>G�4�5& ��P(*��F�zZ��><���INd�ej
�@�{2ғ�y-7쒕�8�FK��~�H�;��sm���QrI�����k�0� B~TQ���z��,�hvr�ool���]�_�f3��V��#�k�q:�� �NI�:F�.|�[�%�K�}� a���h"`���[뷮�R����"H#��]��+AzzF�m�/fs��/� ��ܳ���#�p欝�Dgw��+a�G�Ǳ6Œ'��~�v���\��<kaT������A����>�T�7����!p�P�y�3x��x�WS��0@�a�X%D��Ë�hP���]2y� J6�:g�� �[��a��^ӿ�2_��	��j]�~�U��w��F�l�P!.���ug�RLa�h�ȫ�w�W�$���N�+�19��tH4�n��-��+k��$�*2��(����*E�E��O�ڗLo4Chۄ��o:�k��z�R��)���&Ԯ0{c[���������~���M�	N�@��	ߣHc��ƚ��*�{l����]������ۊ^�T�K��F��u�0;�;歼E�㣗�~�=�=laj)[�Mjվ��3���A�2�{S^��f���i�X�G�㘶t֋O�jZ�*~��v*��*�%�n��������)X�9��g�e�^��C.~L��/ӻ���\�0D�����œ�n�	��lQt&�$[n��:g/�xR>K#!�?���j�X���Ƥ'Z� -U��Y��Eͻ��E�{j�Y��Z�
M�i�l�;���J���iag8;�����*|�NϺ��i1�>-e�
+�bB��ރ�/�4-y^�T1�0�l�'q7Q\W�C��;x�NHU!��X�	�_��%̂��mw�W���A�?�j��B�$��Z�G���K�H�H�-���,��~�-��O�Nk��df���3[��*Yω}�j�G��B/ٯg�΢a�;6v?���;#��!nI*�ǘŠ�U��1�ھ��`���E�eB����<U�����ng�^�&C]���J������:�M�ƿI�= ��t݄�껫FE�!���
@Ы=�c�xqAX��;�N��Zv�/Z�q�1MY���;%C?�oz�-伥�0��� c
����b�E���evY�G�B��e�n\ h�Q�� 7��Ő�z�_$s�-">[~j�h������@�A�z�r��0V�H��b�ӑ�*�P�#��U�Á}�`�w�a O��y{Y����P)jt!`��}?��ՔW�HRwϴ�`�F��u�T�F��4�^;���I�/Jɍ��-4�ҁ�-��j����ɘ�G�*�[	x;A�k� �x��Q��0��>H2��T]�����*�P�xC��/j'눪��ÛM 
M9��#A�'�D�y7;����u��\L��ǡ�MQ�����]φ�f,����J�B���N	�FSmY$rb���Ɂ/P���[Y.�;<Dϼ��Pʍ*�k�����.n[G��cD���dǂ�B]M��l���щ�؋����ji���ڕ+y-l���~ٰ���E�[t����E`�>���Y<���1ȂJ��C���J�-j�Oސ�Y��|IEo���ӑ��	�uI�8��O���JC�?��3�
�$j@m��|Rz���	/��(�L0�{[��E�员��Y8�KfnUb������ۥ���n&��K������	y��q.��n�R�}Ϯ�Q��xzzdwH�8Ά�`����O�q�p'�v?\M�bc<zdI����7'<�n�3��L*W,[3�>�$y�p��j�XԄw���t�����������xkDê�>�5�&jo��/4�I5�,�<`W�R �uIQw1i�.7F��/�������l���dr��8��+�P��pZ��WH���[���`w�J��:m�O�)�UG1��T��o6,��M�XA���3�N�$o�i�������rL���o��S �z����V.%tJ��+��/�sO3��+��<!)�#$vy��WԪx�cQ��߁�������W{V�9Z��<�&��u���#�l)��;���$t,�d�\������xc<Ě���]H8�P��x�E�1�9�3�n%�s�\z((��2".oG�G\zH#�f�n��O`�e�G��7��i��L�ld�N�D[ڱX����%��UCip�~ׯ�_��嫊ܖ��V�}���<�`��LP�8Ӛ��O���o�m%�9��S�	��vk8WTm�r���<$�AR��U��Bo�c^媹�bj���װ�Z�W�4A3��-bc1�������u�G)>�A���u�N��uM�<�jym�u���~o��ItQ�+3`�[s�v;�8Y�����\7����1��s��bA��t�������̺m�!����>|�B�����D9�<�P�DHs���tU�?[���2Ч�g��$�I�Jv(�Sܙ�z�+�
9*@��{T	h �9��+<�u��J�|�E�g�I�d|}nD��\)@�^���O�FT�#�+@m�蚺h@�ئ�1*IN^eZ��yq��T@��׋	B!��x|i�P�o�*�B�`2� ���D�+��Ԟ��A�::��|��=*;ʙ�pF��Uʑ.+��g��vB[��b1�W�ᇼs��ug�E�+�o�zA�~� ��0��Ih�*�Z���S�ԙ�߫J�0�_������w|�0'_Z�(�b}�^e���w(	}N.��X�e�;W�eњo�*F��8;�qΛ���I�JCf���׉G��p]r!�e.��Y�n�d�}��n=��8��A�_Ȥ���u�6��M��THr�U��Ha|��zl>|��d��K��5���v���Gqط���������4}���O��.��+!6o��M��V�]�e׆������sn3%dE�	i�E�!F�ꮫ�l�]�.m�q$t��ٻuw�P0��0%q�^^2�d���A��%�;fB� ����}l�H���"���U8��,�W�4��@�+�=t�<[�L�=û��d&�"Im��C�%l2s���ZC���[1?��=o@�tp<�[��jQH�QC���s�oK�h?����Nn�YQ~�{�;~y��¶I]��;��/@ꪳ+�ڠ%���+.w���V6s��$<+�ҵ� �L�1�Py�{!79��	�� x)�go3�h���T�nm9�ރ��׫'T�H��h ��6s6;{&`9�c��7>W�ճ��v;[��ث�q�T�Gn������Ҏ��TK�flڤ<.Ǻ��#:��½j=�'�>�����TC �oѦ�,��
�<~��GW�ڳ�joM����RߣYGl%�tQBк�:�=F)v��Y�`��,��-��6#������M&j��/XT�w��}�$��d����&ɾ!&Ñ�:z������45���HBu�݀�z���P~Bs#�F��hV�
���Cf��&ˣm���G�v��!�|
t
��41<2%ւأ�Vt�x73W�����pH��Q�W�y����>~���I�����x�hKP��E1��I�E	#.*�w�R�`�au0o����\ҝ�йΚ8�N�C�.?z#��M���;���O�ڢ���:��~F�<B��~VF�ۮ����q֯W-/��qn���67N�>���5oo�[�M WHe#���ؔ`���귏�-?D��,�G����d䢓��Ɩ�Ys@NH2��]���k�]��*����!'_�{/��brP�!���<�jJ������t�y�ԅ��A��NM�k��|�7��(0�N��[ݲk�O���5�Ō��%A���X�3��{�e���]�O�O�@!�5l��F6O���2�K+AMW[���y;o���J��ۄ������#Y���{F���sծ�������l�/9�v����`YM�(�j�ւ���1�+1x3�PT�x�B~�����!;��aIV`���G�xB��7�5ln��(�u�A�|k8NյY���eS&�郳8i��v�N�*X|,��Nmw��a.��VH�*
oo82�̵p流z���+()J���ً��S��d\�H`���^��2:�=)��t�\�%�lSiWƐ�O@Ȼ���ף���.7w`]}�����<����!�2�e�������r:E:�1��;r�m#@GM:��v�Lv4<��n9��/��m�Z�Y΄�Ců .(��Pln��.Њ�K�D�0�ƃ��AA�"&��U�'���B��R����GrI��;%��ɍ?�����"�E�\}��l���ok*+��6X�=���{\�P�Q9���^;����C�*�(�RHO����j�&�Ż��	�������T�������;�Ѱ*�1N������v��$'F�^�H�%�­gA��y����ikD�A��Tσ%M{rX.x6��l<z�i35�2F
���[�̖���X���-o��#��f�����u�]�Sn�P��P͙и��D�;@й��7:KI4�x���^6#�3}�5_$��g����xU��c���CXy��e�#B��a�g�P�'���2Te�B"}�+]P��Z�)����u!YN	J����a�����t���F��(��o��	WSd?�.ǫA hJ��ލ��XΩV�MR�D���'�h�2���WCP�W��ǽ�I����T�\�!	L
q'K�**A���-ս�J/�![���P�.F�1�������Eb���$�M�ѽ= F$���#����1�쒾��E;#���*h�2�k��|�|����⤈���*d��=�C~
{�r)�����'��RM(��ͪ~�g�᭝��!���P�G������yc��]�.SZ�a�� ����=��a�bp��v�=-8�J����-�9H��R�-,ۥ�?�=Gh��Q��:�15\Ã��%�td������\dM�$�$7�� n�߼E�>0FMM�ޤ�}%G4�py"�T�mym�l��
K��bPJ=��#�\���Am���qRz��>�(,��lrZ�-DOݿg����ˠ8`�YKP �LN(+t��$T�����*#�R�3>�Lc�����i�Ӷ��W{��m�)ʅ���C>�������p��|6� vI-h0�hl]7��VB�`��p�����\������=�΁��#7����H��C���[�)�4G��u�H�;N�R`NMX�04�e�Od;rd����F`Nt8e�fju����D��7���p�?$�W����'����IG��-��K�C�ɩ��Xą~�JBd)m�P5�hh�$"��Z�`�P����Z�9�1v��Zx��1^be��;�dپ�3?��p����������փ�s�Gqv-�"�yԄ�3�ɠL����&g���l�U[��(��J�LD�L�ʤֻw��{��4�
���S�?2�,�H�c���.R�֗'1����߀���m�y��{kE�ED�|	���k4�ɋnG°�e����<��[��|��VY$V.y��@��{�Ҫʑ�˴+mKڻ
��"4�9�YZ�ú𦴃�T�z|����7h.열���6�,Fx�'/
�p�x{�1A�Y��iC�rgc#á���R� 0�M랤�a��d�Dp�y�
>���q
�^���{�N:�Σ�c�GV^�w�lI��T�e����ͺ�����ڰ{��W�Mf�����3����s�GiG����S�V�-\�Q�$�#I�)S�[a�/D�#��M�e����[�����C� �/����q�ȫ�8�ڐA���D�%�H<O�M�+2�t������c։7���S�# ��e�����mN�4���#�XJ���c|(=ض�3	 T���!әS�K !������.��C��1W��������ô$�>c��NDۙ:���?���U$�ך� ����U�=�|6C��q�8�vX��zQ�Y�HjD�Ə�^d�GiV�Y��ށ[�?�[�c��B�#��#2C��@�o�țBL*մjv�q��1�����pNB���=9�҄M��(xQ�Ձ����ל1����?���d��]�l��6��a7зzJdS!�Hs&ѭ(� ;�8�ag��>��5��V��x�R2���PQ�ԧיA]���uB�ieo����`<0U��i�[d�Ѡh�N]�N�<J/�:N+q�)@)��!'��pč#�I���<%�̤�\��1�4�;ڰr��9���p.fSĲn|��j|N�4��G�����h�Ri]T��@�Q�ܷ�v^[���[�)��_��+�P��յhJ�n�Eii>X*��V�5[ߨ�t7��!H��ٶ�y��H���q��%����߹pz7~`�G�4MҬ��j��"�g�O�'�gt����j�b�4�ՆtRu< �g�,�,��'�++��<w���0�z�Oڌ�z�@7aqX����� Ժ�8�W�۬�#�?���a�����&O�*�􅷶����`�
�X�q�I�8�����SA�^��<��T�����!��n��?t��,�8�g}�b[��m@7 tzV�ڲ���֣X�o0����*	��q9b0ϝ'�%�(��]r:�=Ah��� q�Xa��{������X�䩛�g�8Y\�9������j;#��h�?7��	��>,��S��>~Q$,oo;M(�~��W��hs�UЫE6�e��
��م�#^�lщ��.G�߃1܁JXy[W�����Ffw��S0�5"�k�G����<��jҿX"1l,�":ڱ�ná�D���3���t���<�f��u�֊��t����c��0��9^#bo�j·ꍟD4���1���y-Q��v��� �!zZP�j��<���i,�`�z�[�#�z��А���x�LFM�ץh
���0�<N+��YKXХ�Vk���!GPo>AV�K��!�\���VE�uY�i�h&ڋQ"�Ӹk:��&��O���E[�D�	5ˌ?`>X�a�EW��*���<bc�:2��I��I���T�ElI��������6p?R���Ge�ȺRˀ��ԗ�ة=iܰ �|�c�=�]�Fu��P��F2&as���m�r����%f�X?$
�J�vA�q�����dO�M_��p�pc���l��^oc�" �gj��+W�"rF�>�lo��� �?�9l^�g�T3렬X OY��i>A�e&��.�$�d�.�3(������H��"�ؾ#����!�5oĄF��@h���@VR}u<:'���u�i�Y�ԣ���kY��~b�$���Q���2л�:�� ���Ơre��x��a
�ɺ��$��s�����r��
Ã�����������|}�o�R���ݪ� ,"�qTw��D?Q�����C��Į4T^ߗ�D>�&|�������!�(҆L���ʍ���x��0Y�r�w��DT�n�E�ls��a���9ִz���n}�R1���j�������4�3�'���Ź'�H�TR4W�H��"⋥�d� �;�?���;��w�&h��nC:j,����-%oBѳ��Mо�c�JfG����#hm���t�x�}]��W�I�a�MA\�����p�2`��j6PO�h�A�rU&�:Q��k���,z�:ı�c���4B�'���Ϥ��@���Q�n��5x�;<�F�e�q��{��튉,���5�c$b&���$�=�2�&�EF������kM���UD���\޴B
�����>Uj�)+j�>1;axID��_ڽsSB�?ܕ��I�FN4H'���`���m�FH�:z�{}�<��<�|��qX<JX���1q.ol���4; ����������83�?�,�ѫ������i����J% x@��
��ʿ�0�	����j�d$Z��J�bjb�x"$� ���Mxj�������vŎ��_� B�I�_���`&b��{s$�{����7�KM�"퍽��	 b�Лj�����Y�d-��k��?�T�'i��8lS)5�$��i<����09�&zx�DweV\UD���.T�?NfA]<]}߅��� �p�P�a���ǯ�{�Ѷi�Y�2�w1�'��e��2��k��⇋��k��H!@���(}��k<:�-u��u9EaA�9�>[_K�����F(���vЎ�wg����&�*O�8J�#�d#�w�<��o���-�.qEK���(����L�,�"�Ѻ'�̰���I���t'U�x���$��뎳�6��y�l]�FҘT
�x�f`R2�Rr�M�����<6�q���!��:��3�϶{�p8/=b|} Y�y���q�E�>�)1o9��A�K�/�K3,��j�{Բy#�ww/|Z�����S��l�(��&)q�C ) ��`�<�t��,0L�ƨEȊM
�g�zc��+�Ó�I�y�Y82GVew�1�׷����
X�o�����m�f��鉞�Ye����e�P6���%T�����BZ&l2��D�BS��� Y�y�Wy���x�Gއ/IGd�z�%�Z4 �@����g֋7>����8���+��� _O�ͥ��x�"�j�")�5m�oۼSS���Q�Q��dQ���I�� ��2��{� o���'A�c�U��8)�v��) E	�-���jz���3z��c�:e��a�0
A�=�.�^:����r�ޯ�'�J���񚃏��KQ0�8!�M�@E���<F��������4.ۢ�T�C��wDv�6
7/,�7��ra(b��>32��!q�����ٛ����f�S� 25лH�!��˞����ykx����1ܸ��(�P1F/O���18{�/�D�G����vj:Vɵ��!$�O]�r��V)>�+)��zFk��$�@ru�2�^&� U����mjr���噓�,�<	ѥПs#�x��'L�@Ҟ^�.5�`�9 yA�B6	�&9<nЩ,}X����z�&��C����?K���D�O�^I#Z��mP��Ru3"�R�v���F�^^�W2�Y1�hx/����$Nc~[�!��	���q�����(ڹz/y��o\0I�s������^���W���%8�H�N�t�9���1��0�[ķ��B|̞��h=����4w`�R���Y�O�w`��|.;eK�Z�Z��
�>BDڤ�l���5'x�j�IՕ@Ý���As����*=kq>(������)�K>�Tϋ�L�߿j���H�Z1��|F�],���R!;��_E��hHoD\&��x{�'"�����l%��z�5��R�w�� ��Zd���,�o1�ĉO�{���+k*(GAVv ��
GC�x�詫���3�����-ޓ� �^��M_�8f͟�Hy�0p���e?ݗ��z�J���.��{e�r�C���r�4xCj~7���@&`���9�^�|�icL�
|n�4S�𒥽HVH�)�P��`��1����Bu9��>��]L]�D��L{7�֟:Z����a>�iݬ:��'�9s_��Ǎ2�Yu�_�7e$
]U��ҁ��6� �M��h��3��1��ï�q5Lm�����#Ϋf���κ�݊�	Y��l��o(Չo,��:Mq6ᧇЏ&.*K� �����-��a��5>(%{x���5���F�oD<�?�ĩ%���!�3��,KG|{�2=ݢ�8���$��!�r)$��w��m�ݲ�V��n��Q7F�Q�cU�Q7+���1;��ތg��Vݺ8}��%!<���P�D���0H�l���R�9B�g>4\�u����{Z�¸z>�/`�M�&M�ce!I�x��>�f�T6���7��<��R؟ﺳu�.�yi���jii>���'��~-���Vy�m��vQ��^'�x��&�j��p4��k&H��y9�B��I˝|Q^�w�Ϝ�U�&;{1L��n�������g.K��B:��qY����ȋ�K��x�+�w�{�FyH"]��+Ĝ��i�ا/F/7U�j�&����`;��Z��6�҄�rA���d{�_�9� ��a,��^�,���Z����(m	��>����a�d��.���pk1�[FM8T��1]��%heHn6��)%������C�^�� ��8�1u�6��@��/2�$'3�%�!m�����Ƅ�(��}�,���VL�X�$�x�|���ke��J=��	,P}�s`�L=��.��Ky�l!��<��,v}3����[��k'ܐ�}x���Bs;C5Q��/z�'z�#�%A4�b[!xDA."潊���8RF���C�t�����
�^lT�n�����Z�y�	���Ț���+HN����O����g�H�ߗ�YbB�F6<Μ��1�^LXv��^��$sk17a@Ś���.����I�C�o^�j��=�(�d���#[���8�OH�=��jzH�[����j�����u���Te/�?8n�=Wŕ�E).��9l�ff��gm5�%��lF��� :\#W�ʧ)n}�X��S�5 D4��'�c��))f6�=~Ĕb�_�'�|f��'��aVX+����~�f����W�Nں8U	B���h�"����͹��r<���|jE���8�^�k�γ��h4:E�3Q@�J�� {�g���Q-�Vr~-�׃ �7l�շf�}�Y���������tY�cPD�K�V4٦�&M1�ַ�L��	r���sĖ�.����{��B�ve�&��nY�|?�l!�Gl�#b6�k�EW�(Ee��W�لj9~���Z�/v>-�����3�@��pN��2�����1�E�) ���V0$Y���|;�3�Xu�T�����}�hLLҦ��4��9j�`6�m��:ڷ(�W9es��f���C����S�@)jl��&DEK{2�ћW�+m�f3
�)�S�|-�$�W���)��_C��Yz�D�8���C�k��
�m�R����a��p�agpC<��/t�"��RWo�?�DxXm�T�3#"��Q��U��RF�l�_67��Mc�{����/��(�-K��D����(E�H�z��/��{��(���v!9�?��n�Ƙ|�|lVr��t|޲�RP�,g}�2�p�F/h��긹���0�Qk��v��7>��B��Lr��#1sC1y"��x�I*�|��_��/�$��eC�".ls���)�b�R�4�T�u�@ b���#J�� L�9/t&�_�\�0��NX��;'�����L��c\'e�K���F(��Gt"���r��u!h��i\�a\����F����y�uп1?8�&��@��֔s�)Xc٬��/ث_ل0�X��K� C8o�Uv�u��1���K���@m�7��A�a��K���n)��2#���Q]�Z+k�3�GA��*	z���^+�▧��ls��D�T�%T����w\�7t7�7(3	��9�)���~�*�t/��*�g�W�j���涔U��׳�廩���׸s��lr���,H��PN &������7�7��$�a�8_{�ZP|xsٕ����#��#�l��jP
eQ��{�A�em��`�|��gۙi��#܍g��I՗%�{�����[��w��I�ٛ�(=yG�'�o��\ɯ�g� G���s�za.�r|s�YI��Q��_����¨��f��u��=��=_рl7���+��9	RD����.Z�CB��S���$�J�	�?K�u����ă4Vǐ+����\�����4�����R�{�mTk�m��3oO���IWb2����=PN���*�.[��鱕I��"z��]+l��.Tn���ht�1�Ŧ<���Ű�*�V%��U<v�x`��j2�Q�����yR���E��F$kJ��x�c�����+�1�I^jδ��%a��!�<f��؅���㞞	�W1 ��꧐l�7���h��|L���'yk����hk
m�������xg;�3�2-�O�A��9 �(|��P[�!����|g�� �d�T|y��Gl/=���'2�����g�4l;�O��.H&h����r�9y/����T�~�����}�[ޤ$���(a%N����ꈠT=׺J���M!4��C�*&�ulq�����~�2��w^����e-%�U�:�0�Q�_6�g�"+��Xn��ʢ���ǀԙ3 ��o��l)I<�6���dB	.��l��J��0%^�̀���f�6l0��'�iRی����6/۸��S��]R�\�c���w�yگ�u(z*��Cy���ĵ�Ww*��N���&VQ����Ww��<������y!X$>���H,�^�1����h�.��pT�ǈW���kh���&J|ñ�c�[�<WHH._
z�h	4�o�_%��MIN��8���e���;��S�x�zl0�e��m��k�$���W�?��.���U��V�e<�����t��h��x��z^�r����D?��K���� ���5
����zsF<7Io��#G�y�`#Ad�й��³��!�T�V�Ck��/v7|�f��e����3�?��1m��˴�D��`g�ި���B����1/򋳫�`"�9��w��9�~%ҟt���:q�N{�D�
h����w�C�3#�\O�.5�{��9��%X폼Ք������ڲ��G�6�\2��ش�k6.�.�T<������W�(��T�#]�����m�eN�4>`0u�Ʊ6
wVSx{�kM+�w��S�開v7f3ޛ{�MD>��Y���u���q��VpFO���scͳ_�t������O}JٹR�'Y��١�燸dr�֒	]S��}�1s1�3&�����~�,廬�l�������#�΍oV*���������� �8�m�xb��A��} x��߶���]���*��
l����|�z����Z\n�\��tO�x���+/1r�����5R^+��N��������	�[��;;0��3������	���[�ܚ�j���;�:��OgH|�z�����T�T�O�O�1ey� 5 �Ͼ^���n�#Βn&{t57a�ƙ�����:bʹF� ��o�I+�d`��is���E�D�cY�i�vs��@�����r-��JH�$9�s����/��|��� �M�Il6���+ߝ�%i�����'�i�i}G��#���␒U�9j���_p��h p�Gb���u�-��0�����Q��A�W�
j�:Ok�N��1�M���[뜅�\x��L�&��$'v}�V�*$��X?<YKXp�GM~��X��A�(/��8���Fo6G8Ǐbh�^$�3�@�p���l�Y��@
�UQ?�aE}�����u�N��������	�(e��4!V#r����-�n�	GD���G
щ���������vK���3�bP�TiM(p���'�{ڵ�ܪ�xm�{~�V����ܥ�'�����I!�I�S�ႆ ˎ�Q�'O@��;��f�l�BS|Bv��W��[�SHPyĿ�=���pd�+���P�GV�7�=��Ѫ~>���Xi1�+ye��H�\=�^�ɷX���FQ��H�Sn���FC�tWJ�㟺�.��p�[eo��u����m/��8�z�Q=��|�13y�����.e��E�_W5UI�[��$���o��Sʘ
6��mlG�����u�{P�ap��g�1�ERJ��Ⱥ"�?���/��d%��:� "�m��d�P���|�7���S�=qJ|َ���Y�o�P�����2��4^>��v�0�Y��g�($�8��:[g$&�PRV�Z��Kʁ^J:��>�̏$��3�Ni��HMo'������u|"ڌ���NTŻy�O��#��n��`c�z��sN�G@JK�y;D�#,�X� o?��d���T���
gOS��ܶV&6��GK�d��Ȼ��GlĢ�%���{ef��h�=�U��껓���2nRt�)������$A����e)B�'�h�a�[Tx��`���_Y�[64�����ύ��)�&�N����>ZǇ�_A▖���=lyc`��4D������Q<U�{N��t�T�Hͅg	�q��c����+��-��$m*Rr ������������|��x�+��{��70n&�SM���R�����ԍwɟ¥-�Uz�.0;�h�9z��V(U
C4���⤜�^=��g*i��U�Y��,ʓ�h�r�ɖ=NKR3���\c�F/Z�T}\1��;���}޹��0�0h�NO�����FǧF���<@\�c&,Eiŷ=#{���q�ifHF
��;i�\�T#)�Iž�?��n	�p��c�bv�>��Z�y惺�i��_b�(%#�Ʒ1Y�xS���fG����⣍�9�{�X|蛈G�YCH�[p���-L��R[�0�����Pes��uZ���y*�~76�1@�� 86�$ؔOe����c򾩰/0�=�HR|�Ks��(:�4<����)_?����MN��~7 yq����'7��9��h@w�X��h;{W	����tI?��v�W����n�.�6�u��Ykk<Ï��'lI<�:� �ގ���׏6Qr��v�g�c�kð�nn9Si� ؼ���:Z#r����%{��q���<8��)�������ա�4���͌������JXV!�UX���{�b�t�FT�ϴ��N'����1����[5`T3H��+j9�)�6#�4�BOO̏,��+�w�\�1��S�(*�Љ8�5$��)z2�{/��z�u�ry���
���ߕ�oܣAw�0l]���k���"J6�hN ,4^�R<9ӓ9�*�~K65��qA�gG���@��5��n�g�
,�QC��h��=[�ex-�r:�f�R�]���Af�*��~
������6���1�Ά#�<�W�F7?�|U���]�Z����������"؁(<]�I����]4���١�x��jܩ���þ����C؆_�}zP��H�6�?�ףP�Z�1�И��4!��=�X�9w]<->���!�mZ/�*�-H4�Z�s}��Ye0�����85���>�4�Uӏ��1���%"9+�k�g���Az�]B�g��L �����N�-"�ii��0�� ��ǄS%ˤ��:Z�v��y�B)�a�ù�Kݳ6^��49tg6��ӹ./Y�4��n;{�f�"q6�T�P��<7�ް�rreT���e4r��b�lzɣ�9Q��ةبrw���R��3�`Waw��b�����
s����sb���C��]�x\7�B�ߏhT�����V}m���\�gX9���'�?��r�e�x��@!�O��#�7��<Q��>�D�?��gEr�	����~��,|�[j3��Pi�C=����r�����ӊ^�U�8����O�u�&Q���-��r8�q~�lt�?�7�qA$y�E,
 �s�#�$7�(��sЇ(�૚󒒫��pU(��������2Qe�d,*PtI�*Yp~î\ �y�+ �����S ��q��Q���Lv�3��f\�/F5T �υ�9u��ܻ�J�r�|� ����n���CE�h�mC�S��-o��R�x�'��8�2���m��%����r~7d�r�Y��Z�X`,n�Q�S~m�t�sr�>NG�`<)H
���]�D�u'��S�*>�<ˌf-��n�Þ��o�F��b�։��Y�G�K2E\�Թ ���Y�C{+��}�D�ߧ]H%��Q0I�l���p�6�<I�K��8կ�)���$�$����:B
��Q|�0�,����T�aCn*�N�����tY��(�.}) ����:����k��,��q�$�1��r.ގ��@�z���p{�����"��g�^(z���y^Ձj�j��,�q��%hI&�^F:���ʰw|�O3Zn噘`,?��t�8�*UFRߌ��U����ԩg�9�ު�XWO��T����Ɯ_0��x�W��vV&��%�S.�9�u�e���ʾ�OC��[wE�*�L�9����Z{�È;�p2�d�`�}D��8J��\T�!#z&%���#��P�n~���bN��	�o9� S�^K�����ԙ<rE�o������jk�x|͜��J�su�]b]`�p��#N;������l���w����r����Qc�.��&'�l�H�](ʙ�s�N� C$�OC䞺���l�֣Sh����-�zDW� �Hf�(�t���)��C�Wy�7n%��z?Nj8o?�e�6Vc�9��2�!�T�����P�m��b�x��wj�A��R;�M4xiC)�l/\do%�j�н�
��V����f �+*���y�q��-�.�w5'����2���ޢ�]�W�������;6qw���m�}� ��j@�&�!��v������+U�\��g'��]g9����R��K�'Wj�������R�+���"�x�[�oa��f�MF�<��j<��?���SY���b�|O�0��Έ��"������ڐGk�\�E�#�fZ�:@���ߔL��ǩ�LJ�,��#��kyF�%"U��C�4Ɉ'��(�b��Y���~o #�\�W>�n�ގ���̏���{�8,|U��,���T�`͏��P.�S�����\�Wel�Q������mpbk��eƯ��� �H )3#�S�LΧ��V�|����\��m���:��]��@�ɶ��ÿDȿX-�z���Ą��/wB\�h��a�yD$S���])m�V����D�Ģ��k���6zm\e��d�Et�VO�7���%��2F��l-�WJ�Q(��4��k��֔b.�FT�00\5WB�>x�{�/�x>�T4t�W��Z8h��\\%Rn�] \�ޕ�e�,�p߶���ʂ\��^�Br��!U�����&�؂
�z��:z�j ������ݎ�ё���>K���N����p��K��������8T
ڟ*�~@��t3��y����-��W����%u��ه�^�� �}�a�{l�#v̩�S�G�
\�_��H�Q  �Uqu���O��FvЛCZ���}��-��w}�3N2��`@�z(�gr����r�y�ꢔ#NL3�z~���0����'mr*�L����`\��'��X��(8qYC��F���'�k����� e�{ψ*�c���4E�)_�(�����s8��n��J������g���VH���X�[%�VS��;�CG�ly�"�`t��:��x��,P��O���h�-{��C�@x=��L�A�3;����Oi���!:o�M�Cz� ����ϼ`��ע� ����]s;k�BY����1aK	�P�_��}:�-���'̈́S��dBb	�*1�є���D�`� A�Q����E44��8
��'Y�<�m*���U�S�*�$�}̾�(�̤�X���z5A��C��g�%m��0���v
eFw �Ѱ��a4f�I��5��W@y��bCi�A�v�{��T^�Dٯo�].���ބP��9���mUQ��F,��
���G�d;˘gT�U����q�z�ߋO��3��
��QkZ���cP솙{��h�fj���`��N���b�,q"34�t�*�㩋����G�;l�C$6����<P.�]l�����{�0��lS�S�me����dv����o� i�ҽ����+�K�d���Z�� �:;d��TQ�-��N�cS�0Q�a �������.�ݐ�[_�S���jy�@]ؚ�}2PO*���]��X���g��r���J7�-S��9Yg:>����ơ���$mߡ�l�k�{��V���8>YK�:>h���J��5�-����C�4���~�iF�
��]����䧿��^QԴ���<����$$7����,sw&���a�8��j�*�E�kƉ5(�����������[����G�|�}'���-_��U�ܤ��8�m�m^�����}�7�ө���?�>6 J��m ��hlD��x_0�޵�͐J�u�>[au��Ȉ��a�"�<��m>aAE��WN$�0��?���xx�R�.�
3i(bb��}�����߇�Ph���v�c�"���t����BZG��Tї�nZ�h�	X
s�!�
Օ���C�%<QS��!�E�tk���/�J�"а�D\[��v�o"���o�7�V=����=-����\)(h��­��[���3���ak�ᠨ\<1�������u�F��7���<�V�/ρ~
�����O�jq��f��v'N�SJ$�7!&4�j�oR@��dآ�۹U<t9��\�A�`_��ұ+ �'���tk�=�;��U$��;�H1�3�UE�#fP���(�Ī�%�Kk"6�]�NZ9��i܅�<]c��i�&~��(܂�QlW6�f��F&mv�6��]1�N@��Ae����wL\���GV.�Dw�YOӠ(��R��&���N1g2˲Ǩi�ݔ������$��f�&��ݼ- Ɖވ�֏��Eo�+�6�}�2:Q�wS-l`3�1�J
�59/�EDh;��D���=|�a�B�=��8veOI�=F�9e��ǌ��܂!�{�MZ�a�t��������4�SR�K��c�4�4;�ǸVYW���d�Wm���p�����/��".���-C(S��V'h�Ṡ�'�)e�L%G�8\������Ǳ�߬D\E+�H�D�$�2S�<B��Zq�Au��E��VS=t���T���
�u�����L�<�ǵ��'G�S�&pUz�:��T�_�~ݟ�l���4��A@Z�۴9B�G"J �.B��M���۳�\P��M ai����s�{(n�%B�J'Y*gJ��k�8?Q�|���i�d���/Օ~Y��u�b�[Gf����N����=��pk�L�:Cr+�I�m�����V���r)ޙ�������b:^����B�u)�A� ��d��j�!����-a�˧ط\�o�æoF�������0yX�Wϙ�TF��
��@������1D�Ȯ2�X@�A��:9�:�Q7�`�����Z��FBXُq����?��%>���3J_e���G�2I=�T;�X/^s�a��억�JE�7�V	DF���.Rk�� }���Š�y�b��c�� ܉�{t��x�( ������j�'����ć�	�=c�c��i�5�צ��I����8Η��B��3fa7%Q��[�0�<��3+x��;\u;�
H
ϪW��h����@�r��F�$��bO|�e�^xu�ϋ�l 2��6V��Q�E�S�^S��?r�:�ݕ��4����!��=�lFS �r1\b��<�D)v�AN*y���=�c���;9�כco���Na�;��xA t�R!���9�^ݻ��
�m)�[�2�V���'J��\Z-��=����^f�<>��I*u��T�K"��5|�w��� � �E��=G�QZ�P�{�UF,o��?,�����l��9��x�^3,��G0�,�xVN//���ܲ��N�1V�"t~��H�ȯӌl/�t8�0�3� ��Bڞ����{�O�N�����*k�ŇB��ր�c�L@�ʍ���Q�z��	�x__l�}��H
���HG��x�!���& �GzϳRg��:���m-~��g��w>�/d�U�)�t{3U�:��t8�e�"��Y�l/ȻL���Bc��D��_�=É�~$�I��h3��)���Dԉ��m��p�ktF��\'�s�X�� �o �t>���؀�� 'ټ��Z�ڜ�`��j�������W���pcK͒��D��@m�������8\��^X���L��0M[�W3|v�o�M�Z�kMس�Ҍ��8K3�4�3�$�1���� ��7bL�In0�y�u��l��!�r�����<?�8��TQ���t�m�d���mu�"��]�PYr_�I�Þ���V���\H8���"�$53u)[�6�:��qB� �9��g����M�E:d��Ĕ�;�~��9�^蔏�W�]����KgV���P�q��dT)��.�u[���%�!�Of1-����i�3#S�`����R°Nf~�6�9�T$$���N�wP���"������@��#AXK�*������H'��w[���Kf,�C	>d�0fT����v��:�6B���Ĩ�.!�n�8�z��cc���vl� �D�零*��[�9�q��~(l�ߠ}`Qȵ��M�������r�%b�RT�m�5�;9ą�W�TPW�O�]Y�_����_�E�>w� E�h!g�1/�b�ܮ�a��R�7���O��{�:[���n$/�4���d��~�Iw5�Ƶ>❹�%C2E���:���N�vҊ�=�m�'f��j~��z����~Е,[�ޘ��6F:�}5r���J�[�xnu�@���T$/�z�Ɉ������m��bZ���еWM�۪�ȥH6����|/$z���[��\�ʣ��`�0 `��'M�h���τ+�7\���yfR歇;52\�\z��@�Ė�����{���`pŎ;��v("^�gd��r-?E���+ln���R�1�&�H�	��/MѨ9y�g�11���>r�b��k͗��ec�<���caV`9<�s�%KE�Ɖ>�×�؂}�1dIި~EXhz�zP�����.��*�,ƙ�N�C�r���L���Qt�=�3=0[kx���f��Y�3E9q# �kW����5#x��W�Z̯�'B,�i��)���E���t�(gl�`��!p���}�5����)iF-��u�0�8RqcEe�~��xv�Xrgٙ���bg�P��K�\Sn{��|��&��)&ɚ�iզ�v�o��؊�o�-��iÕ�/}��K?pQ�{tI�3���\LQ�&OP~	C ��y�KDڐr�:p�WM�6W-ŀ5�J��n
n��e~E�V�g��R�Ө��ʔӇm	�b�����t�ڳ��(n��t�@�w�Jt������I��H5���q�lVڍ�u��:fϏB}k��O^�LO�q�/u]X`�8�|ܘ��+ʕ�g����C����ӑ2\�q:ݰn��<��fA��Ф:��A�"l��\^�P�ʧ�!�
��2e�����"�賬�a���G����0�YiJ�����n,xۺ�w�?�%햨�� �
gs٨��*�s���M��U�Գ���̇_�7q�+$���
�$���*(Y�?L�k��ߛ{y�h���%���&�ֳ��i�
X7�0��w�B�8�������䈰��Zj�eK5�9��{�k�oi�*5���W�-���o��u�4��Xn�\���S�E�hS���[5Zx�!1O���dh��Y��~o�<������QB���OmK ���4v�Y �`�^>^&�\@2F�)�stPs�܊���@�� 	���*==��
�u"�x؋Ѕ���/���D
����h�9>�` �G!f�V�V�gC ^'Hk1��6�ѐ��@�0�)U�R����9�6�,��TG�m�hUal$�Jf��w���:�[�j�ƚ�`#;��+�k|Dy�r
FΏ�v{��+ٌk���z��Tyf�WѪ�P��}��+V�Hm��[c��EKi�T����r �}L������[���y�b&]g?3Cj.�B����?ݤ�\&��0y������D��/���,�ܒ{����n�\�Ӗ-���ds�oOTl4[tw������R��%�Zw�D���u����K��U$�@�K�"6�@��Ѫ�xɉ���,�y�N NK�����C��B�Sq���t�͈��;��4�`��RF�i_���ۍB��h��ǸӮ��6���O�g<�7�� eu���M�s�(�/���y�����0v؂�Q4�b�=!�L�)�!�R�&�UX��)��V\�Ć��+�R֐���G{��CX��!����(��GuAR�a�K�`�]��n.�����G�\�~�+>�y�5��{�cb2���3^_�N��{>�#*��My������F�9��F�H�#�!��4e5Z@���J۫��O��[����굈݊����(r��L�*��E�-p>��>�u�A��r���]Hs��Z�˜�m]�(�XU�cS���Hr+nQc�@��V`x\�����[��^?P���&'��5T�v��%Y�m�Bќ2N&\�Vt ��8첔C���x	�"��j{e-�P{!���/C�a/�k:��%[���*��r�T }�:��+B�ݻp/�2�٤�cG	���^�v�IO����d��=]=�&ԃ@ZR���=��]�a#��ȥ�h���v;D4��&[H�W��tqo��0�kC�%�yY���a�SLf=������¼�a��0���9�r 2�,��AT���S���￲T¬Jm��!ۣ���4�&�f�`Q��{�;�l��HQm^πT��ן���.N�6e�%�@={���#)h�����D��s՛�w���z���ټ�z�R��Oj�E�!�:�)���ɞ#BPW;���|���>x�����*2Y���G�y�������G�~@�߆ʿ��'�¾@Zr^��1*Vz�n�2�h��9vM+�^[�E�E����?���w}`2<%���F�A��>��hO��(=o��}�_"��}%S�!�dR�t�mи��tf?�����nqw��}��E`ު���rK,�13H���ĸlVsf1�*�z�!��M���I��)�b�?�P�M�,�� ����@�X��E��Â�l��U�,��T����گ���v�������m�	Ͽ�`7�r@��nܰ":/P���$�=�C)#��*��������tm�w��U;Òd�^k%����"��HQu�;��-\~���������J�r�e�Hu2Y�%�XH?{yܾFT\Yچ�"n����3�do�J���Q��4�K����0�6�ݗ6N!�^t�6�^����B�ߩ���~+Ƿd������r���.����B�ę,%b��pQ<�{M��kP�~cC�{�^r>�7�G!�Q�>E�N�Pl���C���N~�&P#J�l<ضj��r��|��LSVA�cbKE�Y�4bc���ū�:��&��*����%I$�Y��\�=��uȇ �-��r�A��>�1󋡊\�'�������|��4�gн6
��͚�N�P�	8���s��X��b�Bz��`K�fQ�	fÀ(4�&����C-�J�A.¸��4��V}(d���'n��1������nǑ���ɶ�5��HG%���6K�`ꁩm(C�R�	��������w�����U�eK�"&�1oK��^�\M0'�F/��}���T��|��AL�fb��3
��@�]jb���E 1�����%�L��b'�>�o�l�ʞT����3�����;#��[H8O�.�gl*ZSP:`c���T��@�<�Ī����VJ��7.��h�bq���
Oĥ�t�iNӮ�;��������R�zF��.���$�4�W�U�G	�0��Cq����[m�0���>*|۰�W6����#�2ip�K ���H3����d��9��Yz BeV�����@'��)�i6XBи����WC�$�g��6�3p���9\i�@���~ݳ9���i 64�f�}e���i��XFC�f�m�m?r�'�Λ�*Ww�9"�B �v��B3���C*��[� �pH�ي���~*;�j�._����[%BhB��� Z+/Gwwd�;cM��?CV����H�C)����SC�� �W�Tc+#и�wfe�� [� �4�^��D9��M�q�O� �]�	1b�e�3+����]2��� ��E��8����lS�޸��`�T0 �`��q��V=���"̉�g5>:����زdC����kpOr���'�`���p��W$�.]�g��ەz��,ZS��
�r���|y��TQr8�ν�t�y'�)`a�c�ʋ��BT�7��(_0B4 �}�{�W,�d���0�q�2�O��Ь�g�С:���E�%��p�^�����E	jZ_�o�:*f��7�5�V���K�Z����5! �-d���!6>�ݍd���oD>
BYR���R1U�!�tT^Ҁ��4��|���������ȱ�m�)������dx�0��H!�F�ES��0o|z���6=��i)tK~�3�BԷ�{J8�0'K�o#GE��˹�0�n�gօcQ�n�nPeKf���[-A�L:'ܢ�__֕��g> [oW�B�M��&T�2�PZ�P�����@5�����������P&�/=���G�m�1�����Z����6��I5�V�z�P�fH���|~�����"�-�����n�P�U<a o�ݕR�0���p��A�b�~ߑYʚhW�@��{��AǍ�Gj���*;�=B�6�*�,��V1z�}B:AYΌ9�8Qi����e�sk���[6߂��R�0�K<�����~C�>*��pܙ
/]~�U�aM��*��V�6�j��\ukA���)(�y����S�}ʰNAu���K^�d��^B�i��p�+ro�C�^i$~<�da�:�7C/l��,D��#LL��ni�G<G�wa�}�����M�|��Z�;��,��wE�k]+4 �\GΚ�*����H���׿a��7ƪ-���bQs� d����s�.h@{��AC�i��VN�� ,��b�.+�Y(����Y�ǉ��	U]�А[B1����J[7F���aQ�fI ���;�a��H����&-M��<Q��X��9�(}I��)�0>_��f���뉍:�ȈD�/�W�"#[��t���I���ʧ��dU�t��IA�{cJ<��X撓3gi*ڄ�O�7�A���~d����d������r�=s�y�`�m]���MS�=��x��_�V�q�����d#[
��:@T��IfP���$Ul�.x��w$QW߼LM�Lmc-�'>(�����g�a>g�-R�GHݹ����Q/��N�+�q�����+�수i�[�����a����V�۠3F[���b۝:,ɳ�g�J��t��$����f�����e����yJ�ɑzɜ{aӝ�ԒQ-��y��]����YibY�L��<�q칉O�'ƺ�lUN#��~\�aķ2+_��f^ �@��C��w��Ċ	����u@(b��K��׍U$��m� �tdy�I�W�?��PdL="��\Tx�Ā&�Cl�I����:f����#�F��z�~��B��}�C!�Eh�Z�s����R��������[цd'�}�!�.�������vL��05·geȚa�*�����Uӻh�0?��owK黠n�Þ�H�	�Xbr�^w�?mlY{��?�E�B:���Lmc�设�~���<j⚍�S:��k���z��w^�f�o�<cS����1��8ǻ1V
�
��>3Y��+'��g������~f_��b��[�����v(�r���br��0�M�����4c7��^�f�@��9��J�R��e��;��9��A��lu��г�[��+�]2��/^;{jkv����{
���(H������V��q�[�?|�8 x2J��\F�)�	���n/��T�!��v�>LV1��[�wTX�?�s��Z�����sM[M |"Ĕ���A�X���+�&72�;�Ż�Z?GV�P���V�H�|%AF�JJ[�i�v�Տ�ҿNx>X�|��0�$�$N��[�y;�	-�M�u��RV�����*�{���X���U}��UY4&*竸�M��_�hF<U�1c��y�F҉��K��z�in���~;;#���BD�������i��s�8�����M�9�����|�Cv@-�No,8G��*�J�[g���|���͕GG�n�HN��氟��_E?[��fQ��{9x�TksT���L���.��s�	�����n)>E%PV.�s)��D
7�+��:��?S�4a��hq�f]\��d�w�yl��"�f�:t��^1�Ƭ���@4B��6�O�o� ���%�V��n�[M�'��#���n����*ڪ���b[f��㐖
��3�SЭ�"�ՁM9��6 Z�ƶ��ڭ��=F_<Z���M\>���d�E�z�� U�OI�Ixp�"u��1ݷN��oSy�N\*�M�E�ɇ�������p�D�9����).�|��&Ϝ`.O��oh?Y4���;���֨=��+����g��U�8�O�L��{@�a�t&ą�z��Iv�Dsݖ����i��ʃ�jmQ@�i��Y���1گ���\�)��קU]1e,,-�	��q��:����V�}>y��� ���Ӂ�z����r|�[L����f�����	0i�]n��BR�I��v��!���*���ږs ���Cj����o�M�x!VD� eD���$U}J8eaXM��?F���n� ���&0�bσmk,���|S@�İ	p
�.�<���m�$��?'~geI�7h�I��� Wf��yJ~��%�N\Љ�i7����m ����]$׈���%�>�}{�A�m�C4۟�;ufQܼ9a_ 5`�
(����u}	�1��3s�H:Q
O��IH"��@�RmS~��`36G6P��x���-�Q!Z��Q���372�"� ظA����W���p�xI�#ٴ��,`e6m��β/��ֳz���Utn�/�:H+o�	)lt4���M�Ԩ��R��ŭlG@��#$�ī=�'������qmM�K�+��yi|X���nw�')s�1��3E�Q?��7Mq*|N}�(�������S��`[��3+�q��y�sw�<M� ��=�o���9I%�upD>���d��Gm|�ӓ3�VbB�6��lo�r3
_tD�U'����c��?0����¿��k�]C����lMH��G&$;�s�}�6��b��ڽ��1��9X��G����/UDZ��>c}ݫ�����(x�%�m�)�{r���|y������(�WK�%M9DyL�M��z�c��iu��%~�W��D+"�b�� ޟ؝�!�=KQX��s��
���zY���W=�t����s��=ohFJ � �p��Ë��FK}��n�D��E�F�_HI���ؓ�;Ӣz��/��ĿL�=����|�ʤb��q� �B��A�,U��5��^M �*$ XX.��#g崅���m;��\*W��;X9Xo+��'�"�x���|�
sq�|�ϨMle�Qq#l,��F�.���6J�_�l��!��"~�V�TPvb���#!�T��S}�C�* ���pcs�d�P,G�M�h�=D�H���r���>q���˧�>8��y{���KMZ8n�4x�ņg��Oۖ]+�3'��S�ؒA�Q�nSШ����Sl��;���/�����*G��ti��D1R����ׯ/J�0���A������������"JeyE��1���},!ct�G�N#�	�Ν�q���a��u?w��@��mF&�b�ۧ�9=�W���l1dC5j�pN5���Bܰ�סHWk��]����K�b���
j��XbB�w�׻�PϲC��"�% lb@�"��b壸C�ݬ�4�
��05G-��v��k2�}m��D_j_������dªS4!��ll9�oٌ�n�|c�����E�8L����.�l$�Ib$A��QJ��3���[��|�!��):��Q��FhL�e�NO.tq�6 N��LާFe)�Z�����oayJp��}OF��-Ve�/ҽ>w�	M�48f.;y=pAן�a�I=ryk��� �c��_���;۟�C��#��������}R��/��X5��Y@
�&;��CR
�qF��B�f	~.h['G��$>�;3�EU���	O���1��E�!�!̈́yH5�U���ˇv���l�9Qe����g�f��N z�ODLa��C2a�l+���9�!�#>��r��6DlmY�?��zVFB8@B)j�v�Z�ԕZ���z�)&�@Ŵ �Hk�^:x�-V�����}�!�
�5t�E;!5�O����s��S��)p���g(O��a̉��[�J�ߎ�����%��-��_=�쌃���8��,��˅�6n��7^���%rA	f�h���+J��P�]i1���MMX$�@L�� n(��v՞���F�)҂R��5^.G����a��D�يW˥��a��@K�+W��Z��d>k��-1�u��`�}t�m���5`��6��D�e����K^��iBF:%Q,��ܠ	1���M�
c� -h������?}.��z��,�\Ҝq�$]s������08�~�>�Rd�����&:p$ �^נ���Ma)�����o��S�N#�
VӴ��	߇��c��B=���y�	�	�85w	8|���/�~8���� 07��!��՗r�=̂�7OE��ߖ�p* �vQ���_�3��g�2��R|�v�1��������C���r,r�, ?i�6��C��.Ӌ�ʞ�\�w.T�5�X���X��*3��:	�Sζ�K@@���k�m}�z���kf���$kh]
���Dyg'D����i:)�1��^�8���k0�4�ȶ��`KU�qJ�A��tT���*2�h��:}nY���u�9���<���@)XZ=8��s�qwwu:ý��\��T;�9�J�=Q4w�_�ߥ
�"�^��T о��ys�_1�Y�^g_��aj����'G�&��oK-ٷ�:T�[$��M��\�]�ҠUҷ�9 �j40ٚ�w�/�9�.M�6z�20���eF����8c~���4��(��I9����N�)+�AU��_b�x?N���i�6�=I���F�&�QH#�����~eM�ՋR��˫��_�O����*Kk4��|�a��VϞ���z�"�i��Bc��/�x�p#C�����5���)<Ɋ���t����l{V�$#�*��_��\B��D���KI������$���I��SN�������I�6qE�繎�[���tm��[�U��}���ړɧ�t�@YnۑW���wvf�3uԵ����p^݅�ڿr���y��:�,ؑ��!�U�$=J��>��i���H�ӊ�����i��*�/~���$zA=<��l�4@�6W������a�ɊS^u��6��x�YT���#^Fܖ���7���L#���M:r5�&�����hŊ���#O1!V��Z�v1#~� ��������'	�'T�u�gU��5�� +?�iA%~�Ae�a���5�i�U �`�jJw�{���1��IC�ʱ;P��5��]���3dt NF���u�a�n�+�ߨ����fKKX��c�y��jg"n�c#�.}Y6�=�|����3#|�e��R��T���"�ft1¶"�`O�E��j�~?��G���a��2�o�K����i�^��lR�h�ɡ����g�H:�7Һ[�U5�)	�G���X�v,����� ~��|�R����p3v�lj�	ġU������#<�a��l�G�R6B�B|<$�SJ��l�{O��	*�ݓ�%M�!t}j�".�5^�Ѱz��a\P-��Ax[Md6��ݴyV2(�__S�!�������z&�l���� �KL=
�ե�x�.G���LhJ�����'��^����w$��o��s��� �aQ\nJ
pC��b�1���q"|J���oѐ��6�El��0�G��Rp�����ΨN��C{��ڐ�a�s���6?2:����k�E6�G�m��'�^�:eY-u;�^�{iţ�~l^}��B EԿP�q��R�fdsY��mU����ǟЧq��J��p*�EK�N�2�zȎ(�=>�+4�����fd9��F�s� r����A/��4����kCV���AW�1&$�2�{�Ĭ�Ξ� ���q@��])�� } ��&#e��E�=v~��8�	���#��iX�ʳ�5���:���s'�5CK	\d� �B��]��Yx��P�9��%ۼ�{��b�@�-<̭��um�#����ph��H��g���kvw:H����W�#h*�+c�0|�a�!���r$rY��}�f� :4�A�1	E�A��J(z�!ӊ׋a��y�M]T�o�>sN��J��o��+:ӣ5�1��bi?��@
 b�[xyx�I�F�JE/����""�����V�V�l�avrZ�Su�z�s�y�TyC�n>1an^�C��������f[F��ີ����g/��u�7�A�g,��y�Q�
�g��s[�ч���E��9�4Mt��+��K 1�8g�hP�!�m�.�u�z�����y�'nG=�Y���^�bQ	��Y� '̝G :b�|C/�]��''�q��I6C��rz��X���K���U��X��|��mC �M�z�/��e��!��*?D\��=��\w�E����G�7��P��v��b��q��ʤ�7�#�^���	�:r{��p�N͌X�.tt:
�͉�2���+��0$8�9���j�w�M 7�j�nq�S��t�e�����<c�H���7�1�yvG�u�HDb�HD�l9\��iӞ��'�
�]Uԝ�����⎁�Xx�Hi���ȥ9T3]�]�N}>���%�٭��������
σ���@m������[�JlZi���!"Ƃ-g����7Z�*0��\��ܶPϠ\�����\7$�7����t#swi��B�I�7\e{��+b@�z1e0ԝ���ĭ�5%2�U�T���96[Gy��U�+�!Qm��ca�BԹ��� �NݺD^�[f���������(`0ѭa��k�@���3�),�+���M�b½�Ůd��N �.���V�H�o�R�����oew~���9T�3$���I���Zl������^|�E�:���2Q�UQ��>���6ñ;���1���<����������ox\���R��N��@���xkJ�t>z�F�<�e��E6�kp0�V߹֪R��wJ��}������s�o�.��?t��3��l��q�~������,��m�y�X����'� ��%{Éz�Sg�4�����C�~�z"���y�:}����(;�����OyY�� �Z��7�[5 �=}VwXp{λ��d4��k�[-W�E�X��#jE�SVg�؟�S"4�	Ph��O���?vwk����8�VV��>P�:�1�Q��XNB���p�ʙ��P��>��c~E2X"��R��ۊ�� %���TT��CMc�o��`y���Skty
�$�1�Y`����G:P^i��D�p��݋A)�-!tI����5L���@f����κi&�l2��v9�DA4�܅��n�3f�����><��Ř����Jõ����E���e�oW�r9��Rmp���WdX�%a�}Ҿ�KI�AA�?9u�Y�,���k��A��j��,b+���z*���.����:�n[�k�A�'t*�\S����1b�ݏ�wR�zX�i��;Z}8Ouݒ�"�g֨���'m�@
D�,�HV>�}�\���@�E���:9N��["�b���U?�8�EJJ:��)��>��R�2�4#��w���'d�/%��X8gK�R-�@����̈́�X�%kO���M��T_V�x�i�ȧ�
�}yѓ.ȣ��Y�����	C�z��һKZ�X��w�G�1v���3������S�@��v������g�RC'�����S��������������Aap^mv��������uX�L�b�ͅ���A��	X��N�%΀��m*Xp���Q��~.ț�y���.��=��G�߸7�%'v�
���W�q5����fH	���qDep?��l+��m
�l��"i���Ɯ�e����銎�	�ubFR����R�9b(u-��9��&���G���0{����#Ψ��x'�����Z^��j�m��r��*r>��C�얣@ޒ�|����Yc�1Dh�ޙt���mAg\�L,�e&����8��
CjSSoB�_{��[6�m�O�� ǫ[c'��/�ay[.��hDm��`ı�B��(V /Ck.x��*�]���i����7��1ӹ���E)_�C���>�N������QMR��z{bp��Ź㕮y!���6�0�D��������4�F�$E����1��7�/���]���>��� .�0@�g�)�_��l��s����_� 4
�ڥz�k�#�	������i	�9^��`���da���%�q�wt{ "�L�b����\2Y�H^����/{����`��;��^��R;,;&r:ç�q�~j�H���K4���%��'rXJ2n�~Qf(*�?�;q<9cJ��ጉ�Z��8:
%�ށ]W2�����I[|U� �/��A7g�ކX�`�ܪ{A�P;��Zg�6*Dx�R�"(;+Dg�yV]��ڊĴA�o�����5�Έ��}���F<׷��fe%����������7|�i ������ba��i��~{�x���%I$o/f�3����F����n(n8#�Z�"L�T��獆�g�����݆i�*� �*���_��s����s�}T~�~�f𜲟�}J�l��k��}\\Ѱ%��j��@I(@P�5|U��aJGdؚ?����y�7F��X^Wř�Hd�O�ן��+F�ӶE��œ��%�����b�p�)��S"Kd��2?�������68{(����"�*�2K���M|3����?J}FG�I�m��hcԙ�� �3�-CK���H�r74�4ߋrg�Oa�!P���������uz����q���Tv
cF��m�{"*j`>�63��"�kS�S����=-�Q�A~�W Ӊ���ϩHoP�{�7��c];�� |	5wE͊���7){�����b���J�܈�M�6F��A�<��`��c����$���\t7�*���
a�	jhG�s��Z�q6�-̐i������Q��o�>�%��hcY���_�FH=(#kHC�����U�i���������k�5A�wnFx�]���lS�v��|�S�T�&��dnD�;%|�(�M4�����K&�Q���V��yu�*!X�#>7=H�?���"�h�7}��WW��Y�y|:-{��(���z�%.K�̾�O�h���f�}w����͠��	*8��e�y	�
DR�&{V�5����?�vI^�l�ۣ��bG�
���k ����J斑�9AD��:��|2����K7�� )�r2��r����;�8����- I@,�뚕O �b��w+[��z�Ek4�G���=�{�����-?ӳ`��8� !*����#�_�62K@������ `�&[ ��`���X�Ź�8�v;�����?��g89Ɯ؏KzM�"UC�N)tr�.Ʌ�Y���!y]&��0g	�/�G�F�B�Z�ڦ!d�J�K��`ro���?��� �M*�T1/c�]��"O	D���	К���]��R�kh�j4&@��+Su��Co����0�,��YR,���m������m��Pݞ3�5�H��p��sK��w�@򿤩���_�CH$�i�r��J�׹.vS�-ځ2��0�ݫ�g�q��d�/9��p�,��C�_��?����ة�X��Q�A���h��O�}[�?<TR7�Ĭ�DJ
e�q�F7n	�o�MU`=�%7�q�s��(d 2�C|c��$�-}	���bzw�p�������MԒڿXj�bOv�j�(:\�D�΢@ �];�A�������>�~T����1�沚R.��o�'�w��^�*~��v���}��(���9�ٚ^ᝥ�k{)b~����h)��s��{tM��T�U����}���6#�
&�a���H�Ⱦ�ež���GvW͕����Q��0GQC����
��ϼ��$��M�@T�k�"&_������q[�.Q��<�_V7Vo��uDf���+ӹ\#���9��C�53�Zc >9�����W�Fỽ����W9!.u����l:!�@A¦�����b�g��dJ9~��a5��;7��t�����f��-/�*j�4 �-�ݗ��A+s�	0H� Me�OH<z8��v2��O��|�QI.:n5�Ջ�/��p��aQ"�y�n+;���NzN"�����`q# Rq$-0ê`Í��C�xK�ԤE �hv��o�:�-��?������s`+7)�Gd��u������JҔ�||ѵce�@�߶��z� ��T��m�ˁ,�b^1�9L9;�M�uA�wT����YV���ڷ-��񜀟�����!wQ7���Q��z����ϖ&��B��e̒���[��%�U����=St�����f�Sn��*��:�-��{s��Ʀ��T�l��-��%y��3�(�!)���G^�E���|��P�yy�Ŕu7T����l�������/tn!3��j:E��a$��9��=U��?���u�0�c��e���d3�4i����UA=&,�r�_U��!�Uw-'P���g���&�^�(�q>��m?�z�cgP�υ���At�`��ѷ�EZ��zG�h��i.m�2��������t��͍�zBr���/:���S�`L5o@!+�z��d}�s�:�]���\ʀ6�4i��½��_S��~5�����N�+8�(�������&c;<o%���U[5����[3	�33�kU��pjF�����:��2Y7M�2:4;���T@�\�j�����?�Hˆ�adY�1;�
�j�,#G�S���,]j��Ǭf"��T��NL�zDC�����QPy�s��x>�'N��B���dFg|?I�t�=��T�`��Y&
C�8)��bN��֗����O+
{)%��jQ��������Ht�:T�KM���"�_���Ҍ5RQ����f8E�
�s4�eV���?�7��M���`Q��v�2`EO��Ǥ3��nQ�tQۄ
8PRڢ}�/�IM1���ҽL̆Yk�7�o���&�ÔY�H�J�h�z��mqI�{�^u��;�4z4�H+ϻ�Kۧ+�^Ԩ�#�N��ޚW��6N<>R�]T�@��ϬyQ0|�#�.:�c3�a�#�s�9F�×����KO����<zrָ2������a�C;D�!zS�S[����'�����O�vnR<�ȧ��Cl�P ����N��Ҳ��i��l��zD�&�^fB���S��:8�W����:��:>\5�cvϳ��?c٣����U\���+$9]��!�v�к�^���C���2��w�hV�*A�	�E������:4B!��@���+	犺jVw�0'��P]pHSb�{���:���C�\����̮�7ba�Q9�qG��|�#_�V��(cNu����S�x���G����	z�����Y��L���[�^�l4�����@O���+�K��{�_�ڙ<n�J�����_PϚ�����wE�W������ed ����~�i�@P$eq�IW�m2���Wg�r�����~QxL3-l6af�5E��TQ8X�Kx:������������å�l$�9%y+צ��VJ����L�bD� q�-Ӏ8`��$:M��j=ɳ��|�+%l����[Dg�Y!�g����?2 �Cl�I�������<Ͱ5?�l/��v��Fm$��]|c��5��&��������������P}Q�:8QET+���>�@��`�m�f�$!@���R�N�\J�š 5yh����H��� �V�����p]�� d=�'���|�3He|g+�o���jE�An�e�Ύ�;����i���D�,�
�&��ӶN�oY_h�5���)i�7K� EOSٹD�ZY��"}A������s���kd��Z=R&����+E���%�s�0ش�����f�z��l��-�`�*o)w�9�{�l�n~0'G�ݎ2$�k��ȭ"���\�����_Z�C�Kp�wX�$L�F�^����!%e'	޵���z��/�7�{g��8L�����-�U����Ղ������3�DzO�9��;ƌ��	$�&�}ɒt���]�'a�'�p�?�S"yz�Y�i)I�,�M3-�b��~2���Sjo��A�>S��	~���g�݊,Ӆ��"�9W�^M9� ?f�ec�G�T� N1�W_,.,ꆊ�S�Q(�Oe�9��!�J��q<�b��M�:���W'��|_���;rt����� e�gH{=��W2���Tϣ�KD7.�'jA7ס�3]ʫl=,��0)�Dh�x���$�<%gT�m��0���ƃ�i�L�����]�F�6�4l���8p2�1�ࡇ�H��>���O��#H���"h��m��WM�N��m�~-��o�Ġp)�8F��/���iN��8T�~�w�&?���������ߞ��A	�𶠾���s?M熙;i􈲬!/���'c"[\�m�̾�ʲ��!�'�:���y�˨q�q�?!��89<-���q�t��K�<������=�b*��p��tKi��%�,�,δ/�qN��~j�-����I�ۀ�6r��5~.z��$Jp�sI��Z�A,o���5��)(�NVtm[��	����F����f�:GΌ�8�(������׸T�E�j�lZ�iS԰5�5J��5�+��Ibnq_�-W�UN!N^���@3�"
�|�c)�(� �]�qU��(l=�t�������l��S��|��Q�D��7P�:��n�H����`��!p��Z&�:B���C2\hg�6w_qT���ڦ9,�T0��{YR9�� �Vۃ�P0�Ö��2��Y��4�#�����p��s'1Q���ȗ��B���_P�ܫR�n�W��W�SWR�\K�ֲ$y�'q u���M�d��w1�)v���(����"�`>m��魴��v��+X�ln��$��52Y�L���Ao!%X���d8x����є�zx+��
,ϔXUy`+S���U?z�^;
�P2u拉@Z��$�*T|��.����n�icnX	H��ɮ"�Ed&@ǲ��3Yo?�`H�>��5�h<�0����hK�xHp��ؑ�tn@޶�� 2 �B�.<�2R�R�(�\�� q+�r��Jhv˹2<�]p{w�+�<�θ�U`��n�9���/ *mǸ� ��r?6\��O����R�u��o�|Υ�����,k�(:F�M|ƅG�nC�)��=�jh�ðʿ�M{�=�Q���a~v���P�0V��y��|ٜ�KۆP!�<1N�A��&�eZ[\�fiJ\������}<Z�U�o4f�t���Z����a��|�!:��Hi�&3ɳ #Iߍ	cADu�=� �t�_�,h ^�=�ŃT�ҏD< X���<Q�Y�oā�Y	��4P��|\͑�a��åi2�e�%�	��V��]W<!��5��Aŗ㎙v�>m� }!�t����¸�T,kJz�.�2΂����/�;/S�h��h#�w[N;�4��)��P�Q�lD�]��iԅ"����8_�a�A��Ć��w/�cZ��|N��b��:)�0;$�K!��4H�]O��3�w��ǅ���`�w@u�Q�h������i'�D�ȞJl.*.�H#���cA��Z@�b.ZF\K����/��8)�V�_��.���+bÂ���ۥqé�5��L�t��5�}���N<�K�w-�Nn����RC���"�&���D�PU��0�.�B�l筊�/�El��>,v�q����2�T��[��SN) �5������bЈmY7���,G��z6��{�E�8��d�q��?�ߏ���@{B߁D��r�����j�Q��T���M����(��F�$R+��(K��� ��.XE�g��a*�#̇L���ۤX�F��>�edo�t�Fo�E{�}_�١����K2�A�	1�aEF�])|y�ztM�%��zԤygG��A�j�*{F��� g]*�'�!"-c^������/�.�=P��xr��y�N����I��$�0�ʉ���1E� b�'���TT^��ƣ�~̩�cU/kB�>G�k��x.��M�u�A
�{]E����,����><P4%�����)� 0���Ѿ������
�J8�n>��n���x�E�Rr��O�#xy[��_�WF��A�˘,�(��CuMH)��yW��$�{e�8k��.gm�-�<&78<l�n[E-Z&<�Ij�8ѡ�\��̭	ȯ%l�hϸFH�R�vuG$4>Yr�s�t�d��UdJWnf�Z�oه�=%�PFƘ|�m!�JVX�(�f�@��!�D13��za��r���3N��:U����9���ޝ�:f�&dϰ-��dzo.[?I��?׶$�����Z�a���Q��Zl�os���蒼�����E�����Xvq�B���z��L����5}���`�P�} �D:N��ҹ����Ϸ���.0q&�q�(�AE�ZY�����:���k����'1Z�T+z�NB��T��Kٳ�Ч$9�3�4MRy�8���(��C�� S�D
 �^�^(	��OQ_k�mB��%��A����Ў�1�W��%��69�Bx6�)X1l(��h�Y�thl�����@��[E�� ���}�ICW�S�1U��K�a��($��׍tb�x칰9��S����o�a�oA�i'����m���H�b����������X�'*A����_l&����ǥi�t��?���^�g��=A~�HA������h^<��]�I�O���w$k�y���\����?��0�3lғ3~��m��P~*����/���v扬E��K�jߌ,l�n��P&N�m,U����B���٬Nݕ��u��lU�b��J�cH��m@ߐ'�L������}�rwH�	�\&�_�x}C!��f.U�����Jy��	T�%л�d�,��\��(K�8'D���q]��j�G�S��
w�Ý�Y-'��3Ex��7��@1��QM���J���LB�L�|��W�.O��!�LW ��2����t���9�S�&Ю���i���=Ħ����gҵɦ	��9��l�91�q\l
v.��\=r	��7�eА���M�%R��3��.�
�S:q�Zͅq숙�x����5�Xl���E��#Њ�"`��Q�)� ���l5�4�%���A�OY ��K���:��[�V&|8��n��˂�ϟ_-B{���'>�I�*҆��9��~��2����q!ҵ<�*�{�H�.�D�'�Mz�T�O�!rpaa��+@o+Jgp��cv�=kܫ��`�¾R�O�i�6�61�j
�5�>��`)��U�;���F�,��;6��U"�>�H��T�/e���1$�=5sw��1NC3��)"�mp���p�����	���	�$@H�Ӊ�����f��Rn%�ς=�?+�J�aX�z�U�x����Z��<���zYѓ����Ab�!s��ͭG)���=)�9���k�ަ���T� $��"QFE����ۥ��n��獴z��wxv:��W�2�l�]s'��=�w��![�S1W�_��}
���8u�(7E�7^�H����]|j��q����H)!Wbos�MuI|���	4 �	�੣��~fO��[rC�ېup|M�2�6R\Y.���1�8�5���T����4/�P����k=�Nĉf��4����`��`m�;i�-�������L޲;�З����
@�=1-�!�������bwj*h�z��ʛҜ�ͧt�v���G3#8uf[��Ac!� ϱo��C@y^���EJ���̈���a$po`�Z(dqĖ�o���u�<@���z�(�"H00���y<��J0�����y�4a�ozb;����d��B���^F��T��m�q���%Ro�D��,�R 0,���꒍˾c����}Sm� �CǱ!�M4�/��r$a06����d������D.0�sd�q����f�@:x�7�69y�ؑ��}hH ڋNx<��Ɂ��{�5�.F���� �ʟ-RQ��\����o��J�E~�:����p��(&Z��,)�9�Lt���������p_�4Q�)�X+5s�ѪO,kaC"M	�bop	E��߄L�-��x�ݨ���0�&Ax�5��ʯ}�5�L�M�6��v8�S���&��"�懿L���Ԗ*�W�R�\	{��JD51ۻ��t�wFL��d�R�i;�,�E�B�\������9F|QA���]�/Y�d����hxV���S�����1_"~#?����|	[�bf�F��{+��D���L
��'�,�[K=<u3���9)gxrhբlg}EҌ�nα��U'��b��TK3������X~�̃_%J嵦=����R2�l�%mr�Ab�A6�(���?�F�1���� q��feSϾ�2�=���yw6o�B���
( f�hϙ�"���V�W����t�_@�'��F�ss>��`\brU?��=þB6�,�;�=	G�W-�n�^z��G�j"�9�>�1SDSsq����L��|�>&��lycJ�G����,��RT֤H���I�����d���a�r���?	�~�Y��+8�Kq!��^ n�Hlk�|c(�n��p��{���r+���	���䑟Ä����������Yb��샬�G�Q�Ϟ�Xp|.�Wd��Xk�`$#(}gl�/%;�ac~f���s2�h��F��t9h�a�^Q$Ϊy�H��;�7GP������6{pQֲ��H�v���̴\~� �"�#�(������%1o}[4f�
}@%�п�r�jA�ܐ�B�����0Ne��o�e"��W�IKn�/��sV`���)�:�J�祮����K?5"Xqw��;ŸDQ7�=���@�������,A s$���w�3`��5ϰ�|�ud4֢CG�ON��}H�>�\���e�AJ��(��X�
K�i��c$|m�Go=����K$�XjU6v���mYX���O����p�:�N���8�vf{�����?�|�h��R̽󗑩m>S��0��F�����Gd�O���6�*eF�q�e�8�]:Zy'	�뱽��j�]a�ڨ7�8�z7�T���v�J�ጼY�P�|f/�xYRE� �j��*X4Uk.W_5���_�m���C���o4:zwi1��:�����Ե�G-b}pw�YX9�\��l�R��jq ���9!0�"/u�%2u0k��|�R[\\=�ry9nt06N�P���q	\�~UW�V�S����=`�ha����B@�W#lD>|��E��O\�(�;�y��5��. ��S�&��Mɯlr������͹�2|�p�X�}�q���x�,#�g��%��PlZ~�I>eH��gl9�	`$syU�o�u��)�m�^1=c�'�r�Z�,�\�諔�l�ũg��'�B�!2��t`���ߚ����PL/��?�en#v�|D�|�/���$D3�T"_�h[��@04 at��5�ƖT:�����P��G*��&Ƴd��L糬�Oؖ���fі~u�y7����E�����O��n��y"���2%���;!���#���V*�J���V�F�ɜ�3IY�濘��R7���!�i�e��b )����4�����6aȦY���E��//ǿ���;4����y$_F�F%A�����k�L��A�a���~A`	��7m^���,/I"Ws�
&»�!X�#�;���ܷ��_�Z��,�TL4ܖmU�m^�ӈ�d#s5Q${y�0�_c�^q@�:�
=$�����#�Ro�e�w�W\M�;�����~���-�}�,�b8�<d�		@O�
�XDց�^�He:��
{�
l'%�v,��	B�GUr�����R��2�h�B����ToeC\�T��l�
�frLW�6�"�]�N�˗�m�ԕ��o�������AG ��$��c_5��Zӝ�xg���͎����Y���l{YoU� ]�oX����O���]��,��Amw�9����m]���Nd��]��,�vӢ0��Z �.�S�x^�4mxv���9XۃJ�<Ղ�8)��-�o���^{�����e�����#I�zLaK���U�?悲R�8풦�P�����$��H�Z_Z[~����c�DP��ْ��3 ͐0�N��+�Ĝ��#sQNpl�I���������%�J�QC��t�.V=�4樔N8�����2 =�D��f˹;�{��,�i9�0PHh�{���FzH76���4�{�Ԩ^VA�H%����9m}�yD a���6�b2�ט��� n���&�a�&��;����*����c����U��յN������0Ya:��)���9ɄH;$�z�|���f��0�L�4�9nh���Fbz�(=�V���:�$?�{�Cۭ�<�:Q
���]Gy:"~�Rj��~�ޒ��#�5����b�?����'Ϊq�R���R�����1�++b�`zI���=�([�L�d��@"1n3eˍ��k+4���I���w���Y��1S�R��*!�U���5�Nf����.�4#�Rw�YJ[2V��|oq~��lX,�a������'u2���B~�"U���C*D�����l���{���W��-������;3���}�nM�ز�����$P�W�a�7�}"��jY*}�E���ڄX��e7�A��W9<��=MxO����S����,�������JV�,g�pz�����s{�����!�R|t��:Rok������gp�2�� {�k*��+*���>�t����ϳ�>���?�S�*�Ê���l�	M0zy���V����}g$�J쐟]VKO�h �2ϭ?ac_�����j�R�� Mէ*E�Q1�/R�� m�՚���	�=k�{r&O�������}2܏;�����C�`����#�#���d'x����f�.�
lM�^n�	O� ��4@�]J%<mh�~N���덏�t�b�w�C����s��=�ܝ7�Fo��9��I���d�(�Ws��w�W��j��f�L	}`&��ەn;�����e[��|f�ր�NN�����A{�����s�+�*�;�ﳯ:_�O��B�#�ED@�[���r��k��T�����x��P���a2����I�4��磬�f�AoM�FitP��?ԝ��ݏs�]a�>}�����[,7�gEO'����^g�O�R�#�P5��(!�ж�����O�����w5��,[�$�O"�K3�$�x�� ��&�F�}�Ek:PM�I���(��O�%���`[g��}�f� �M��$t��|�3I��P.�����gq���}���<9�E�<4*<�1ȈX�3 �Xl��ݝ|�ohOm�~����᥎_t�V�a����"�U��L [MeZ��i��h(O��I��'�V�fv9�*���|�X�=%��=8�G�'g�eA���tsd��@qx��a�5fʾ䏪e����Ԅ��^���fR�@�s��k{����!M��ܥ{*�e�--�J&|�������/�T:��[.� ��5����R�4�Z��%��`�jxS��6�B~
�@c��W�z�<z:�IH��Ğ���vE�ȢS�kS�F?HD}�ܮ����)�"�3(i���S��$��z�y.���>���s��u�"uɓޣ!��W��W�ã8=�?��>��f?�`�Y�����rl�!�i/�O�+��r*J밴��z��oVu�u�<��T��W��x6'@6��~�r���]Xu�Ӌ)�rF앶U���D��bv-fD��*t�o9W4��+�n5�d3��!&���RW%��4~>�yl��Q��A>�g�ߞfe�݈]�Tc��sz����_1����G�z���a�-
_h� �$�qBR����:~�z�ǳVL�qN�\R>O��8��Ga����3�`�QD׈�a�� ��]R�@c�ص�ݓ�����T�ǖ��_���U^���[���:%K$��^�U�K�[�n��+�4m4����)����e���1��4q��0_�����^K��LF{�?�=R�6JѝW�� <�5�r�b�4�ʇ�Q#��T�B�b@%3��oC��9�f��ʶ�������!J��&�!lگ���wL�RCh����OA�)3��W⏑w1�4�g*��)��+@�w��:�e��_N��B��ׅ��K�&E�n� �k�� 3?���Г=�F�V(�f���
���Ƞ��H�O�9�䢒?y��zsv��B��Eن����}��{-Qͺ8��v�$��St�s�F�[��`3�	���|�[(���V���{{1FH.����	���cg���D8"jr��%srt 0;�۬_��o�sC�+�����;3�COs�+h$D�K�z�!�ya�F�<��#i*a]DU#��^&g��W#Q�[�V?}��#yh'����1 �Pˢ�UF�����pv|�ng���]�����%U�Ux%v�˓S�*��*�+�B��Y�W���ΜQpU;6L�q��?8F�P�!M�-�),=׾)$��S=̖�4@�;�D{�$��ں:��"P��
[���y�>fM��s�o\7,y��ce!��͍g����e���P�N�|�^��k�C>dP�����D�^A�Z���y]ſ�ɦc�>g���h*Ŵ�#��q&��H�Pvf����W\q"����:J�Å<�hƘ�3�7dO�����4�^y�7��U�%���	�� q;J��&� (�=�����\Z9eJ�TvJ??1��sA[t6|l�˂NG$Tm�&Q{�1�����N���$1u�@&̗h":	l��~��ǝ+�-늌;][ꗆ3y?B!C�M�����]p@�l�"h���s~���MI�PP��P������?ao��o��S_���pN�ĩSbZQ�����E|��{�W�F#w�AxC��ci����{퓍 �g��װ��h~�W^� 4�j7 ��thP�ա"�~%��c�8%O����R�Ū���l8�>�|�9�s��|����D�O��!x��5J-���\�1x�h��k�n�bS�:��Q�?���p.⡄�!$z�.��"���� }[M�����b����P���� [��Q�����)"��9�֎�;�..ƅ����>�oP�<�HXx(Vzw0j��%<A!ߖ�����ɧ<}��{.�k@ϭ�~�ʾ]0J���P@��	�;�U��b� �ʧ��+�����ӯ[%� ��Q��jA�MQʠ�şPsn>���	�U�'�S��=�����B5+em�,y��M�r�d�T囹r���.�1�lb�~�⠀�*f1����U|f�o+�h9���}.��}x�5�����Hme���|�������~���w�斝�����U�s�+����*�o뙪��K�jX!���3P!��K5F���M����Z5��թ�nvW���;��'�����S�#Y���S��7��q��V�̸�^U�9��Y�tj�z�����]�숰��L>�Y�$�N0ba���'�'��TM����&�H�~̸!O�7�/����/ɟ.�OĸQ����I�&�����6�����th@�)ڃN��� �1ǯ�m������݁8��k��ۺk��=��$����B�?� �k��	u����0�f�\�ۡƿy��w�]xѥ�k/d
���`���rSRI��t�ȃ�t��%�.֏�ml�{յ�?9%΁)��e��mE'�됞�����=�`����۳����@m��F�X\��<��?��$S��r�Q�W%��_a��]�HY,�iR�r�2=���(D sk1���,G<�՘QU(��xӌ�a:���΋bP����1��n�蹽p��*ݻi�qaAb+K�Q2��sfM=�(J$4R���	�U�'�m�c�i��a�v�ˣJ�����2�_�t�c�^y{�?���P+{��v�֡)PG&��5�;SL�ɜ� ph_é�nF��i������ ]
�x������&zd]�Y�|j�v��85F+��H��JO���pکT�k;H ��~��P ������>�ҭt����u��H��k�ڄ�t����e���48�Q[ՠ�B�Xd� M��,��\��$f���G5������ԛǪ�B���$��_���ESyP���:#k�y�=�ABR�n�u�mR�s��d�Q�"���n��ζ��;ᢟ�׵����2�u>�&������e*5qK����ء�u�F7�TXԖ(�u����\fjWםo+�Ϳ�z�Y-@�W��ϗ4aya��ST�&5�r�0�$+7l���H���t�B2RԴ�"0�#W���;s�%v��xP)
�:���Kc9���?#��V��K^���:���UV��ïj^��A����.V�=^�ɫ�Ԗ�r�щ6������&<A�Gv��g�h�kҦ����P�3�a�93�<'�6���P[8���:�y˃��������8���*"c�L:�H&��P{=�<�)�'�޳���e�%�]nAYZ�t�����O�9/��%߾
���sbgh9�X&5�f���E�z;ΰ	N`3��qr�]07V����:@o�Q�f��D@��e�[���wB�WĤ6�Ջ��6��"�h��Zغ�.Rڠ�(������
y���މ�����^� ��'��������r+x��<���@���!Ә���`/4��d�3�L �7J�ǠO�j��4=8:�G����g����cȏ��><�ێ��~����M���t���LIg@yw$���4�eݡ$�k;k��.�Vw�g�hn�U��T#���_ٹ˜ϔ�T��U�}C� ���#4
V���Â4���"�@&L�-UV5�T�aq�l~c��sϠ�xߔl�e%�7ږ��c	/}�� �o�̀f��;��N�A�J61�w���~�3F�G�c����GĹ�D�O���!��(�����eg$"���̌�B�ӳ�0Z��[�2�2Uz7!��U@��:�eBwSi�����d�Cp�XM�����*𗬦ڻ-\��T����t�$�I|�&��tώ��4c�^7M|iol����M���i��:YZl�x		� ��:n��Eh�wql�e��d�q�� �	z���ʑ7vN	܃m��3�8-���ԙn�O����b Z~Ou\��ΟP0ł9a�4�� q��`mS+O�/3^?\�"'�K���Z�^g�ݺw1���[�c�>6��ۅR�u��S�@Q��LTC8Q�M���Y�/o��.�I�o��r��oЌ��(I����t:&�kiO��é�"t"1͞�}=�P��s%R�6�4�Qł����_�DȘ�,/9���]��,A��B	9u�6��bw��U�δ���Qj�>�\i�gv�QA�h8!me�������N:� ������4�dڜZf��� �����Gn��%k���k��B@-�B�r�ŭI�9._I/p^I,p�ܴ�@&�حZSFۚӕ�a�]�Z�(�zxK�� Ӕ�(�����H�p�.�_�OA���6Wb��J�Om	�4��m��,��E��Xnֽm�ͩE��������X��%b�i�D��O�@�'v7(��4dL�[u������#�}TU[D,0��r�s��%nND?@g�q4V��A��*�m�Z9���(��҅[�-.e$Ĕ���.	>�������Џ_7�
����Q$�矂���_�zHQS��hR0_Ŵ%��z�2���W^TӲ[�Ⱥ)�6�d������SNK���XJK����޾z�U��Mh8}xg��*����B��]�p�*�Tꡐ�a��A�����1���$jy�q��R�xu��:Gz�-���0s/o=��*�9��hs��`~�O�Rr��sI M2����:�X��,��}!�W����ր&DIC~0a��H~؈��{bЅ�Ƙ"���g���S��╕���� �¬��gyU~�5�F�cLb�*z�:pbb���Y�:p�ⶫ����G}U��+[!5����vgyl��	B[G��n����}P��V�}DSg�����#Q0tI�*w���P�3/c��5^�#�U��K��c]�L/�nLª�� �e�:�FPn�y�k�	`Ύ�q}D8^b�|��>������������WmLP��ū��d��S���#�ڬ��3�΋=���+��qL��7�a�fi�?[��:�Q0��x����:qf���Jߜ��~�?�Gi�������u\U{���[��Z�����?B걵��Y�@`Ϙ�"Ȋ�\�{��W�3l���H!�U��f.���^���ѪDd��#�Q&#Aow�� �s�������pmPdp�)�S�8Q�Cn�ϷJ�3�>���$�1�`�'^9�I_nyK��AM|�fQ[J��	~�u��]�S	�	�'7��8b��$yO���jP��{i��p+��4��ޕfJ�� �`��$�[�qI�J^H�������+S�}6:/*��_��er+���k�A��8������|�*��Q�q�}7!K�&zVH�J��kh�r�%�EE!�!C�PGF�EY(�a�������vW��Ԟ��e�)�#Y����j=��TSş�E�Yc�Lu���B�C��(�$��y�|����$�$�PD�}p��Kؘ�h�v�ҷ*_������4Hc�[VN6�<��
���!��i�
�YU�w��9��U����H�t콐�s�`*��S���"j�N�����^H���ѴVl�\�;�M!=����ۄ,g�X
?͆��3e�	z��	�f�f��P+gtɶ�]Ӹ�&�x�����L̡bA]�}�W}���2JgIJz�6R��v�x\��w^&A{I��;��kM���%����H*��2|����%2[�K����Ԕ�GL�'-V@�H��}sf%�Ĕ�Y�@E=10���y�!��s��/��}$\�����S�����{כd��=b ��0�"��w��1�v���ْ���(<�oX�n�L�.YK��l�6�ڑ B_=ԝ7�_@@/�~HG�>�������e��"��ĸ�|��=L���}�u :�Ƴ\ܲ|̒=nŘ���[��=r��u!`�|6���2���.mu�%�g��]+#�<eQ]���1b+iV�b](����q����n*�}!灞��p\����,JK���\�:o��^_y�˷��c<SW��e�W)���>�����ǎC�&a;f�ΛW*�D���4}�e��ɪG0�)Y�er��#�W��������\�e��jȀ0/~WɅ���2��9!A<[�����xuG�� �+G����l�����"e"�J(�*�9�]'`��-Nܻ�t{F\% ���T-�<)���;˻����ү�СA lV� r��Ⱦ���#��n%6M�Q�V����ت�GY�z�t8��fJ�>p��|O��x���Gc��^/ߚ(!뾞���N��Ϧ���8��^��h�I��T���4\PF(��j�P�o��F��O���2�����G�+��i��	1�=��n�"�0��e��y������V�@J용�
�����6�\raZ,$���F��y���+ {��yr܋(��W^��;� X�Gx���%��T�+4�_l�j6M���ψ��M��hط��8��D%a��{�scd'��a����[��x��h3W�:�הD�.�Գ�⁶� IT���� ��ۇK_�J��U�twAxJ~5��!��.+����_	��\�����@ ���D%Ʀӂew�B��{��F<� \��3�_�йC���}��	M��bZ$a:��8�Y��ƅ�a�[*�_�Lv����F��#?k � �8�̒=P�l@�2�V�N=�V��,��{@o���:W�U��b����+���Qlu΢T�=P��Cv����S�.�$g�@� ��}C�Ƌ�����>ǃ�?����������[�/���D��`�v���a��,Qi��*o�J
��M��E
?�B�%3�T[@���e�=Z���eW	X������Ă�T-S�gZ�&d�\�])E���J�Wx<������Xɲ�F-��2,�}�m]�(&vX�=�*{<:���o���!~�F��F��i ��{|��#Y��{�2W�_��L����%���6��,W{/�i�ws�
^[,��5rv�~l5-����ԅ^U��G&=&�m�7=��Z}Y�~i��\�,������+c��iXL��"(��2i	�L������D�̵��{�V��S,yum"_A@b�[�ʛV�I�1v]$[X��[<EE�e(�x9�o�z.��.c��s�2FZ�4��*�?R!��w��	I�#_�����h��|�6��62V�s����9N���Q�߼�p"�t#�*����񴤭�`_�6X-�WŊ�
O�`�r����!̹HbR��0'�h�͹�4p�o�y�M����MBEy�҆=Ĕ٧����� �gM�^��5׎
1�;&,d�;����.$s��_I\Q�OvI.��a4����	<@CT�&n@���k漛F" ;��s�&�x�׏�!t%��c�e�A.���p�,����~D��-��Mu���S�1V��4��	$�?zj��Sm�s�t��`5��_[߼ja���b)}N�jZ��{��?X��;>J�0����[�T9�V���d���bU�ff�� ��m���1�����LctH{Y����g�l_����n�O�=�ss��6�I.�C�2�������[3��-ٝ����*Ǉ��3���[�O��+؟��ޠ<�`9�J��*f�+&��$���C����^�']�w�srt����a������%�i��>�`���Ei�l� �+ĩi��B�Tc��Z���P��\xq��;^�VG����f��_�T�Q�g�/s@��S���Ì�H=$e�7S=�z�t�����I?���x3
Y���V�,`��d�Ij����3[�	�9�c0��+��yÃ�GǕf��E�F�@��mG?qE&?�y��
�bS©�ao-��\���*r �{FGI>���O:5�?�<J5lo�rP�Y�B�3GG���-�~�����\2��R��t4(���Ԯ�vh�B8�l�1xE2d|)1J�|3���$T��u�Lq*�N�5�ڳ�.�E�eT�lS�-Zòd^��]���E�UġF�[u�����m<|b�-��H�0aI�:�m�:��B�������������UU*	�Q�f�(H9�GC}��a[��v<��p��v��5� �w%8��ф
Y��'���c3җ�Ť� ��_ 8�n)��i��\#t:����0'摌�o�6b��^7ϸ��=aT
j[ʿ f*���o���ٺ�\���!�w{���[Q���uO|p��C���0ef�hA�ϒ,cT"��Jo�9Y֕;錾.]Aɭ�����
�yV��]Tԃ��<F:��ٕ�Zߨ�j�8�=�B_UH[9�hY?�xs�1��#���2_|��He��Ԏl�zX�*�-�S\�9U���J��X�P�u4�d����_eA�
�B������@8W<(�X�	o�u{��?p�y�74DD8$���;��z�L1ٻ����,v ~���ɽd2�I�sfe/7n=����h�7�2�u'뽨���q� �c�!L����'C�E���zl[���b3P�Ie<tXu��,L�����?�t܅XS�izrO�M�-�ޣ]��26��@2�F:��`��_��9�c�^U&���i<K�|Y���{�e��+�pG����_A�خ����$����T�#�ѪD�j��;�ћ��Y��h����ԓ/��L��{Z��Po
!���}��r�@��
���p�Ѧ��N��YOC��c���E���"֬���7�c��:����`c��#�.F�I\c���Azqs�ao���Կ<�B2�si���`�3��
�V�.o�"�xJs_�[�朚˾`e0MBj�c$JF�j䥪�*?@�^M/kj�l;�ǀ�"�����۰+qi�
#��Y���oZ���|�}׈O��Z��z}�~���A��¤��Ï��=��>�r6� V�M�	�7�G�v��^�����)�_�3��
��e�q�m c�7�ل8<��l����2��m}�T��Ț'��#��2v9 l�V��q[��W$�|g�c��×�����s�y[���Ω��;�����;e�B����1��=��~oP��N/�M�Q�Q �������JŦ�E�C��t:�̖��Zٹ���?H�5k!�k�1��L'��^w���RT�Vg��� �78��$�B +3�W[��j?
^����Ѫ��йIZ\,��s��6��_���H3ۧ��o�c{����@��]<�����Ͱ)��[x�`� `�i��ـ�֥D�K;�����ԧ�:��7�n���Y�D9;�퍨[NiA91m�R�8���xV��o�G�|{P�n�Խ�}T`�����k���Bl�6�^n���Q� ?���:�0YP[{��?�R�.j�яޭ	��*��ߕ�QN��
H�I�sƮ	�W�ެy�p=/�E��$�P�<�ba�/�������9S�@̸�<�Ƞ؃'R��y*v�/� �6�(5q�f|Bm7���Å�.��5sS�{��+ӿc�pݦ��AQt=�e;��YE+���kU��aބ�Q.aXć|���d-1Ji�ZB���".�[~b4g�0�@,34�%C]M���2�/����tgnkͯW�ZbbK�ҜpFda�#�P,��g2@>��N���R|�sb8Տ{\���富3����7�o�����eGJyt���'J�s������Cab���2@�,����V}��`�0���ك��AC�Ք����n�����@���J�cU�2��Z<��ߦd1 �>�S�cpc*��ִq?k�z�٣��+�W�]-�����!�f�>>�h�珃�9�٫8doԚ�䕶���|���跶_MC��j�C!�քV�0���~�3e0��@�773&��N�=+�*J|�����y>K��V}s���VG��x%���_�?O�5��'jN�;��q��E�B��˽
��z���-��
���.HB�� �m�:l;N3bi�����I�k��=�2/U��%$�}��7��7�YPXb���l�An��2)=<���ٌ7ue����]��	����|ˎ��,ܾa�c=�  �$���W�>ߺ���6zp|�����5R���؊;�y���9� �a�֑��?R���.��B���vъ�e�RY������bڴDH���ߖ���R�)��m�Ǳ���M&������ʒ���E}�-�㌣��l�`�����ƾ���m�j��օ6�_��:�G�����Z���PD55��/uC4Pۂ�I8�`�+�^8Y��<l7j��,��}�'P.��z� NX��ʇ�$�w
rX�����
�H��
^;�gA� Џ����R���N�u9B�L��V�G7��$}�ud��u>�
�{d�I�`�7�4+&�{�Ӟ0�k�j�ݭ
V|����n�ڲ=�Χ
A�1�{7tn���ۇhH��à��̔�	[z�H7�:��|��D� b%[C����DhӃ��矩�lbN:�Te��(O�z� �h��S傡s9�*�,)��ބ�i{?��|p�(�as5�Í	�Cx��"��o ����t�곍��|�-a�i3�������ȹSМ��«���b�� ��E��m{"Rb�'0���Y��ʻ�2�h�o��I��U��B�v>g��U$c�qN�XC�tS�k���|�5<y��E�[n.y�0Zh��X� �Ds2R���A�,#��D�	����l;�k��[g@u�H1E��q_pF���\��B�y�F����m;���f�س���L���|q�-���v��!/Ѹ�1��f���#�����÷�"�j�;�S��'��x���'X��F�p�v����`�܇
$8�3&��_zl��I&��+0����g�#G3s�
�!2�+H���B�Y�@Z@����h2����EMb��g8Di)u�	� G���va��d�	��hՋ��h>��a��TW��z�9�VccG��Y���9q��uk�y�q���%��+;O�wA,
��=�`��66^�{6�؄�8�D>��
���\b�$Nr9�E��:�W�"�%v�A�����ZX0���/�����㨁*�	�K�ɟw%���ܧ6�����M���y>~�Όh�v|���Rݿ~��'�:���l�����*�9p�k���6����aj97[ t�"i˜Yg��dR	�iV��")�]!�ޱia�(�2��\oncaB�1@��wÛj�nJe���H�::v�����y�5�G�����f~���� ���F�^�i�t3�#u���n0?MS<���%��Z�2�r���5�D��� zU]����m�N��ru+DͰ<����_&��R0(R�#��I�ާ�v�a-���v��rk�H���v�T�F4/K DdQ�D}�y�����Z��64�*�)�u� ���|��/���b��\�vzB�H+�a�"�Y�!S���􌀃ѳ+V�Pu$S�̧��Q����h'	m�pQY[�^�� |�Kt�#Ƣz�����u���&�k��n-���9]�4Bp���i�A~Ȉ׾9mJ��c��Fd���F4���`��nj2!s�r�[��ʉ����dl�+C�K�9�l��d��DI�+0��f>t��l4�8h���F>��	�wÛ�w��k���uh0��jt��$e"��r��9g
�}��l�'�jJS���*>e��t `�A��kԶm?���AWT���g�N7�ΏK+X�2�@e_�Uq	���N����0w��3S��(?Otq���9�uE�e�&�Y�򝉪@=�&�*�>�p���;�x뿢� 6��%�p�8�i�S4��
�	��|C��:Df�eL#�R˩OG��]���LB���dR�B����&�  �A�)�]L_�3��a�xj�"kԠ�U%O��mz��ԇUF��q�r`�CO��࠭�����`O�W��a��Yl�N�\z�f�����:�~��Oc'⸂���Jg��D/�H��Uv�^9�Z���-�1���T�V!�]���;ll9gS�O˻�,^��ʛ�l�QpS��4���\�%v�/�G���p,*�EGHkj���"o^�fg��?��N=����0�������UE�O�K�őh((��7I��5�������9�,�\p6+��D�����>���XPy�@mv�G�'��:�c���m�n4�}����Kh����������\��ʳ�r�R�۸�4��9��?��׃i��nt�E-zܙW��Lgb�-��b8�]Dס���m�6��{ڄ鴾{�) �_�����ќ�g����u;���1���b_�W�T��B��X�W�C�i�:����y2�ҶRv�|��:!���M��+ЛR��C�}��q��o�T��0��3�'�w�)2M8��'�b���_K�4��O�nܜ�&V�)�-Y>�<[�d��4�M�\)c5�r� �\u5��9�0����E&�m�8�3�k�~(j���!��hI.�i�N5����|@.~f�R��3���w�~�<ä�"��xmhP;@�����XU��W��mǩ�t=)E������U�;�Q%�x�8��mk���d�Ѹ����pv~� ���i���, �L�tУ�s}��L���9��Pc.�+���oy���h�p��3�\�Zk�D�=f��t��7��׮�� *��+sA�F�=�K?mp��}g����ܪpc��dE�v�ќ�8$s5|Y�q�tMg�#9����o~�T��"/��������Z�8�rn���n�Lq*�����<Ba�f�=}G� 96&�շ����C}R�t��5M2�Kha�O��N͸�l�l���a-�w����@�#��ݯ��+@��z����fB�9�n]��U�M���k4m/{����%����rXl��ͅ)F!pv��W��I���`O@�^�l4u,��l���=��䝮ȧ-��Ng	�l-�%F�%%ƛ����&�K��(���I$����R��v& dJcŽ��麛�U��}��~���x�I[�N4���I�$
6Fǭ`]Jzr݈�:�aϐ��1��nh��ǂCdK�ʡ�5�-�Ј'�C���0#>�U�
��:�d��p����wL��*LAx	�O�^R�IZ�����*Ca�=[�*[�[�W��������i���k+߂XU��DC)�sTSÛk8��%A�4��Iuˣ��έ��l�
�A�g���X�?��R�T$������ ���)�N�>�0UЮ�	o���s����L�f����c	({�V�C��`�h Ɓ���AL<d���|�7�'���r�
���g��?��}�mjS+$:xZ�B-�b�]c˩���m�fј�
�a��9�礐�y���v��Q�˰���h���{78�)�.>�������BT�@���/	� � mW�_�z�� 5y K����G�A�Dg9�U�8Sw �S�6���(�#/�,k���|^8��.���Ӆ��&�Rf����[d9����i��:B��@�;iD1�ꜚ�O����)�_P*�jy�������BɁ٤2�ޯ@�0����J��M�t�|rK�c�w�t���=�Z�`%c���%��?��:׿5�S�N�L-�E=!d1��å�������g��sx�� Ѡc���G�V.�<��8�w���{�hZ����菵����w����ס��%]�z�1�i�5����Pڛ����M���A��7��^���B<t�s���:a�;�R'�e��8`y(`��y��A�V#�P�*�	�w�J���j��NukZ���`W�?b��"oGOE}=�(�BP���NY�=����/'+s��>�0H���q�ڂ�䂯��r{#ݟ��}�D�WL��������(m�A�-<���5)�U|��N������|tᜂ�N`���i�x�!�S�e����,2�yl�0v,E������.��[Z��X�s��7n�Dq�Υ�K*w%����>���"grLu�Cb_ ��w�K�B�6#�0���|���"nz�	�)e�O��|�5{_v�zǅ&�*kC]}�?�0���u�֖L��άڭ���$���������Ꚋ>B6Q�L:V/lZ��}�]��
����������myq��KPC!�T��;��ru��`�1�N��so����F^�b�|�)�!"���v@����"RZS�t|=���I������2�^}z'�#�խAʫ���^;�$��	����S�^ӻt	�u6a7i(�xC�<K؝8l~E��f2�����3�yoL	I1�2�-s����ؕ\?�U��I�1�HE�$�o=����h<���$�c�\T�	�Oa��Aݠ�%��ח�h���S��I�.�k�^t�8��N�o{����-��@���"�i�z�����.���Gm稈p,�W�+��g���;����@�)�M/e�)�x�/�Acm��!ʷ�L��o�K��kk�,��*��F)�����js�<�½�\-�p�'�@i@���a�|'���*Dh�ɂw8�����}M~8�Q��l������ ���=���0{<Ri����� ��Qd�QlE�?k%���ʨhv��.z�w�$�ˎ�K��z�j_6A�����F���"W
`z����fXb|)���[����p�\���A���,�pz �L#<1�瘽��'6ĕͶ*9��H�_�ZI����	�,	0�M��<�I��k"2Hj��w��8x��	 �+%q�^G��v �<�xH�(>�=�0A�$��݈\d��rM��I�L��l`n9ӓޓ���_=�+��|�/Do� ú�.j�>�#�p�����A�׃|!����ѥ�Vf��3�p�@�p������"�����'���!�f���[�~��Ub��%�/^�)���n^������o�{S�����A�p�ջC�@|
��;et�����Z��!��}�CB
wa*ZDv\�v�W�dϥ�c�������Q�]�V�����-��v�)����F7�[W:�^��JXX�6�3g�3<�R�&"#-T:u�����i���41Em
�W�ℷBD�P�v��5�|`��p-f���ٍ��!~�+��v��nCbe���.{��5����e�˞Z�[#ne;���il�� �u�oq�r�e���C�b�ҍ:VZ���oQ�_�8.<��n�t���B����T(Ķ�H�dk?�[K�O�\J���K"ړ�d>z6���H���0����D���c��,ք�f��)�W>֎�'���R�\����.�`P_��T��yX""�W��-P��N��rG��]jVr5�0Ԧ�Ҋ ���x�Z�����v�ģ$�@��Ns���G�z��O�1P%_�י��ퟞ�2@�����n�m'޽d��"#<fI�a�[˾��2L�8X������!�h�k�S�4�3�0t��J��{�>8������'L+n�d�Ҍ���+��F���7��M�cb�*�E�[�qj[.�P�j�G�m�Lm6��j,'e�Ĭ<�G.Q<J{c�Z2���MDk�7��܂����@ɢ~S����t �t����A*$a{�j�� i:�xWj������'��oM�VxxN�|3!�i�7��%��t4�N���Z
W�튻�x���ԥWqac2xR���W����d�<�vɹ��s���)�^�}ob��<��4�Nkv��5�
o}X����\����A�B�(�:PzjŇ�ԫ~�Z�W��6�N�٪g��#en�:3�vn�<X���R����ٶZx�	�����Q��{�¸����_�hGd�A��uU�~1��w�@!��S�v�*��f��]���lEI����\������u����xQ�KwȘ���ﳟS�R��ͭ<������3(���jn�}��t�_�|^��粉����8?��4%;�>m�����]LT�l�j��z�9;]͎��|j
�Z�
k�X�5BE��!��U$�شB4���j�P�ʸ̣>�7�2N0�H�/I8:��QֈY�t'ܯ���p^�9-N�Ǔ�ڷ3f�O��3_�g�	9�d�s�spz]�>��K���j�9qJ�[Jbz��Bÿ���C5�X�	�,���RL����+� �����e�3���'�RT�E%C���d\o���8��$b�1�.WbK��[�%q�J�uSE܉�;8���v� ��#BM������k��h��.�S7�4�E�+%�
i��l��-�)��g�a��;����E@-�7h�97#T=T4��IjC�E'b�f��a�E�ʍ$x�2����.�F�������GvN��5�<�m����5�a�R4��[�V��G9��#k\5���ٍ
V��V������3dH���T����<����  iD<�m�9�|��	�<�(����?�{�bK[r-�����ѧ$�G���$��w�KD�}�Vmh�Re��
o�{�Bw���R��N�Ƭu�P+��4�!�Pʪ�m`�JZbda!��¡��_(��2�I���,�`�BEygk��i���� �]�����&�E�&B�z{�Ձ�6��{ Ky��"�?`��X�q��#��"���h��`������`�C:*+^����04WR Z��`(w�K�~��e8r_��
�$�m�Si���=��
�� ����;�ฑݻ^@�>�9��?qV�'AO��1���Opfx�{}c���fY2Sq���?�G�}�D��B�"���B:�tC���x_�f�|`�ã�o�o�z%�z.� [D=ݻ�\z�">����{�Q�KٿV�C����^iJ����.�;d7�E{���S�]����l�|V �E��n�AA���Q��	+�6ո�J�\���޵Kc�`��c�,���H���!sf,!Ź4��J�5��߬��5�%:G�T��%�L��Q�G�<E�[��:��Ĝ��wj�R`�O3�)<Um͠��z�^
逸ݨ��㷧;[�H���
_ХWr�O�#-#S,?��'�V��`�!�Di��-�<���ߊY֎7���nw��u��-mE!wn�=����xN�T�U3��ةnI[��\�]�R���+���t!�hg~%�`�kq����-��1�C\�U]{0��>�����|� �g%�������;�I3=�߾�#��.�)R��#[��#.�:!�GخG��X��MyP�
�_���)U ��h���7V�hл�F���D=Y�Vw��E�P~n9�)�ܝ��"X�؆/�a���x���M=���{�Z��Z�!�~|�q'���V\;��R|�A4/�pý�$��#��a3��r��Ij+���;:p�T�Q�ٛ
��,���0��:UX4n�M��������d"�3��74��$ ku�����:�Bņq=B7�G���;O��oZˀ<�'`}4����O�݃�Gr7�'����Q�Ad��'��A�=�A�D�دNz�Vd��7>��E���!�An�x�3��b_�K�q����˜�umX�����Q���Zڰ�M����/:��a%F��d�����-5d��������M2, �'t��՚���,�\i�;j�[T��=� ��t8�Ėt��M�*2��mfM��%	:�(�)�|�l�:X��鍔Q(�i�}h��mopq�ϣ����Hcw�f����y'��ȟ��-#�g��7��d���ʩ �������L��n�s.�[��+H]I�̶k��OҰ�0�Q�������l��kW��Kd0)J}vઌp�f��,�DG5�Φ��zmt����H�N1+����آ�z&K(�����B��r�л���:�2�&?m3�U��j�׵2�44��\�y���-�{0�"%�=a9d��P��n�n��{q����I2x�fc��ב��-H$,7I8�Nյ)���q�e=��~ ��X���>$P�����7@�P�ԧ�N�����H��ؔ[��Q�6�Z��݉�ǃ����驸C�ʄ�`��0f�Ό$U�]UV+���fx����ʪ�X�k^����hMbC��7�t����U�zi]0g��5"��y_SL�_�km��R7�W�Q��cط�'���ݣ&>�"_���=�/�V&���N���W@�U�`�H��OЮ*�`݋p5 R!������:ط��O?��ݮL~����$y�=ObP/ʘ��X���K�Fw��=Ϭr/%��Qt�v���y��M�nz�9s��p��xst�P;����dN�3��/�M$IHڹom���O8�:Y�G�=U�XS��>ٰ��5�м���e��֎�tjF�!��࿺C�Z-�X�s�
�_�ȉ,vS���M1�G���0e-�]w�J(~���B�r����� �z��(�	�n�В�\2��X��ȕ@�7�zI��e�0ft���Թl�0Q���.������nͧ$�椣>>Qa6{t�@o����_֓G�ؿN>��*kd&ɹFЮ��0�k{!�P�{]�=T7�m��;%�DE�+t�q�?���0�߫+���*��&�7̅ݷ�>v�AY�ͻ�
����rE�H����K���z}���C���G2�	`�ņ�Z���C#�Fu��gN�H�
�~j���1�L�2t$���F�C�{�pLγf��Ƚ��w�jAU�
c>�|+__�|�/?{�Hf��(�F�G��x?��0+:�Q�TZ	)=��Jx�=x3�Y��E��P��Di�z�;�x�Ǭ1g
�NI�Y�֐i�G��� �����8����O ^�f�b�'6p+,����Q�A�U,j�D�8,"Z�SC�=�S9w� �>[ɧ`L�g��q�JR�&������	S���a+I0iQ�[~�v>�HU���5�r�ws��ĝ���N�G��2z���O-�<�I"p޼w��i+c߮>��%l1�A oʵ��6A���IO�BE*���k�zQ��{n��c7F�,X4q|���Z�����Tj��W����O�����ybhy37��N�F��x����H��Jb�0�zm�s�?������� ����w<���N<u����ȻET�Z[��'�n!�3B�K��9�]~߰V��B���؎a:D(�Ð�x�ׇ�\ہ�>������#����x���sSnz�xQ�'�ٌ==݁�������^ξ�����B,_�Q�c��}���7׹j7s �(qZh88b=ց@vk5�B�3�=��_vi��x+#���)��%�3Ãqpe��J�2�2|X*�+�UIX;7QX�>d3ŵv벺�'L]�>E=M>��+tT}�� _~��pE޿r��8�;c��|���Ĺ ��2��d{�kvK+�FA���x�d\�lӎw�)D��q$8xtu�FO�H����J����۲�� %����W�@c*錩�=p���V:zv����	-�Vp�t��)}#;6#��@ꋱ)
�x�;���l�?�,�XOpZw��ԍJM���;2"���'�ڈv1ξ�Ր���3�o�����E��ߔ..H ��޻��2�������1���R����g�[3�ɻo�D
���+��i����5*T�h|Eʲ:�z<z��P/�2��dLٲ?)�f�^T�-c�&Szq�_�v�0/�*Sò��s�*tj�W�#�&>/Ǽ���3��1�I�w+���!<����>i!�	�u�l�NRo�P�D��GPQp ���Ֆ˦�'>6�d�{��M ��P�Sg��~���9ߡ���O�N���/|6�	��v����`��~�N�T�4@@5H�/�%2�Ĩ��`��, �'Xt���)�ל�,�H��~�|۰�"/�-���bn���w�*~���f�ph�ށ�� uu��И� IoC?�]��\��D��b���F����;k�<4�eWWĦI����֯Erϒu}p)�N-[ԫ�=��tp@H�{<��_��Ք��eF�A2[�|���f-�����R'%qL67]��jڶc��LY$�1�ƭ6d, u$D;�����o>p'y?�X��H��1$*�j���ӥ,�~a� �	i�_L�T��l|���=ߙ�J�0���	L�cc��(2�J�H2�Ns������b2!"��#m�UY�u��I��I�����o��)��9�65r-�j�H�d��{]�DC��Vn�x���*����j��Ov�S�ō[j�� ��X������MiM�Q� ���@PDU����o�ة��"<�R���Ы<Ѽ���O8b���Zl�r��<[���N�nR���
Vy�L#��/���{�v3�ޗH��L���N��L)�$��h���}�]�u�V�����w�"�J�ȟ�@�TI��C�C��xAc�k�#�A��aO�{Me%��"���98��GtB
��f��5�`���gW�0���#�i�,(A�Wմs�q�=�x�@�'��96����囜�Z�l���T<^Y�7m��! |�aG����!��W���
Y5㋆nk�� {\��nUB6	�؍w�nb�� >9��&��'�Ke�Ӌ!�Acp�� ��z���#?@�X_��#U<�L���;y�/��F&5	Q��4����b�.XAxBc1��0q��|���|:�L��<�D�  �)0���k
߭���[y�o�rkl�3�r�=���dqi�#n��ã��~�����C��� ����KC�Xy�Y]A5�6C����r�|`=*�M�F���
vӅs�9�h�������=��-���؛��e+;�����1e��i�c3T���A�}�(�q�W�p��`�<�Ck��Y~�����J[�f�XY{�S�9����0%���Z@�����k��s~?�$u՘��B�IF�tD{75/j��!6qw7�%η>�p6P�v��H������� ���iC۠W���B)�xw���%b�������F��v�^K#ڶ�vۅ�&"��Vj�\�k�-���Z�GҀ��#����|h��\�CN��-�F��\�D�bQ�$YwfX�2eM�>�^k]�y�a��ZKX�
w�M}r�aٵU/H!a��-r!��ɩ�I*�TL�Y�m#�\%��(���6��=H�� �zk��S=�QxDCq"`����Ö]��B���`~<��q�DJ&#�x��=K�)���7p��'*��9�ҬW7�����DR�9q7ȁ1H�)3���~+9��'.�8'�ëvE�d�S[�p�qa��<{���`)���^g���~�3|x�~�,*����k]$c:!��$UL�
����q!��X����c��!9`��B��[��MO�q�u��|��4칌�	�V�{�=�j:�����ߤgt�VB�ً�|rW�����I?�h��Hg�ψ�Iq
�Б�h`�F9�6A� Om1�/%��L��X#��L�R�Tb���&���0�u���>��1�\"C���xz���	������K,����X��bV�\��	�����]st�A�_�/(d~�=���,�i���^`"�I2B�U@4\���g��!�`aܥ}���@�H4�����~��U��ɮ�1�{��S�㪗��ҡ���=fH�4�k�%��t����!*�� jz>����**�
"P�s�b�i��tNlj�{x���A��.������`�0%:l5	mb���O����F@%٩����������O����"N������ΔV�a�Ɏ�_H�;�iW8z�]
��959+�ł��e��|�J���R��v���#
[[�c$!������T�p��V|Y���'�}l��4�(,I�b�>-�[���ȡ9���KV~Kz�ԣ ���XQ�������L�y�� �x~^�_m��h\\����d��4c�l�6&
G,j�f-��˛=v��-2m$����E���1�i�AX��U��m�Ы�V�=Al����[K� 4�0�"��g�'.�}y��T�3%�-L@T�i'K+�V��x���"���mkm��T�e�-��xwD���'�C��Tʥ~Y�H��{�H��5v�)޷W�ԌɃ~����s�Ѕ�^ψ
�`�(X.�B�R�	E@S]���sCD�j)S���=:k]��M��q�7$:��~��P�qulɮ������@�	.�-�TbY�I�g�x�8�"�t�%���4_�d>��c��r�>�N��̏<�k0��0�AZ��B�p�%��7������E����@�K����S�IN�<ٴa��%~z�`}�)M[s�,Yb1�����=�8Dt���0����+�%4%od���m!%���&>�_��8���_��u� ��A�)�|暏��#m4 ͷd8�toK{�Dr�����
$gpP��Ah?�FJ�DH?�|d'���~�!��2r��F�8˧"���rR�ϯ����]aY���C��&�3�U����L�� w�x\^�d���.o9*�Rp�qZ..P%PS�����>�A\b�U���p?��)��F��,]�N�4H����i��������'�����B�����]":yR��E�j�ڔsDb��I����B+o!��9��zC�	p�V�(��4~FF٥��(��^��q��_'׆��N\��bhS���]ƺ�����mq�S��zۓ�W���N����e��蚏UU���)������ n���ܼb���	�[���D�����òO����Xǌ�f�&"�Z2'V0���0�2�G΂/�6��[&TX :O��F`32�HC�|�BA6� :�g�+��Tg�.���@8㲑�����s.ἐp)�ߢHʯ�VFޜ	�2��10������E��9����k{���h�F?󝗩��*Y�w����;��bg�|`Qh�cʢ ��i�L�U�5�tp�6��4�_�8�����=I\�_61�cv<K~%�ԋ���	[vh�^�C��4����r���Y��{���
�����)��#Sw��Ͽl_�0�1�П���ʖM m�Ty����p%��ج"]?1��̝±콢�5z�_O��+���,����	g��2f����&$:��(z/��Z���mai�3������q�(ŎS�����d)ա���ZB�N�VI�a����[B�Ez�I�{#֜�YL��ِ( x2��%~<�?2襶����B��¸�G�U�x����i)����1�_+�N�^�@D'a�KkWbfxA-��zkma��zԙ7RMB���$V`w*��ڶ�1k8�IT���Y�P�=�G���&�,�Ld�ʂ!P�@=�K4<�`�$ �ٺd�t0X.iP��뇟���R꾠Zg�t�m�X��^�(�E&J�r�����`"�0�f�,1�������i��IEP�W�ϋ���V�0�<�]}sȤ��,�x���n8,��&��,�,��p"��x�67F���܆���F�&4xBd���5ˉ)Q�(��j�z��%�Gik�$=m�S�)&f�vh���I�E�5�0pЁ�Pe�c��u�>)u��.!_z�f��wn���>�3n�n��=	��h�߂rT��#�j�|J>=D]���0 hE�}���HYT}*	Rڞ�*c�Xź�e���$��`R�1���)��%�����7�l��U��J���씩���lX�#xy��4�q��N��y�0L�g@k*�9�hE�1�ǖ�ї=�6h�S�u=J8�Ř2��`C�fuNe�(�W�m��48�}�9JO5�.wSl�J{����*�.N����ZE�n���8����+.�f���+�H�~�K^���4���O���s��M2K"��M�̐M��^�����݀j�ї�U�Zb��IH^�}q�@�|�^ S�?	������r��_Q"���IdvN��T>L�O�;����*�γ���4���E�{3da-O�]@̩�	\N�Xl�3w��_.b�[_I�}*=�}Ug�f$`.]�*��4��T2�d�#����(l��Pc�m�R-��r(#�A^7�0v�B�J�3I�%��.ά@�3N���;_�!h�h1:�Fyf��:b6ozzp�C⫺�͋Ͱ����R����Nv%4Ur���_j��:���7=��ĩ��I M.�	����Q���n/�2uS����q�����eHp	2Y��,z��b����H�����`�e��T9�G>Z�ZTx�����4s	�w!5��qS�!����Zo�{~8�� ���گ���VO��9a��EBVL�� ���'�2��E]E��_J/�mz�#)�/Gup�q�17�ei&qZ@����Gr�iмjܜY��{��E�ٍ�'�K��KC�/���xB�5^��"m 7��+�ܻ�u[�
�UN�����<�\˭.ɦ༮�4���qt�׿��"�����u��Ųj�1]	q�X�����-I4*���b�����ƻ=
!ƑC�f��:;&����RzӚ�5Lކ?ݝ�h1�N��9C��S��,�֗�8@�v�A�����!.!�{��0����ߦ�e�>.�orJ%�^�����p|� ,J��S�̂:��}ӈ̉;��j��mE�vt@G*�#nG�����Fx(�Su}C� 
/PP!���q�[;�g�ڜ�Ϊ��U�VG L�lZ�B.�K�+�W�(=;S�/z��Űm,��O.'oѢQi{7G)�ˡ1`�%�;�r�P޲sp��i��i���~���������aNL�&$���3����<�-�wV6O�,������dt2���E�$ �H>A��ea�KZ�"���K����ݢ5S�a3 �0>Ѫ�K�%�q���&jU3�m���-lr�tEů�����j
C�'��'�7t���'F^u<�4������,�\�X�H"]���tq�
�T�ٮ=e隵��D�.t|�|qx/#9�Z!��-��w�c�{��#�c����_�����	b����f(�tUV�^b��r��Ѕ�=�jf��,['v�sRqص�P��y��a�kD>�3"^�f-��=���G������D�͵G�PrqT�	@8�֌u����era�w@��N�쯽%���|�)RIǕ �Q(�KWHo s�Hj�p���Bq��,�%zŝ��[�b�:�Ȕ��--yV������.O�ѯ�>��^7��R�
?�*B��
�O.-ͦHX!����c��"k�~iHf9�3��\/�����@��\|}�<�ށ��l>	5.6k�D����QT$2��t?�����-F�*��.�jA�������c����v�2nz�#�U;��Q���C�oK��;�xG&��F�;�Y�bP�����9 �0�F[RZb1B�!$ܦ)	��Ӏ�0�w\4��}����ⱆV��&��K�T��pX������5�+)~$,��)i��!��OI+3Ӷ�l�{�ӓ�41,.H6���|E­e;4��^�a=@������K���uK��l��Rv�L�j�T�7�g�|u7�Oq=l_,]��������H�;)���;g��
r�?<���OR�ҋ^��P���HD"/\�ǑZ��ƁgBH$m�!
��T��3O�n�b����T��D�o59#���!ǇC�iHf	cbo�q�>�C�?��!�)^��8�-�Q�fI�f�$Z������y<�B0�SK['�nT3��㔫QFV4^��pL)I��+��׽�)�\.��V�;�$�F�+vu�%�	�_)�R[(
f���~��7Ϸg���ww,�'X(2w6	�eT�>��k.a4!eI�t��c�9fЎ��rM���E򜁙לϼI�bg��f����S��4�eSFK`�j,rtI�4��I9��D���&Q�����2Ϸ��70N�Z�ʰ�ZU4�������'�hNL�
���苸}�Ŭ�[�2�#y�O������}wK�UO�cw�����8J��k2oT����� �O�Ev
X��N`�ك�
�'�w���`�d1�=G@sB�%w���U�J�si�����E���	��s4�K��6��h�(`� e]֤��������@*qj�ҋ�QѮD^�)�gG~��x��d���Ohb�]��ym%�?W%`���3�wX.�B F4?t����b��o���`5�^��PB-����x�:^��{Y��Wc �s5I��_�D��o[��ӝPt-���)�Y�uɈΘb�!5����C�B�٭!ss�m쏑<g�����Y��g���u���x�����Z�0��D��Sm��������Z�ЀY`ꜚ�������h"�)�L�ⴅ߃���LuSaA��=�O�����)����� �O�T��0��&[mIf�*�jT���ow��-�Z5M��^!�W���`@�����+�V����k��[Y���-� ���6BjEe�jOp�#ݞa�2����^���({�8}�����-8����$V޶���7�2�m9�����3�V��]�#�u?��:�X�X��_&��kqɻh>�J(~~�CC���T��IWf+��n��L��p͛l���Z�,/�e��	�:�y��S@@4W:Y۩�*�c埓#%#���R��m%��w�x�K�q��PN��5FM�����4���T��SZ9���U���n�SlΜ��Ez:���.��";Fdb�KNz��85Z�+`x���x�n]P�:�.���&�ڰ���Ϧ����z�~���^��H�l;ڕ�볆��y�7d6�CT<N.R|s0�������z
fԳv>�í�d)��4�?�G�q���&�_@nVn7OY{��|4�kP�=��0�4�]L���/��[�����|���:JЯG�� -upo^?�
Zަ��-���/����>���֜�O��r<�w��p>��8
%��y��YG%Tt����Ѷ�)�1�/M:�r��?��/�1iY�U�����0�=U����ʚv����@�Fe�ӟ�ڦ���D�qPͷG��9,Wܜ��ȡ�HwG��3IHޓ�;���i����QuX	s3�ǣ ���'����AV;SFm�4h ���=���D,"�Cؤ�&c�t!�m�˵W�;CԷ�j�6�~f�&��C1媱�t֌x���w恳W�!��H�4�~��?Q�`Ǒ]���87��H��k~�:Wa��4P��^0��� B�l0�d)�o���Yo���ԥxC|���-�}7�����Y��J�.��i|ic!�ɥNd��W"+��_�1�{E�`���a�yાQ��F3T�5�϶��%\�dNI	ȼ���\h����*�͊�iA&���AG��;�)��_��擄|j��9}K�L�e�t�Ѓ��6E�q�C0�Y���~�˷n8��S3kfN���{34�K�������'AT���Âʁ�jPL���O�S[ ��)ſ�[p�k*���̦�D+xЇ
u�/�Y>�K�P�0�x��QL���;��y̃Z�߮Ѫ[��h��o@lbb��أ�Bc#��w�N���L/Ý3�F�w������eS?@\+��7���z B�sئw�ЦqI�x�R�MѺ�k��}v[���<�=<�O�؆�8lB�}���Е����]맟���8\�	����T3
�\p�xA�;�FE�ƃ� }��_�M�$���qS��K��ET���s�:[r�',NG���X�pi�ǚ=�j�C�'���-�����(wx �&�ŋZRXg��Qf�@RTR� ���Hc������hҩ�>�b��K��yz�����a�%��w�|�pa��:�`�2�
8����b��êў�\��-�0��§h�Q� �x�(��ea��gqK�<T�[JH;[T�]"�3n��V,�K������Y$�I2���p�̛L�Šq�ʌ�� ���f��cV�v���B�YI�w5��O%�8ks�L`��Ͳ{d�y.���.� [{�b)�˽��G��v>$��.�k�D�p"��O�~�A�]����=yV���\��ka�Ԫ4^�4"'J����Z7�H�'�T8vB����h,��&�EV�;��U���h�4�Ӹ�8�8QW�ŵ�}yY�e������t�׊,w��)KCH�fh(��;�����e��B1�D�a����,v�3ݼ�+�n�.r�b�&)��`_��=�]1���m��B,F3P�!���(�6҆,O��z���`���P~�H�8�-����� �,�R_�K�
C` 7o�� �g�����zǙ�\��8)�ūyZ���@Ť�����ǹA|k}zN.vV(��s��2����d#G��t��nL�s�)`u��]�+	:�6=�a�g��H���1�\����G�ڣ9%�5�4�fM�h�ػ�k@b�ġ��]3�b��x�]�}��qbӒNly�F��7�v�պa(
%��%	nC����[}�*��4X�"Lcp�����$�?*�5���_�?-�mh��H
����ڇ��>Z�C5�`�${���:���n��q�*��Y�E̋�R�P��kW@Z�������i�����1,m���W�ݖ�ƪ��J��^]����>���R*3"T|�UHv�vL�����tf�|Q�a� p��^�у_-�<��D�#�U]�����{�B�֭�u���>�!�����`T�q�L�N��R�ސB����ȕ�,!�ԯMsu��|?U��|�\�
��c�Bv
�qP3��I�r�2ZKC>ˮڠ6wi,��6�N�� |�v�x~ �ͳ[�6dY�ry^I��+���(�8%�LW28�1c�LŪ�Q��.���[��T֟F�L,�t7?'�U�s��-��l|�w��{��)x��`�����{�?rF���~7`�����|xF�r�����9�YlU�w(�;�9���^e�MLqn��k���T���w0��Ë�8�̄d_�R��w��m�0���N�M���Xc'�F�[Ho�\p��JqM��&� `x���v�J�HA��[Y���3�uR_5U'�3�P��Ӂm#�©��w2�A�`d��(���6�w�.�0!����K����x/٨��l�Q�z��C:l�%���(ֿ���>�.ܭB\Z�����܋����G�p;�-Xm����.���ߐ�D��A˼c�o���6h\�/퍐���,����TV�`o���5K�t<�t���V}'\}����3:"�|�!�2��n����&	��8�O͵�s-�o��Z9lhc�o��l9�߁qq��T����s����>$#�=1f
�dޒ� �����wd��U���h`{rM�& ���z�e�N���t��a��`SJ��:;�E���5pMG:]����T��g0�#H0  ��v
��1=�$b(��c5��6n�{����IGPx~:����[��ft��������3��D#���=��,��@�	��.(
,A3W��c��w�v@K>`�"����z-0���V�0�cq�]�s��'�;j��K?K�qh�D%R {�%]��kY��t���q�'�^�� M/�_�BӶ�a�|�ͣ�⡉;z`�X�L�O};���+EHv�$��G�����9���&ּ<�GF% I�z ��6��x�y7`���"IZ6h��󗫄� �h*vK�d���r4yb��6�l��~����,�+���e�*I���P)2�7��CI����D5��\G��Z��p�>̋2��eH����@^��Z��W�΄*&�t����й���q�"�>�8uMj��w���!D��7`Ѱj��Y(R�_���&��e$�D�MG<���aE�����ʪ]'�rՠ=�*P��T!��#�~3:�E����K�h���FJ\dA��K�L֯)!A�%�o��$i����_)�ꘃ��:r��Mm��(���t�zA_�B��� �� 㧊3-�FK^���l�(��Jd�@d6�+AT�FB��%�M�*�yP�t�-L�;��S�t|3��=��UCV+5f�@G�O/�r��$rg����kxm���s�d����=��,ٲ�� �$�%��������:�Y�a5�V��<S�)Z�g,hv7{�/9���7P�(�R�A��J�+�Ɨ^[מ��\�R?�ʇU���lC����ܞS��z�T5��U}2z�~:�8�/����ԧ�,�����pB�F"R0I��n����S�R��Y��>�T9ֳU���e�$K| �.e��N"��d�/�f��詇�� �<�1d�
���x�rh��6�D��J����Ǿ������Ԉ@�f�CcL������͟$|e;���HHEhj��w���Cy(M>�gp)�
�;OM���z�0���Q���!� �uK㔿$*OA���mx���쬪��X��ݜdj�fV���n�x���W��5�A�\��ޜ&�r���]Y	��6%��<�M�����IAx�=�|��K��L_ ���$�͵��A���=.�\�J��{`�/?w,�B�L"?�}=I��f�D+�S1(~H�@���d��3"���۷�K�G해ʮ���ᲔL��|�M�����mz�;L�l�(�<��eW��;�.7(�?�|���P���a����+�6��n^]�G����]���!JL���D�C'�(�Z� �=�T_L
�ahЄ����xB��50Bph�q��Q	Muq�lޑ=�Q�������ɕ���s5�
���s� F� ��-3ݞvk��M��̖{J��`������1|�ɔ.=THK3����hV=ɫ�����e@W�#�>m��_� V3iSko��y	�D#(����s�$�,�xK���쎜Hz��Fi����.�~�����m���B�>�����~�x�'�e쩺q�L��$J�)w�"[Y��%�����:�����u_�G:>�ʳ�f�ђ���m�Ё�b��#��;IF��F�	�&�@�Bm��/n�, AfTEY�q��i�
�!�F�'_�{@�_�E�l�ݒ�R�]ּV�{!ync�Q63�D�L({�zb��V$���xI��L8u���3��o�ކ����kZ�qD#xSG�� ���F�m�Ͱ���N���뒛MEƇ_��y��WB?�i��<���k2h�)c� 	rw�xS��wx�g�ޜ���j(�o��w���?js�p�m��@�Y�e�� Qsh����6�������#��XɚX��0��Ɖ��|��xt�����BY@�?パ}�w��H\eROb'j^�sB�n6G�[�,&���S�t�� �Z;M����������/�����lp��d�n��㐦�RP� ��2<@8CQ��aS=��e @s��E���iHp��5ΩnFf
��;�N')G��U���,�mCo�0=����;m��%pglƘ��moY�kc��
��)��9�*��-Oĳ��8l�����t�4"�R�6w����eO�N�OG�8��3:�yU^��7�߉B��|�h|x�|_z�"�F��Q����*�>�F^�L�|���2^LJō���o �B�`)��-s!ۄ�(����u
NA���iϽAӾ-0բ��F3�홀b��V6RIħ���N�m	Y�r���A�m�EQZ���``_,R� ͰC_Pf]1�r�+�헕�)�R��6�l��c�RDtt�grU&��;RT�y�O ����^�)◠*�xBtŻ�5#jP�^�M�� ���;�<8 �`��|/aVS����?��!�Md����1�@"��9J+���%/��~#�2�v��PϹ��ݝ��칁����\�̥���Y\��햞�>#�7W���<KR�d��x��Lc��0hg�#
��^��e�y���uÒʭj5��'���N�@ �uW]��`�h/����Z?��o/�S ]���]E�.D3������k�#�������̡��,�L��+�d�9ٮ�&E��w���|�ݗB��)�k��ٓI�f��#!j���j�G�8xϟޭ:�����#�%4�K�~�9ռqa[����\>�!��*X�.(�h=�LYD��r.�����AI���������n��<�V��~rG��IxL&b BK-�OML�i�ή��>���h�(��g�|8U��Q� R�e ����1l%��J#�!m�*�E?PG�.�_��<L�ke�^@���c��}�g06-y�,!�4�'m?Ub\�R~|�Gt��%�[%�
g�PͅRc�8'*ʤp6{n��O�G+r��yFހ���]���NȈ�sz]ꖮ��w��ǉ���0漥����f+�Y���_�T���b�[׆����s����9�eᗨ�!���w��<\��Ga��?8�->ݨ��0SJ�=�Gn$~������k��'&� p�B9�O^�&���V �|���,�gr?nJ�2�Q��
�?�f��=�%)�>0�ml�hc�1FI=��.h̛��D��W�å��ߣ�-�Ē�١>���^�����\'���&�y�����Ǜ��� ?j�p��9�=�i�[�%�%xJ<��o �N�]��!�v]s��AK����L��k`�]��E6��XY��E��4R�������ܢc�}����-]�[$s^Y����LWǁ�%b��������*�i�r�C���3@��zՓ�e!/ul��c�_��أ~F[�|��I�M}#y���D��) P���6^����K{�^*�E���a�>-�Q�O��T2���W/3tH���e����bf �Y��0N�=�Z�����d��r"_@���0b��\�a[ߖ�e���
�MΩ�qAu �� ��߹R�cs~e���@.p��ĳsS�$�y�1�ɾ�M���F*�{�`d�99QƤf�ܛBx!�$}�%<[��+�t���d�ӥ�->,%z}ָ�2��%�P�+w[���Z�W��mg����_O ���9N��|�J8ע�j�	���}��9!����%Ǣ�Ԇetf��<��6�G����=�u�	��q漴�A��O��_Pڀ�M����g �9��I!1�I�b=�tg;>H	�Dy��wrρf�i�=�`/D�R=�9�&�g��	,��t�ӣ��Y���1��)r�o���B������X,�:�w�5o<�}�`���j�;���;P�aWIs��»��M���g�'BOz��1�_s:{�>���Bb�&0�!�����'ۤ���(�4���`�%qG�{*�*O��6���}����@��Ol}�r3�'�~S���B-���N����\�5aQ�<[t��!|��.ɠ�����wr��B��O#���"{g����;g�I��ZŒ�+N�g��-ΛK��m�Siۉ;1�uN|�� ��͸��b��_�;��;a�>� ��zǟMwB-��]�E޼!��G.u鎣�����4"�dn*�@�v-��2���S�H����`�z7<0*5�4��$�#���q����}~�+(�`�bqp~��c`��2]��'�$ �'H-�HO��.����
B�@�@�S �f����ޙ���y�BC� �EZ�U)P@Q��:c�m^�)����`�����O���(5o`rS�'�I�U�jJ׏�U�[����`�{)�mn�����>k���ݢ�Q�g�xOԩ>͜�`�YlXJ�:�v�g'uW@t�c���nB�[ЍO����5?>�B�{nː����d�g������3��Q��<�~4v�O�J{�&x� �3���E����m?,���L�V��R�F>���`��a�A���[��D=��`�9�� $�y�q�Y�6� &���rO��t��0��j`ĉ���R�����e�~Ð`{�FzPd�����OHK\}�ON?�\�sT������U�5��;]��/��W-y����z�0W��1g��+��cA�$��~h�Zs��g�dv�I�%��c�v����ߊAҼ���4���+ͩ	�{�E��=x4��1;07q@�yk^��)�h��ğ���f�E�wC��$.�=X�C�Ʉ����3�Eg�!�ma����w�f����m����_�g�W���V�az
��J�T�<*��I� �Mk/�LFl��.�p$w�)�A}�a������*xkE@$!M�e �,�>uG
��7XҸ����5l�'7AABE�v>|&Ѱ;PD��ߗ/���<�Ьؖ��pNbz�u�$�h�a�H	A_/`�u�ܕإ�F���N�{Y�0�@Z�Y��V���f2�e��m�*��y>�n)J�n1���pO���� �^X
 ��In���%j�1�*�����g�����4��×/^*�q;�S��Q܁]�&8��ƻ�il5� ���K[�b�D�h�N���Y���?<6'�fO�1fN ��|��9+���� ��.v�.���U��Z�S���Y�-�P���m(e�\�vr8��D��	
��+��b�/G :=��������A��^�"��'�H#�2���v*�\�<#nK}��X�_��?��;��G�"���;U�����8
5j�k�H���Nzy��J��L"��1}��?XA��MG�@@�/c��4������7�Ů�-V6��#�+i't�&��[�g�A���i28X�*Ȩ�(� �O~2�㋄�&�+�����'8�t�&��g.��4��=�֖��9m��al����zm�_��jwE��c���Ct�KS�Z���W���s���*��\�lu)=@�&�A�QN���R��ԥh������.L�u�/u��VN{�E�%G�Q�p�'�-�Glz���"�+��y��R���������n��ժ�|���!'���\���<�M�sx5�P�^*���Ęb�z��6L�V�Ʀ^�N%Z�XCO|Jo���>>G�xy����\�)o��2<���$��TgZ礿�x��S� C\qͲ&=Q��b��m5 � o�����E�_j��Fr#)[^�[��	��yK�AR�@2�F�=��Tfe�4�i�����ڝ�(�EA3����)`$?7�'�u�D.]ю���Fs��Iv?��F�3dO*Df�e+��zd¤N�K��K��lqϐ��oc��g�SXxx���f �c{ų�_�NƘ�re�k`T�� =�Űa�ŕ��W.<)�����6PR����\[�r�*ҹNʊ!�3^g��S����
�)5`�B��W��Z� �2�g�o�)�%��OÈn��3ǻN��a]��	.�׺Q�=(��"7����K�a�=�,�8�E�S���Bm]�Yvj�P0t������~hy�^R�⮤e�0HG6q�vcw �Ę����~ߢTq^�g��!��8���^� �F�9t~��.Ph�3v�����#Ο��	�!��s��7�N��\I ��s '	��64���Z��>��VIJ��lZ�M�0�q_�?�t�>}��f0'a�0�tod�ɮ0�ц�I�e�ִzC�=Z	Ů6��2v���D�I[�֣��58��n�c�������Yy���֌߄�6���7fb8Nf��<l�jR�	��rC�Fzʁ�h����
�QK	�eRA� ;6G�����Eږ;��\p�F���w�%N�,�d�А ��{}���_�XX�}���X�s��O���ʃ��n�y�1SBv�QÐ�.�~� �L�ζ�d�&��A�N�x�ׂ�s�$@g��%���Y��ޔi�9�#�\]����(�cj)��R&,�����vY����9��n���ua�ƿ�?a�a)���zȤ�IT�SX�a��v���nKh=k��,x���]Ղ=(a�*��={QU��vH�v�D$����L��75���W*��x�H��	?�n��ˬ-�K���P�8�u�������R���f]{T��<8���f�FD�%2ӌ�l]vȼ����6�Rۋ��l��b�Ʒ����뗊}�޿�M��c��E����N�Rh	��/�<B+g��y�#̭H��yJ�󨆖��/���V/ĸk2�������p���ᧉ�F�4A��r�3M>��3������w.�p���������('��YGn��~����*�y�`��h���J�xuSW���B��Jt W$P�'��������H_�!j��n�n�;F�{<#����d�~I�l�
�w��*_��kn:���Bo�(�ϱ&w��V2@�J��D_&>���8��M��os���>|p�C��Q�?w���W����~�n8(����ݖ�AɄ>���Z&R�gC�P]1�	Tw�˜�OG�P��}d9�9Oy����\�^���N����3(�6��MI8��=ȳ�����3����a&�
犴��Sġ��ⷆ�tpk6�j6��7L�nL��)���K����j�X7e-1:����gk(xm6�Ccd�c8e^L>�d#鳶��R���Yd�>��r���d-�͜��O1`�d��O�pﭘ��lW<b���O>�U�]u*}(�|��s~ͻ.��K-�44��愾��j��0���vzÔ�"�]��}�X�H��J� ɺ�gbu�cUBZ�컉��h�mU�Ո��T�����*T"ӌ�׆���؃z.�Ҋ���!XW�����7դb�)V�[���<�3�F����s�@O�֝�
聵��P( �jL'h�X��Åz�~[{���9��-koH!_���L����a�S܇��Q��n�C|p��H}�U
(�3�7%��w�r��$g+~�����ZԌ���M��X��'[ ���PL@�ɝ�y�EĹU�'��ȵ� #��Z��^�(o�� f�q��HsH2�֯`����򋣩sr���j�}_@�?@+N���O��]j=�Ee.���\��ʝ���I<VI_N�,c(�s�F��('�ƍ轻:!��R��n�����Ƶ4��W��Z�6�O�L�#^iUxo�$�d5�J�t�8�X@u�a�:�ݠ�İ�QԆ@G�V"��h�}��uo��M0+�\���hj9�I}_�H˱�?�[��g%��G���Y�ё�m@E~Q��I��gw�E�n�S�e�h�TA�M�&s6��y�|���ޒaʰ��_mf�����z��U�u�]�ӝ�w[7E�������D�]|c ��+,�95��urM��B�y�_��onZ���?c�4��\á&"���?���ʛtR�k`���g?����Ƅg��G�X��:�5��ԍ�񷿚ep���,�Y� �}<'�G{⼾X�|�;�A�`�J��IK�ǥl��C�
nݑ�V�+�z�<Up-t�gW�^N6��jW�{�׼�Nh�д�uM �D�����`�&�Ө�83����V��KZ�V�$»��t��HLu���8��'�������%��������R�`i��*;1�0������ι���9հ��(1��"-e��Q'�����!�eZ������(���%ֿվ�H��~�����`��AO���͚���΅Y�Ԑ^������Ԩ��8���w{�t w���3!�܁'��MBp&km������}5\��@���e�ӣ�g�@e���9r�h��n���V�Y�Mj��ִM������zk�>�0���G'�K�)(�}�C)9̄�8j�/�wɎJnHlE1�Q���*�/q� ��	��Ԥ�0�%�oM�Y�c�2�,Y�&mu�k�~�������L��\�%�m��*3��ɳ�g��B�L�䄷*XC;>8z�ӌ'i7Q�9�Ě����MϏ����ĎWa��a��M�W�$���\���|�A/�h��b����X��#t���}�<��!T�Ҷ[��*�����N豙����3�;s�5�,j;�)�(���D�*,kw��&�p�;3퉿�|;W���Vn=KtT�S>&�R��c�8�oܹF�Kw�����n�U|#D�'y��1�9���u⻙�GaR:���z�vuLٚ���gI+�}r�`�[,P�Û��v�7�?q����6�Z�hB�<C�ɟ�'k]7���
C��X����	���p}K�*4�+tߪ4�g��3���T�w�s��iO��d��ͿF0�,1�:ˀ�#��E6�����dY��~2�����s6��
 ^�g��dɁKd
n��}m�5��0��/*���h�)fLwoONP�Kq *^Q�9`�;(e^j=Xx'uU�m�n�K���'\Ol6W����4�+�=���t�4���m���`"���(zJ� �Xr�C��i-�T��>�@8���F���"qݵGz��V�P�`K�Z�ß�`S���hԹ�݅�
��y���
���1�()k~�)�����N�����$"�0���6��0+� B��6�@�/��D�*��y�����3���!���k���Qf�QH9��&��J��/�b�c��Dc��aM���lke���)�F�Uw��Q�4���25��j:,�̨�[}��v=sM�b�Z���& �	Xݢ��,���[
�4l��0���Do��M{�>0_?��?�(+ּ��/�-���}[����l)�jT�9�_��)��v6
L�<|��gNN�O�Þ�pg�00�k�VWX�t���K�{� �0ؑ����Ho� ;��˰��f��y4�;�{�XL���$�y�o���G�����A	[�i�\"��찀w�t	ӷOn6�}��h��m����iX��O�O�
Ƣ��D:d�|��v3��IMø?"8W��mB��U���NfI*��J�M���/Z2y�'�������L\�tr�BM��U�C%��e�D����h�L�:�]��p0�
P��씶 ��v�A%���%1kB��D�Q?[��+��uܘ�ИR�ɐ6�8F]���@T�����[����i�����43��\zQ'dBRwK|�)(5zB�N=�?*�F6l҃�U���?K�T�y
�J�W	(F/ë��d��(�\�\�;�H�X�R�3����Vc��:���n�������YXoG�P���N�����_��eJ,ʻ_��K��A���Lf��'YC�c�	ax�!���*􋩸r�jߙt��-���ѸD4��$Q��q�������i�Sϖy���h��Ti�丘��?��c�cb;>��Z�#J?�ٗ��ga���z"0���e��Ln�ȧ.$�vo_�W�b�S�"	e��Lq�V�o��@;�y��qV�J�	��'0�u ŉ%ګu���j}�v{:Ȟ#b�\�4K����!	XԤ�>�N����O��7�=����f[�[!�������P��l݇��@�����L�p ���/�XP��I��D�:ډ�~~�%Q�k�}�ʧ\8`PWW~(�+(�_�����.(i�)uz��b�CEJ'�e�%��HGK��� �2_NU�n3I�/e�odtI���m�̪����1�~��k�E����e�QW01ɹ�X Ԗڪ�$�Q�l�'���E\?3H//��=�\M2��L�{1��������b6w�@��xp�����6��$�ԹRU+�����l���S��v��,�W�ɿwD�W��'Tx�K�3�Wvzm�4�ȣ�ߵ��q�s���8Nk蓙�'#(BXX'�_�/ά���ΒӉg2A�~�V��)���PU�c��K:��a[��XөSC.H�MW~�!s'(ʛh�p*�\8p.�'���F�؎�f�ٺ�^�M��l�#\boU�mng�� �>+p��^g��v��4��)pm#Č�M2�5�B�������q�5*�:i3�+(I�S���|��G=���+h\��d���d�(�ǣ�\��#��k�����Q�����K5S���%�����xZ��;v����~�5�pC0�dL$R�Ғ�?���U���`��"�oh��'�Ð���r0��ª�rFzT�f�=�����Ä��Ӵ�oD�RU�ŒN��U�|/at��!��迨rlF�D$0N�l����2/�v�rs���Lkp�B9�b�4IEx�`�B\��{�#��K3P"=���J��s�y�4�{��a���&�s��Va��Mךh���=���;A�T��S5#xU&hej*�4�$�\��xv��Ky@�ؽY��r��Q}�w�6UYh�����>D)i��	��C6���P`�t��N��a����0|�Y{(ھ�ヷ�z�o*�� "d�T��}��|�/d�
g�Kr�P�*���]&-W�����5d�k���N��Q=Aj��"��f�)�6Mhh����xҢۭ�$���������
0{�p��
�lO߸���ՑI�;�AF��c)3kr�$8֔RHvv����gx�9�Z�o�a��R�\�Ss�}�,G����-�O�Y�a�LI�7)UJ��b*�"�Z��5��L�)�8�
;����j�k;n��%J��QbY{&��%����,n	�'"MX���&y����1��k���3�)�ᛣ��:�����L���`�a|@C�n@�YgF=C�܌�]�v� ֗Oψ9��Q]a�S��?�ݏ��.�� �ol���I���Ȋ��ǡ����v��H��N�-�}.S|�P�L�3|=ůEm�i����"^�6��{(��#JTA�� ���eG��'�=#G}g�	���A/��(�ف�Y6��B1�����������|��H����D�חKm�hB���ˬ]���np�>�Xe��N�Zr�b���H����^�d�*�%�,!RCh>1���$��	�׹�9*Lut3���5_�+5k*G�1�T� �3�[}}�\.9������<jH��f�ZOw���U��0��"tY���C<E�o$xh$�|��	?%�̄��l��~��{]<>nj-�٣�ʦ��ڷk{\%:���'o�7�b�3
H�:=���'ń4�w��3���9��}+!u"\�C�?Q�3����<�XY�^B��I?�35Ki~���l~�]��5�O2�j�[,
�"�������ke�Mn�$�	�����UI(�g�DT�Sc�"w�R|6��%�,$}�$W97I����+�I��i���}�#��0��^Lw~ŝL �0t�����k�Yd�R	�/������e��6 F��_#|�4�2���9Ef0Q��a��:���_Ɣ'j����D�;���oC����z�����a�^�v�b�653&��O���G��x!�+4,�o��Yn�{�[xR�2g~8��6���\�U�]���^*�L<�$.�&�	���� 1F��P���D}����frD|doT��FMz�/N������FT_��Q��q)u<��-�9�i��ᒪ��cM<�������G��e^��)>W��jl�8��M
u��yM�t�i�>�v
(���o��c^*Э����A(q5n��$g^���.x�q,TFG��Gל��.��^PC�{���c�.v�hO�E^p���Q�:	���=T���=�0����$�Ҏ0˗0����{�v\i:�Mxh��]���4�ye�]L�G|=�R�Q��=ʝ�����2���A�\�w%�~����P@���mq�_�9�q�m�vX7�M��7pXH��a[��[�pT��$�<>�4Xj�:G��>������3g^�L��Mj-������i:����ܨ�V�!�>�dXo��fB���N�����	�1�R�r�'���y��C�Pt4�0�aR����C�)��9=-4 ��KR�S˦�+v��Q�(����:��P��H������6�e?�EC�'�*~<��������
W�)i/0Z�	�'#by��a�4_�� }<#���oL]o�)�ܓ�2�{"�ȋ���w���jBZ/-]N�[H�Lq0S�=�A�"��z�7BtJj��U9'���`+$nn�:���&y�b3}u g�
M�=?��Kl���e�$�$U���±�e�ự	���s|�r!`����@�v��X���N ��j5��,��ŘAY]1��a��+<>U��\5@���"T����0�8M�5ge��M���t�F��p/��U��V�#��S���s������H�^����:U�+ 9�_ 4��1a����ީ�i��;�b�Y�_@I2�^)$��bo��4��>J;x���2��G����?�Ҩ���$�E&�5��C(�24W�Hʒ����)WL�����O~ųϡ�'�g�]�P7j������ 	��8^�vy��rIGZ����ۅWt��<���-�p���E�GD�&Q��g7���u�l��Ļ�8yȊ�7j_i���`T�Hmt@���xveY-�L&�;��>脓uN��'�4��[6��/�D�&{Q�R���j�ħ� � �U>����_&v�eO��cU��~IB�@��������{�e_h�0w�o0�W�K�:CJ��(�^��'�<ŹfM����l��{�A�AdzM�FHmH#'����=G<�b�Ce������G=�;�Yy��%s�O$r�)Z���:�8�iBK�����9:��\�SU��)�`ѿ�ܜ�Nk��_�4���޶�!wg�?�:����@�0p����	�1���Kԋ�'�N D�f8H�yUm���67Ls�C�-q?����f :�L�T<�lD��ъ�:��:�������݇�j�}�6s��m�o�2W~`#N�Z�f��ĺa���Ȏ!Ԍ��zܜ�b��Ȟ(��Vl���v��69���~P8ɕ���?[��+��z&�8	U�J�� �zp؍¿�DSm��e'��hk�H�p���=���g�+{��&�*�v^�ζ�Ȏ8R�,���淝�B��iN�16���U�G	�+���@	l����b�S�m2�
�D�}4�-��:%���F1oG�jt?je�A��n��r�#�b�4��hX�R�h��Dp�3�	��Ä�H,\����}�����҉����m�R^��B�]qS	�Έ&dN���[�*+��xD~8ΪՄ�Ѧ~��ej)��VcF|��??�\ql(�����:0�����`��?�Юb�"#no��v�E�r���^s��(�̢ϵ�Bs�U{?{�J��-��I�����S���r*���>V8��V�1���by>��RnT9�m�N��uE��
xsU�$nf8��饟�[FF"y�O�P�n�6SDqM�2[_���$X�TO�ȳy�/4��z����&�k9�z�W��
"Z��Yr-�+�ԍ�,�T��!bvb*�N��}K7O-~���a��2"��Z�E�m!�v�	��'�U��ɚ������|[�îx|%yv_Q�
	7�xJ���&����zfB��E��1;��>��oLNu��L��S�����\w�"LPjg"��I�ć[�̜�����_�5�GU�4$��թ�8Z�E6�*/^��: ��>�nÓ�tE�J0�����P����o���l.EJ�	�7�;�ˏ���5�՚I�Ḳz��^��]�,���ڭ����������|�Uqf��E�[X]����>OF��?n���O�v:��g/\?~S�sK Y��~k����ݻ�%�F��~�A����k�#3��B�����~��4[ۦ�C\x�����-���������S:U���x��w��P7�:��ճO�O��a�YJ�sc��-� ��`�l���{�?����5Pm��c:�HO>>��� �8�y	@^І��ڏ���ԃ\��n�6w1�4n��^Ĉ�,}=�XP�)P��*�,���̦��`��'CX`1�G�	��u�3�`VfN���̭�i<�΂���H�y͆���ŗ&�-�5��e�����d�wv�����K���)�(��ř2�}�+�4�GM�eG&Z<��D�@������:vOe_Zd�����d�͌6I_�\��\[4��b>��oL��\�
`�d҅���{n�zb7�:�8֣Byw���+�Q�&�u�t�"-)h��N7 	��g�`�SQ��"5+�+��-@��T��a�`67w�{ڪwr�b*M�N�Ǭ���_�b��E����mD#@�y+���/�ii�a����i�.��kJ��Ԫ)��a=�}�ܯ�;�$ϽhM�+�]vE��(m�5��+����.>�$B���D�)r����S���2B���w��X���P%e=�X������H4��I�������>�U��Uތ���NI�x[��T�^�ei�7^RZ��zy7�-�J��>�P��c�\��t�F)��H��G|D8[;K�����&Y��!�?l9=k"�rMr�`�fUI�G�Ķ)�'����L8�c�fs,�f�}�[�`&$A��׏�/r �7=5m�L�_����^AS ��'���:᯶�����/�w[�N�~I�:y����M�ٳˣ�� S�2oq�~X�f2!���k�@�h���Ǝ[Wҁq��A6��9�bZ_�5w)�E��I?XU1��r�aɊ# =�9�zW�h*�*����΍�(R��`�hwة|��1�X;R�d��U�>nZ�O��]��Q�9Ϫ]���f�䏣5��|��~�YQG=譗���@�5�GRT��
��7�v�6EL�]�^��_����	=~@����p�����4���'��̂�d�Qq��0Mʮ�!�*�AU͍Y���Uu�E���䦠a�T���a\ �^����!�iJ�y����=���y�Ɂ�.��.`2��IR�u�__r�X�S8�,��`�͡J�W~��I~	jr�����FKu���NDTz߅-��h���\z�>���(U�,����wkV��,����$mᏝ�!��2�6��-��ג�P��ܤ
�ޓ�Ӑ��ya� D��#���Y<�6k��IY�������qA�;��.`uV�ˉ�y6��9���0�����	�`J��2bp�I���]�5��N����"]|��:f�T���Ә>�6��t�RK5����aŔ�v��+D��>�8�������**Q�[;w�������2�$�(E�e�m�]�b�'\��͏3�� ���gg:��P�	��J^5��vT��O��/��l�{����=��Ë&Di3�	-����-�]-}��Q��ÞkO��`%��+�9�7V�"'�M�[{��x��{�M��7a�7EE��ub�	������F�y�'B��oN-�U-���!����X�j��x�$;,cW|}��#Rx|��W����n�������67hb���#
�����B�D�D%��Q#��Ai�����8A���"+�lZ���^�W�`?��
�]�rQZ���3km��RG�k�8B�Y�0�N�L���Et�:cLLJy�@�H�������/�bw��:�C�K��y§�J��?zX$�t�.{�{~�l��VTU��&`�/�q�*�P�hH'��׶��{����:6浿�a�(M!�Y�w3>�VF�W��xw��-Ww�j��Vg�r�h���(FXa2�����m�0��ǶW=Ķ��+����;|3��]Fx�ٷk���Owۨ~׎r�`Zsc�/����)OxV�;��/��ٰ���4܇�U����U�aI-��ѫ�]9�����������1�S؟��OE4�GsX|C�l;����e"&?,��b;o���;���� �u�6��V}�&��ξ0f��	�f�9��ȴ\���A��uZ\�!]\�v%�s� �����
�1�]�|�\?��ќ�%�7k��"rY՘�P��r�l�D���?���N��6+@S�8$[��ݞ���qkc�R+ɯbl�_x�ݓ�Yq��a�T���[��
�=a�/���\ZH��p��I޻�ژ�$�Ts�?����a8�ӛR��Z�S�A�-�J�|�ա�?�f�)�ږ��Aў�����/��P/��F��*��~򅗖��C�^�m�u�������z��|�x|S�gzr�.�	Rk]��s|�T`N^=h����n0�b�b3a	�������餆ⳬ��� ���#�SYӀ����_��PDުF[�
�ƺB�� �(
;��!�VY��D"Q{6�a�,5�)�nn9k��j}�K����O�	���G6�|���UY�O�M����$����|bB�Jq���e����5��)V(�^���W�O�`�f;��ՆO���q��L��I7�^�t�J�C�֡�<�{���E�a�FXKc�!���Bb��kr��ײ�X���v�wL �D�u���Zv�k.�l�2i^t>�Ch� �(� 3Ya�	O�_�x�N���u��K{>h%Qa���&��BI�>S)����vq�2���ᐴ!�oo�����1�LS񢲾��}�rd2�*ė�+�7��D�dj-*�;�,-{���d��<H�0����@����XI� jmnցuy���rMJ[i	˕W�_�(l�}+�8Xe%�5P�P��^{$|�����T�w�epUs�( �_:<�6�=���B�":-��ž2?9@�����j����w0�o0m��(�I���I?��=A�,����m���
%����Z��\,T��bxA�b��ra=�Gx$�������Ԍrȼ�a������?�-�"�d8E�IS-�<��a�J��6�/Ჷ�}�����rw����I�7*��� �<����Yj D��?yࠇ|�>n�e���Ħ��6�#u�/#�n�S�����8��>U�Ah�[��vx��-;.������e��"�
���ƾNo#�Um ϛ<�S1+.�m�=�=�)�i=:w`�IS����+-3/Pg����Ӵ�߿��&#��(�4�_�>��f {�N�a6�SACR�pWpF���6�D쭊�	���a$zY��Ɲ��_	 ���fTmM:ʭ�ZW�F��>��y�Ӭ�.��2���|�o�p�6�T�~*�M@��1/����&(ٱ;[2�������x5:~@H�Di��[���[K ��Yy�X�h�M�)��K���	�tz�,W
rk\ͬ�M��6/��F�M�!nfم��D��E+�N����a��!��p��3�]��⼺a���+�W��#"�M0t�����a��v��܀�$w0<��QO��T�aUQ$�� ��j�Ka`X��?pv�;��+=E�h�f�#�ĳUmb'�=ЙF7����x�E�JA��5uAB·-^b��*�ny��]���#$w���.o��K�3����	PcT7�`.�_ˣ���d�mk������n�;m�x��UĠ״_�oi�:3�,��}��^�M,��:3������ʠԙa���x�#�n�e��l�DW�K<*7��\�~���3�Ƀ {�$���"�ZS�ipʆl����S����*�=��0{i��i��<��=�ie�ƀ���������	�]�o�zǵ| �����%�������/"���|da��c7r��~��-rq#��5��E�m��)��bm��`p��{�Q���D��˚�s:ҷ�G��)�q�Iɢ��&��ї#�W��u_��@��=�az���?[��~j�N���0r�?��>6��D�([�s%H�ht��dV��]���H�-���E����{	���\CW�JMXR�畚��v���X�d�Fe����:�ljJ�]����=�V 8%-#�'	�F�N�s@�[�a�~����q�J�q�4/��wH�q�/��֓>)�Y�l�K�<*G���0���\g@��$�d,4� X����ψO��%v��t�E�kS�g�Op�.�wU�!恮�Ѱ :n+h��dq~�p󢄝}�# !K�$Sz�,�e�|�+��V��[��
�X���M-qD{h��Q�'SoNJ��6��Hykf��$I��m�P��/�&�w�����0�7�厀)��C�F�������˧��Ԁ݄�6/�/�����iĘ'uƐ;n��㯰3�aھB�Ղ������E�C:�C׸���D^��-��nzry��SI�8�()�r���h���K��/�p������pT�b���M7�(?EC��};��[�;3t�,#���4�kO�XD֨��u�p��UM�d�P�=�ӡ�3��6�ܿ��2V	~�_�!h�ӊ�v�㴃c�
���a5��&��k9T��5D���͸�����h)x�*w>����)M�z�S����+���FB��MI�]o|T`�ܯ�e�1���WϿZ}���~_-��t�"�-�A�8�j�d�^V+P#Z4�i_J3�*��`�;T��,��{�`�(�h|�n0����H�*&�q�5�'D0�qv��椥���UM���2M�!q%��~�Y�D�e���������*!Њ�����I�t[���de��fxո�%,E8��_��F#�_��g[��z��B".����5h����F��ݶ��`*�n���L�/�fX���e��6x�q�X��]���$�y����V�9�p,�Y,�#D��K�%s�*J6�����{�Y���3�ިU<���[^�U�'lM�Tk����ɐ]���L�����f��Ur 6GJ쓢Y{���]h��Yv�ގ.x�qx����e_�a�*{�י�Y/��6���'�d�-49�fq� FK��ч�Q�eL&s�_�?��A7y�]��`a�I��1��8@!xHy��&�P�6 摖����(Q�
�c��*�`��A��b_��N���C���F�9@*u0WqaV,|������{��L[�U�!,Fz	ͫ&�|R�۟7q�C����B*[?���StH�h��.�u?J=Wd�A2P�M�f�Qƣ*"�\�2vl���BM�U�E�\hC�lê����oLk�F��F+B�~�jޛ0-�NW����g��H�f�\���_fŵ��14�#�~�Pr� aWn���,q�+��d֚��Ti!rPl�9���Ȗ��L�&�q��W[��bM����é�w���0��Y���W/�N�屿z�T���<(6^C���%���[�Հ��$9�y��aU@����-�j�~����F�����,�BTb��a�G��3�óŐ�C���8�>@�e��n����p�|`����A��&���ӑ������Э�MMsNSЍTW��"�q|��.���� ��{����B��o��o�T����9q� ��6L�/W>�k��f=a�NF>9�	�� *"�q�BL�
`0�!D�D ��]9&���F��m}�8)� �-2�K6nx��<�Æ:��_:-x|���pn҄[ӑ��9�'e^���R)8�앗"ky�܊M�8���<�Ls<9!���ధ,�E {�[ŵ���h��/F��,���$}|��|4h�W�"�$/�v^Y��@���D�NEJX�H7%���;�:|��nOFO�!gx���s���~��#䜁���b�A��<N�nIޣj���i?��W���A�肠x��r�U�g��� y�a����w���˾Ot��	����?��s��	ysW6�9�e/��`8D�J{Mŭ����!{SeYD���x���~ ����l� Ū���2�m`�u�g���l������Yx���q�^���k��ieΎ�_ͯd�i?9O/^W-6�5�f,Q�;ȉ��L����H^'ܥ�d��1;������������Z�)�*��%g���Zρ%��j���UW�(�ψ��ߛ��ؙ�v���7B� J�v%�����﬋KG y�1L�8��߰-��
(kmgr��l+��6g�l����K7_IC�&��Co��m�{�z���Ɖ+lQ��Q��<J�$��K�.[@޲�������+H�Fy���lxNl�#�0`k����o���9����nڽ1 �gC���l�E�g�'���MD5�6�俣��Ԁ#9���"�+>�O��@*.�!v_�U�{���2�w�~J�C�݁��y^/{"���׹H�� K�%C �����M �)u�x�y)�;B;d.D>����'l� �����������a��F}:k��ǎ�Vx9��@�ӽf"�H���(]�#�z�"^u���H=!e��M}�~��ϟ��?F�GOQ��선~�1���Ɔ^r����҄�1W����u']��h�����!Z�W�E?���e"Yd�e�r+`���r�A���� �HۤAJo�����$���曤��Lg�W�{]ٯ�V��[�J^Ny�d��Y��7��F�w�)I[H�x�f� �U�N�|�-�x����4P�u���?��ʠ~ںQ�;���!��X�\�-Ż^��(�i����|��)��;6&����z<%�ܬ+�9%.X�x�vDXD���]���E���&���D�p��v�<=����j� <F��SqZ�WH�;��d�l6 Ru��� �E)�5p�.����+�!��gc~���0 �=ҘuI��!�:���T���y*8�S�H��&�ªck�o�Q�_�R�K��|�VZ�D7i���P�)kگ�q�	`{>�T��g�^�峴wm�������(ꆚ��q�z�O��{�-�����+�[ �1�.0�Ƈ�v��<��X#��ʮ�ٻ��i�\w�f�����p��y��(b>PݝLiP2`r�{�N�j����<��[�"1:j�k����'5�',�;x���oN��"?��^�G�"�?��������yg�g/�Nִa��ۂp���x�X{�R~�<�?Q� ��cV�5g\��Ħv�w��|z��V�e^��GHǔ�X����P��H�z@�V�N��}���͂�Ek��Ζ�wZ�ӄ�|�l4�LY6��fM[`���~�E����,>;�#e���.�,u�%�ᛞ�_��ŊS<<1f�8|N�rl��"��� >��<�gL��I���A䴰���>6恏�l&h=<�$k�S�JO�I�&셜�e�� vY�da�5��#�_%�Hl'ݑ$�8�Q��9~=�����L����N4�2�R��֊1��>���������9���y	q2�'�E�}C��l$:o����ޑU��%m��V1u�>�,P�<U f�;�Ë�ר\��B;��y/���q�P������'~�B�b�x	e'n 	�+�9�R��$�N��j�M�.�>U�#ug����{���"kT���(
ڨ�7���=Ho����#j�c:�AobϠ.:��oY�%�ɀ���?�/��2�m�9���Z,�q���wC1��?�����χ�%Ȁ{>�˶�{x�L��. �%���!nQ��j�a�]����y�h�r�-%�=��W���O3Z��,�F � �3��d�؇7�6��D�ڙ4Y��v|��؍��%=/�{h����$��XZ��/q�^�q��6M9���� kͼ�k�O����O��L.��5p��t\1I���j|s����;�0T���o��%#��@��]�y��l>ͧ��A���(�
�ЕiɃM���x�+]ȱ�`С5�?�г+�\�YƬ%�Dv�4+\Orz�������N�--�]����+�k�f�t��VW�h�L��a�Y?�y�1��=zk
[��T��iu��r(�=�BL���J��zCz܉�M��F�`!�2���O���=`[H��h�jp��e��q�Ů�.67�1���Đ~ꖓ{�G�K;����)/‒�*1�p�8�Y���I�a��z�Q�_��=�)�!��z#5�"y��\�F8l��΢� t�3^��P޿X���Ə��R�(�����\ ��|�f�����_��0�����J���^�����<B� ���*����G.ː��i���9A5�y'�azYX�/���������s)\gZ��b �3�]Ar�0�(嘄�ɯ���g[��9��bd�c��� �u�kD�Ƣ.
a�����4���b 0�n�7'R���R�>H?��j�dH�/P,(����m;���-�w�T�m�2��g��;B���M��'*��N�Y��L�ʛA�04�7���-8�i�ہ G��q�2��4�z���" H۝,����or�����8��CJ6	�����f�PZ���ѝ�:�p�6i��Ƌ��qn]i

P|E
��11AH������%�jU��[�@mh(�ʒ}To.�Y�}��_? -Ⱦ:y�5	L"N�ӽw�}��j����e���?�p>�')V�a��M�ݳ�=�"2f*@�1Wv�͗���̀�W�E��]��Ӥ�=^��Jր�($�R��ZOK�d��]��C�+��3�ĹeP��\��(�%��p6�p�k`���F��LP:߰>���r�5���ԊԆ�2�w9�f�D�³۽sB��l��=&�O��
��R)%&LV��Bt"*4�L%�)ٷV��Em_]��*�@�Sԟ,��1��PyQ�E_��ز��(\MR�u\m$l1r-��+�,�mqn�C<\ϲ,�s�2&�k?p|�f�xfi�N�'�I����Ůi)l�$��ۃ�����B���$4NqꛭQ���zY�)eEBp�|����r&���M�/#�r qĈ^��L�2�b5up��������s�J���SY-��܋FIy��GvP�=v�GbX������|A�#y���Q�>�L��J�"!�;l��",�쇼7*f47U�0�a������c#� '�?^��_<���&��ŵ�fm�BD�������F�h"���6�13cY�0 y]T�\��P6<kQ����E-*RCq���A5�'�O�%h���cxqd3��t*W���@��Y���;0�~���m��_A�]��:7!�O��n� �w�H6(���
��o����Κ3�#��./�@�!��	���z��а�pg�eD�+:&K��/jl%!��4=I6��auP&�ܩx�������VU��W�M�7�b��p��	�a��FU����{��Э�%���jAչJčeg��U�-0�]�I��h��2�L[6��VNW2*�4��M����a%���'P-�b���Ts�pa��J��S����d�=!#$���.�@R�xHO��|L����>�`hS����o�h�� ?-ʆzl��7�2/���eqO'�)A�c�D�]�N��'��py9g�`�ۂ�{l.��K�n�.�����]-Y�-9{�l'�S�:��;��dAN���E0i���Ge�����eW�^	K�Z��3~�I��O���&�"����jW�M)	R"e�?����F�������G:��l�S�����Vd�Jߨ,��k2�S���X��N��6[��p7�ĉ?:u4�G�=�8�5���GdpK�w[�C-(�� ��׭%���4y5w��_18�.��g�ps�EZ�u��7�T
��������7nK��xP&c����A�ݗ��e}Դl�wٵE6Ea�XW.k�p�� o_�����Ȭ�@�"�y���y���fL��R-q�/Ā��F��:S�R��b�����s����bKk����@t��� ]����[�5M�l����[1�����epQ��GR���$O?G��c�n���3n��' �Wn��I��L��i�<�~�ମ���"���`�E(�Z�[�F9GY�\�� �[���yO���ƝijP�'�M�]��Z+@�]��1�W?���a��t;>F�!-�"���R_���w��7���)�9�
tG�da��fK�P&����A�P�k>�ŨXaj�!O���ns�`x|��ҽf5?ja�a��i@dX^�J��#OY[�ج)1��o=O��!VP/Y
�RP2�L�,�jq�6��Š�d�V�yD��FoGw��@\0fB���N��sC�2%I$�q�}�!<���B�-i<8�j�,X*� '�l-�.��	2o.ZJ���7�_b��%��Ϯ�z�}B���q�>B��`��`Q�Lt*|��E!|�z(�w�F����U:(�Z�0���~U���9[5IA�����S��1�7Ox�ǝ����S�Z-�RX����m��#�PO�H8�ظ�)�w]������'6��5�u8p�F(�U	���Nd��å��C$p�o�B������i�#�X�73�q����"|���5lm���E�M3�m��]�()��[(�S��d���o�]�[
���+��o[��!<L��(��-=9�JpV��`��s��N<c�
s^(�ߵ2�����5wL$PZq�8��m��,�u��K�a�<���ĕ�pM�sI'5���u˓��A�RWП(S�����C0f`��>�����#f �3!��w˓��V�r��(�7�q�oJ�#���`@�X�M\��/�m���dV��%����U�[������z�n]�lR./I��ız��#lw���qMM� X�!�R���z���M���i{K�&��b�i��V|�Zf�i�6�d-ҍ$�@B��t��p�@&R�%��a_�	W�}zĝ�����(oJ��qU�5t5�N�b�`�W��]�ϧy��F��#�m��?�x�AiN�Y#<�:�[����ݶC�Vkp���̈́3@l6���/��s2�1�\�����}�
07�\b�}�lR�W��Xm,�O�Nv��ɤ�iJ~O�������M;��f��,0a[.	�Y����҃����H-�/:;l�Ik+�ʔP}+A�<i�$G	�a���Z�?aqM����O�=���^掔���	>ך0�8�QC��V3QD�5����^ࣧ�R�@{��Qj����4��M�*�>���|��hjy�&��7ʘS����ނI�@6[
��߿�qf��:��]{I�}"��-9�K_��[�P��+B@e�>>��\�T�ӘJO�$wg��	��94?�#9t�&�~�;�`�6+�ʁ��B�?N��f�ĨLm�W����(_�"�^��U�[u�󵅻jd�����i�P֟���{.=� 6l��ɀ�(t g�m�������*]��(�a����Aܯgk$Ec�[���!u�1����]�������e�DY��6u'�1+��~�=����;]��g�-Ҏ�P
�;"O���I��m��`���Z��%
v(�`�R��5���cz'7sX�]UU4�!��2d[jX9����z��)����<.S�C��2702ޕ��R�S��_c*~пH�o�ϴ�6]Y��ҙ�b���z�?�$�/��4�����|iA��pS�S,�L�2��������|�d��3��̨<Lg1O���T�"����&�Fp�QS|"�̍�h�Թ����2�"�<c���GW�(���p	�[�@Ī���nfEx�^:*���C��;X�*�QM�ՠ��6{rN�~��ܘ�0l0~�\E�����v�M�Z4�j��\�D���!:�~�E�V����
��.fXY���|��;R� �	y"�I���2����%�70+Ú�^��WBWZ�	�h-^!���{���W��$ڽ����N��R!{���hJ��B��B_b��e�׮�$�A�m�I7U�~���Glw�N3�N��3S� ~��JC�]SX��l#"ư0��6`�5�B_�X�$E�2�P꡹h\���(���-��~k�=]T��f��3@
մ�Z� 3�T|*~x�����(&������*��-;����5�3��XMm&�M�b�4�t*�U���u�P8�%7H/�[�KJ��`'��O����ᔵ�+���_�_g�?�J_3z\�m0Va���"���f��DD$��Bo�\XCe�d8�Wn<am���<���2*��L�e)�/�Z1��9���e��(��	ԑ!����1���{��ư"!�e}ƛ��i���s7k:�q��Ki�`/
LZB����"�Tدz�i�Oّ
}�����'��gi�z��[��2<���bȾ��U��=7G�,fF���Q��7x���r�K��7�T�2'�D����i2˿���q-��N���ڢg�������:#��^�ɇ���c����+�ZSBJb)��T��cv�qw�p�6�������S����r2	���������S��N�.ҝt@����no����-F�����ppn���Op�җ��B��MԻD�byu��M�^�]�����kD�t�`����:@+��3i<���ck)x��Ȝ1�Pt��LY�2�r�Z����J��#F���z�Y�?ޜ��
�=�z'��L>1�'�斎��~�;�~_l�6Þ�B�N�xxtʍ��Bc�M�Wς���࿗x�}��kcey��J-~���O�Wh,J� ��.��zX}L׼Gi�(]�*f�)�D�x�*���
�=C���`V�g��q��5��D��y�I�`�s����A�Y��U�2�C��V���)�(�C&���w��"�q�*���3��p�.��_e1�)�t�-�i�)gs~SGG�"�U�N�un˯���BX@/E�$*�;������'�^(��ަ���}�h�����~kb�x~�a9 z�&�]bc�|2�R��	C���T�F,)I�xNʳ#Q�ۋp-�T��	8���h���e�y �s�-�L��CODW�Cf��3%V�D'e(sOݖ:k�+��4 ����*��]���#��AN���LR���F9�vm$;L���8�:�.��F�}��9�Q<g����s;ѹ��ѿ��LrfC����;M�����'�:��>Bg�Ty�hOe�tX~�¥�}}T�u�}��N}�Y9��
���B���ƲH�k�+$@t+̚-a�o|5�|��VHL��z~�l_}���MƑ\�c,��ʝq�J��-�f�V/�
+�R��2�[���1�T�~i�b�� T�{���;�-�j���]�nP����3�3y��aJB��y\�r�*�.��F9�x#��3���v�t�a"!깂N��ܭh���O�l�F�~]l�q ���T�6�A��l��H�^o>Î�w����k� ���q�¸I�� �Y��������p��5�/��p����ۺz�$�ś��ҩY`��~_�#:��9kV�&���cz��ĸn����~.�n*B �_&�:@q����|�����1�y��B.O�n��έP�Z%����� (�G��g���*v�\��C��]�����e���%�g-���Ƞ�<d�d����E5�p�toL��hX�쓢�V�l��������%�R&.���?�A�l��b�!�H�M�p�6^X�F߯�G2�����^Jg��t��pyo�E����^k�����vm��~!#�|q_��BIm�.��[��"�m����09��[@'�J��PЕ���9YSIN;�\Zu���>�l����f .��d���m��|�Yn]�\�+ʳؼ�`�	���7�#q��Y��P�>l����;�>�ie�0n��F_&}J������=V������[�{r��,&� *w��8�'� <#���l�M3P�i�h� Yx&5�F� �+��%g�eUSl�f �3�i�F8"K���S��^�;N��h�˔��P:=�����Y��K����"��X6~���̦Oo����Br
z/�TT�PP�v��p�t����z���As8T��V��ӊ��:�9d�{��yq�ꙩ�Q�SO�^��㜛-�"�1�u�'5���	�6�<:23uU��n9�y o��,�c�V����x��+�@ҬT2A��]�������c�� ���d�,@���6�rxS�[�&��N��+���d_i�g]
4�*j���7�AZݒ}� �123��T����vùD�-BP�ݭ�{Ќ�Q��G���~+>����N�
(04&���	��o�]5l�VW`��&���$�u�z��}�+�R�6�O �o��K8R��FFǟ�e�&vE��Q��t��.RN���DU�D#"�+9m��t�����٬�����xofT���,1�[��O��z+���%�h|���g/�Б�w|��� &��	8A�#��j��Gt{�/+��"[�V��VX�~���(�	F-�e�m��>�>��-ro�/"q�	�L������n����Ük%�{���'��]�ǎb�ǰ�����	��۸��a�o����;��J���<W���]r�m�Ɗ�����˩rF�sJ%���ҔJ0i��uyi��x\p>�~��u�nG:}χW����}A��$��A�M�a���'��ā��s9��!������>iQ�0q@r_�P_�lS����3P�Ib������
�.v�oae�p*0
q��VHh@S����uҋ�^`R��`g��Q��OB_Ftw^�*�s�RD�1��­ͭL�y�)�aB�B�#���DIԅ	ϛx�bc�s�o=�C&���F�Ɓ�S���pU$6Lg|Pv.�I|�ҭ�'� \�9H�M�ɹgCE{��\|~���ol�|/���ъ��o�x̎����#�I�
�������f.r�N��5�ED��dB��r��5Yy
�͈aB�L��JǖTO<,k/���E�2v-}�67�"��-�����]iT�Y��`5�DD�r��q�:*d}����ψ�="��F�Է�(}E�=g� ��VN� g�}a�N\�Ɇ�sQv��ΪY����9ӹ����WS � �<�h�K�_#s0��#RN�,3u�<��4��P�;)�#��+;�ڗQ��B�A��)UH��M[4�ڌ�,EHCD�Y�B���ҕ�xbW,"U�M���m3_�ǡ΀�E}\�����g	66��9E�y��P��vWA�$�3	L�+���H-�`Q�t31R���m]�P[i�.�V�G�1���>��V���)l��'�ȃdt�=R���'�M�[1���򷎩�J7�3�t���=d�V��d�t����_�� ����8��*���ތwi�Y��3�N*7$1�M�<�z�C
nf��t�v��JT��0��WmdD~nFMU{����¢�g^��,�;MRq50�z�?S���������N�b�ÙC�}Bt7yЎ'L����%"�B�+��@��p��?E0��f���@�aP�T��Gv�����IMCOۃ-�K���&܃r��>���2�X���L��2V���[iN���OT	M	\2 �� ��
>�یܥ��u�U"Q�ޜ]��[���U�/����{�;���r��@��6j�:]R��T����`�/5�Z�KK'%z0�8!#�ўX��Ϧ�r�ȑe�}��
I_��*z %�n��9(�����S�X����y�D���zDĞyݍ���O�E��F0�?�k���q���E���ȚΘkR2J��$�m
;��}Z��`g�a��*;���\t9���܆�/J}�la��[�DdS)BG��p�?��
����Dm�~�HR�C��4�Ma
�/>�Td#���hT���M��bO,����z^ �2�q�'YR�Z�)�N������_K�� �o�R��o�P��}[���4���e&�llgW:�@1�qI����Q�sXK�X<����_���prw���^Q� _�����.d���k��̆��mG�b1iфH
�(���ER�>݂�=(���\'�����g3�m��y���2�"ӓ�"��w�.����ʹ�nN}����� ���.;�x�ԓi`�E��?4��*��]zE=їͦ�}�XX����2?����V0����\D��ZЀ�r츫}Ua�t]F�W�!��=1"�:��n)���]}c�]��������G �� @#_avW�_lL6���ǐ�"�A���S�w�9$���� J��p?������N��Ӥ�}���Sq#^Ѐ��q���$�?}�a�D�y���|���_���V������M���ky���`�DG$��]��<�`�s�ŕnϱ���﮾S���T{�C�)o[V����N��҅����D����K�C���$�TO�L'm�:���S���<1��a� �$J��٬@G'C�Dߖj�������-�U�U��C'�Xd���K��Z�λ��$�oY+�#����8m��Q�|�.�����[�)!���ι:��>w<�9�H�?v�N�Hj�A&�Q(�ٳwYɘd�5�\��z7�����A!.��(Ý���B����Ȱ�r�t8N;��CuG�o@��`����Q�z�虏���9c${(m��t^�L��7A:o '��t���W��$��]�Dǖ�T2�̹J܂~���k�O��P�y�3�!�}�Ҍ��S�j�%�0}�}B�����)���Q"�d�	��mGM�3��H�,Ă���\O��΢��u6#��O���=�k�����JSC����a�+#>I$2��4�͞�<z|�r���jh�JH���t����M�˔Ec��Ԑ7�&�r|H>ֈJ1����3-��ƮQ�&
Q�����C�9u��������m���#�w�O[1-��\�¤��2�3�CfPrbͰ薧��ٷߐy��Ux�큩�OIz��߼2��ڻ����~�m�i'�J�s#7��
[g|�y�~C:��:!�iVNq�����"�@61fk�ym�	���L�f����\� �,?����T�/�A*�Ê� � ��b�������?�	oU@�b�FE��y��\^��-��%l�?��بYG�ۿi�N�R�\1`�Z-��?�������/ǝc��()mR� ���>����:����� ����f"�Ӷt�e�7��
!�n�L��GK���C!�$�����ƕ�e�k�G�"�ߩ}�(�We�Z!�՛�� ��ZCL>EM,c9�Vyo���;�|PQ�|Oڿo\���Q�lc~�"�4`���@N8��|���u^�/�F�r�4�"w7��IH
����b��X"\���\�v����9D �r�#cQ,��Ν��nd�ǜw�S��+ ��ч�(d�WZ�)�9���!K�ݪ	�UKs4R��nF�]���%�����L�Z�}Dc�v�>p�x!4E{�|X�jݢ�*H��"d]�,�mU�;^g8�p�钮-��%זv:y|�r� ��g�c��'�+�(CY��!;Wc�u)6�O�?s��KQ>�bC)��&ɵ���L��w�v�'mBl?M<��J�O%��X�aM�A؁؍��Ɵag�M$X��(�]Z a�o��y�j6s�g����dO�{� f׹,,l�����,s<Naj��}MLA#�l������Β���,��+�}��].Y��G��s��5]�5�Ci���nNQ�@~1��7LZb�XO��j�g��a�B��t�#���
�{֗p.kpԆ��s�Z5	���u�������v͜(9/��hW�9[��͗+󰎻}�a��Z�A4Oݕ�D�.���^_���wL�4w�
�� #n|�ne��`y�y�LL� RN[!B�I-�"��U�pn^�Up�_���Il0���ł9�E�e�+~���ք��%(@lH�~��f�٩�j���A�����O*J�t����6n���f�=y�YB]jհ�
�<T]g�K���X�SͶb����<�1?��i��t��w�'��[F��~���7�U�!^�b������T{
����9
�?⦔�bm�17;H��y}��*���	ŗ�Tc��n,�Ǳ��e[��8�U� o�a
`��}�U;H��&뒣ė�|O�:B�?���W��W/.�b���tor���צ�W�c�pKjx��ɹ�ŵ�����̵����7�OWoFX2����{t"^��L��'
]���ݍ�H�/f�A��^�k�3����Ƨ�(�M0ad�|����9r�뾉�R8|q������y`�Ė�p����֎��w�Qe�+η.�35��o|ήW�u�W<Y����4��O������������9#6��L]����V�.�x��#T!���j���[	e`9q8��P�,�[B�|PW�m�B�o�1�4n�r	㤸j��^��h$�mz&���F�/��8!nU�/=AVH+��/9q�����Z	�|X�׎Y�"�óYL��4��]O���<I�4ҋ�>|>b�O&�v��)͋
ׇ��	�E�Wxn̜x�64��u���L�4�h3;�1�Ǚl��7=Vgy�Pd�o���L��ߪ��ƫ�ח<�ݓ&�#s�A����Q*/�.-|��2��K!���݇��'�o���.��]���h>��t6b���U�v�6&pW@� s�@��.�(k޺P8M⅏!�4x�am;&$U$F'�;�}�*0��E�}���3�/cc��!�dg�<5��MD9ƅ��z�}�Z�?�zR^y@ȁ?B7�4�D�,g��:Ja'� J1�b��ò�c��@���H�};c��R@�|"α�r�E��)�F���k4�b���96vp�5�kT��8��V�T�}9۩ }!�y*wsX�NXM��!���)��Δ���p@i^�L�|�xhY��n�lx��ъ@Z�H9�T��T&R�����?OC��r*\�Q��>�f8�7�<�Sĝ#i2/Ժ3��	A,/�ٽ�U�8��-J�I��}]|����AkK
\p�{����9�hExFhW��-@M	S�c;�o�7�ɧ��-��u��Gk�X���M.Aw�s�@��l���^p���1�,\f�R�����9@�32yݲ��~v��vsa#D���k\K��"�e�B'���������S��L�c?�BJ%����N�AL���aE�������*F�0�ZK�c�]rzd@h(��Α!�3\��k���ɭ*�E�[�F� V��w����2Ѝu�I��"i+2j����BBǠ�@x��8��]T�H��ij������a!��U�O�+/�_�J�R����	�guI�֣��mяu�	Nr.�.,���������B:aw ;_ �='R !��/�����[�
�؄�0���+����G�61=�iVsb;�=;;��8��Ļ�S�
�8ʆq(�6��H�H5���If���58�p#_�.M��nW�U��KL�D���;l���i+��
;UM|�K�)L7���(`���7�u*�����gC��_�>|���3�nI�)BΏv��'/Y�m��[y�����`��� 1t�U��n��SsZ��0	�^n� \��`]�DO��o�nч���H*��G������kݣ���2�ܫV&�]l��Ci��%�c�HD�}��šAt���;�}��ҖBGHh��EO��)� ���x*p�=�(��1-R\���Sߍ޹DQ?��`;#�{���
Mnz�!h<�t/~�v5�����I-lq����}V�f��{�� ,�qB��sw���q���w�b(+���Hc.��e0��=!DRgtP�GjM��c�A�Tq�� ��<Y�5�u4�m����(�x�Iʏ�q[ˑ�I�@��QP��)�IpHWCZ��᱾5�m6+�NI!��4����t����� &5��hT	�T�s��ľ~�S[���	�%,�C\�s;��hݟ �91�ٕ���眠�"j��n���䬱����p'���ۮ��F����!]Uv���[�^�1�|a��Y�`O��ġĘA�pc���ѧ�������g�U����
�!�8�M7Y�����*�D)������`�:��?ߩ����6"$��UW��}貢]��Sb���Qmw��5OQ>"��R9�ּ�A��TT���6h,^��Ba�$�?X����H�8�"y�GM���Ѯz+$AZ���T��\�	�h���>g+�`�?���P� F�h�$yǳ2<�I�v����,�r�H��`�ւ�vZP9����B��E���H`Q��ncx�O_���?�j���������p��	B'\���y��㨯��gh���P�&x�����
���Ռ�_�-búﾰ��u+]��U��fZT�Y� 8��#�0RL�wž�[Zӊ���C8�O`F%v�������#�wm�W�=��R1�?���������ad8�+��s�1��bЛ���E�F�6��)��`�mx'N���W�4��-��1r?��ʉ/�mؐ�u픾=��Hz��Պ+E��TW���p�{n��"76r�sk�)�WkfIw��D���~�9��g䫜�-�!�A�eu��ej��\�)�t����D�p�Φ�ӉI�?�5x���RT���\�"��e�4�Uc�6�mU�}<�
������C%S-�D��<4��#��itגDG)����a*�h��	���n:�'�ԭ0Q��O?����\%t�YK*,�k<�߄���*ߪ���V���_�j��"�n%��h������F��̄<�����hG��U�oɝ�!!��k~�bGj��΍���S���<��	�x �X�6� ��(_�v��Dt�?�
�U�Q�fAT X-/0d�K���-��3zw��L�b,/�$&@�Y�Ѫ"�;|*f����U6�y]�ɻ̑���U"O��iZ$C��Ǫ��(z�q��%B��r,�y�o`-_���D��G�m?e1��UJ�@&�<��7��|��4HV���i��`7a��6/zk9 �'y0�d��QզB���~�����j�+��|1"ן�
��a�+��2n5�<��� �a����/ �4��a,��ѽI1�����7ǋW,����Hq�s�H��hk:C<T}o?0��t�'��%qEf�O���:5����)�vR���~P���2ǰ�U����72��O��x�����>���
D�4���Tw��+ݭU�I��b���	�n��f��U�x+�J"&ZL^�E����)O���EX�7��@YΛ�ikC�8�:L��=�ұ�e��Q��0�/�4�'ꤻ�\l�G{��k3|9N��{��T96X&��UH��F�6�����=���p?���9�{���g,�W���� �.P68ḀN�L�d����^ʈ���f�DTr-��rg���I�8@�Od���-��s�&��`ʍyu��e$UM7��[^1㉔�ǆ�9c�'�a�>��)�0�J϶
c9>��R���C6t�����&�E���a�Ҟ���Q@}�#��w��M@v�W����ʭ6�N��|-�5�2�Jli��@GK�a�(=K�΋!nʎ,9}�ᰶ%v�a��cwbi�ۘ���Z$};�m�H�D��SF��EAh]/���W�]�&�\+Y٧���6�~6����� �IK�H���6����"�^�y;����~�_+:[���V/)��õ�r+]�Tq=SO��tv+���q����$j9�&�=i�򨦂2=ö�)5n\��9�3�?��3��nëM�H�&�򦯥{Mx4�P�O�5�(FK.��WȶS3�@�|0���l�#4ZH�4)%|����/=$rb� ���=���������MT�L�|pa6��}~�<z����XT�qaN~-M}b"?q(�hp;<��lp������oH�냮[����Xn3:���<��փ�V�#�x�^�\�F����{ ��Ū���ۗh!Nݽ>V0�GkuΦ��0FP�nR{�c=�-�3l��9�
�����ݱ���<�m�%8��~�p"�.m�tj�m:w`�l���0<pX�А��;Y�JH���켼�������9]��7�Ag�ޠq�H	��Cξp=4�������f���:�ʰ�%7��p_��^Ļ5��^L�[X�؝���4�lR�6%C��x��x�c����?gC��ZpTT�7"-E K��ba�kL���7���b4-\`X4�د�������k
��C�V� c����d���/z�X㭷؟x2X�$��>_���n7߈�F��C{9��_U���K�f��%�R=��-���#$���gH������r}Cn_*]h�EZ_�0@bdQ��ѯX�I�@��X����=��`��\���i�Dĩ��>c�=\�2�//Fũ������<}7J���S �J&�?�	$f34�h�j4֜|/�P��]��2���7Wt��=j�/F<�*!I�م[Ac���ܓ}V�2đrG8���٩^"D4�dN�vN�U9�?#Ŀ! O�4���d-<�ӳ�1Mܲ48NiI`�p���+�2J�ɢ�ٮ�+�D�e���oO�Wpݿ��Ij%��oŀY�H��*���"�W���#s�C뽞�C�h�}k����Bļ+JLut��@i���%Lh���H��G�W+���<���Y���&"��A
�Ш��� ��0}k�;G=�/�}�j�t�%P�Ȟ*�a*#ԻA�C�%���;��.$��g�pg1d���Y�Q�MgWp>��J�VJ���c����+�[y!c0LO���2wd���JPGHf�v_�'���'�^�K��8N��-]���Uꞿ������9���W�gߛ�qt���k�� Ci��U�H���1��,��-$ƿ�`>�1/m���K�Z���>K�9f��6vE��m��\p�\ps�i���"��%&,���=����n���\�鈀Ȼy�xY��h��n��ʃ����XV*���G���v4�c� ��w�&�w���0�Y���B�=��0H�RC�
�ipR�AJ��t��Ω��_>�M��ר�	
��{<�=�6�>�z��6�f���\e�<����2��9���z�'ĉ���'
Q-��4a��kT���֓������*։�`�;���S�x�A�����Z(8����ݜhY��!ߨT�)��p��k�3 y:�u�'��E��WQ��ɥ�[��g/�!������.�����nQ��s�R�iX�'B�+��wj�n���܅n����%�ܞ`\'�'���wշ��8��<��`��y|0�8�'�����tUΌ�]�X6��,��2b��xq �:&�{��y3�9����=_~��U'`k)К�]�AM��q���E�ܫ�j��Жq7�S��y�C�]��tR�w���w�	��t;�a��w��L�mG����AC�0Ű~ˡg�-�(��h�b~T������}Q�~�LI�h�vI�g��J��&�4Nm�e~<]�N�
�	����� �N\]���?τ2��R�DsNTք�%�s�R�ï�Q��=Uu�oI ��^O��Q��Q�K6�^=�~ *��H�(�:BW��ufW1s� �ƾ������/�������\�e5���ji��薵fjs�P$:hD{M����넯��Ƿ�	�<�z-�V���0D��QͲno{�,�FA��-T����]���$Z��ʒ�5_)�4�.�t��M�$���?r<m}�� ��e���g��	��}� ���e�[[M(�Bȋ¿��k`�f�8���S'zə��*3�T�?����[戀����_d�n�f5�t��A¹2O�Fr�zھdr#Sa�%�/�c2�p�_���P�4pS򠀧Ϫ;�鸅:7��MZBg�`�/��+H���kI}�-#v���7�2���/��WG&�D��dp�,}�a���Is;�]�!��)�UFTt��V���^���
��oE'ɹ�G����1��*av��$.p�O糨"�aǦ�tt���eS������7��ŕ�~B��P������A��ok��,
�m���C�lR^�}	�o�.5'^��+�6mPAB�dG�x��k�/�h�5���i�#�-��M:�yB�}��� ��Ac��#�ΚЬ)�d��d��b��`G�v�� �<ly5î^���`
S�
��̉أ?_ ��{K��M�?�%�%��r��*XÄ
��R��k{n �n�v K�R4+ׯ�Yw>�}4�f�������61���5Jq���Γ�`6x�'
f�]���~������R��~Y;L�E��]��C)r�"���E���Yح����"�1�������*��T_f�)덐B����]YTӸј���m��$��qLq�m��	��窙xC��'Žf����XWH�s>�g�ikU�a���^�]��@ũ�&K���H-y�
�f���#�H�7�U���C	�ؽ��ض<���g>�%>l������Z�2�MsU�à�R���񮾍���=h�i�7�i�BS��RO�'����dvH\�S��I��W����c�Z�℥�c�n߫�=���3�0u��FI4��	c���:Ϟ`m<2�RHI�0,����8҂R�C����?iug�����)�/1���=.{��ߏ�E�6��-������ :`�b�o���5�5\5OmI��k�H�C��|��]��]�4_��H�3�,�"��*� /��k�0�Xǃ��I��^%��6�_R���{����Bz��/�=��
�(�8�Y
jG�Uv2@��	�EcqȌ(V��B�*s8��:������K�G���|%:K ,�$S9M�s��#�\� ���:�O��E��r���������4��ua�V�&�g�C��0����Ns��'gz&@�Ҫx#L?���1��~>f`B��6��ՕXÖm^���+!�\���7��s���R��IP������?��p�1*tK}uMYW��Zv��4��ldCU0c�۷�<,��d�,E���ՊB�Iʽ���␝�-����'��]�N��W�0�����
|�j��Ѧ'�;H��Ӡd�L���U�`�8;��8�ƿ8��p]	����a�MaC�Zڰtǉf��.]q����ɤ�U3z�v {�vه�(B��Ě�p@]����S��ؠ$�f�R����)Gh�����g���Z!Rw� 3�D��J#�zt>Ds��:*�G�>A�C[�/�a�����k���5Q Y�U�v�Z�?�oR����z�ɕ��툃��+������q3�St�#�)���:��שu���!���(W��m:Nh�PC(��rZ����g�~X�|c4N�B4㦕^,Τ!j�G>"5���b
a�nE�kM�������W�#�y}����C�1����[/$+}9:w���2D��`[�:���\��-�}!tSU|��q�Bo�痺x���w���W�$"J��%'��Sۊf��f�K}��|����\&��@���o��,��i�i������}�9���.��C�8��;�KQ��?"O�Бb����۽rFy�CF�FF^����8aL�90=��`Hi ��3A螷��l��E�])�7��d��9 ��P������?�|�o�_�c2�z1�6�l�*\��M'�|���t5�1���I{�9�9
�S'q�bZ5�$z��ٓ���t���r�O2,�)m�&��Ě���E���6`���[�߶x�.��k!DX�9S�?��y�E|gPg�-����0�$��Mŕ�={:S�i�g�Pn��tν&�{ٵוG0�)�z)�0�$�X����	a�c7(&ww�bu?̛5}CL/9w���O}�*R��Tܞٜ�L��ӧ7�E&j�t���$G���G0�������f�W"f�=Z�G"��{3�xO�-?.:i�.�~��m�ܥSM�>�g�\�'�ǕC�D��`Y�x}�=�'�.lN���<DƓ��·@~y�s+H~���Y9��g!^M�����8;��S�ز�!�����fx�l=��� �r�����I�1��mw������1��ۉk�F�q#��bo �ē�.�=��;�H�=RK�h^��|��6��(�d��)���3G����#q��������qF�������|xI\�uw��j�JV5:���8[��2���f�H��>�93Qo���@f~��U�C�h�*$�76�ڢP�O�h��|힚�,�H���g���%;#�![����f
�\k"�ӡ}�����A|��1�ays������x�׿��$��|�[)�g Oз��b��Lv��~�x�Cb3|-8��^wK-���"���*:��(����n v-t����'�x�Q�n?�O2[���Y��JB�:aH���3װ��&�;3c����Gq�&=�={َx�a\9zT�T����G��Y$�ӂ
�?�յ8��"�ӫ$�Z��o�Np/uXl��mc^���Ӻ�pS8�oe�Hxg�,b8) V`N�4]N��X&�	�FC�	�`C�f���!I��sP�u}�n��
�d>
�;(kI�"p���I]ج$�m���g!��R����6�n����i��+	�A��@6Ł�ygJɵ��<��;���� f�c�n�.xc�͖W��\��|h��P\��N����֌^X'Tq^�H3�&�X<D���f�o�3�؇��n39?J&�<LT��W�{��^{�q׼���-��3+2H�
�adtPe��>눱�Ѧ?���YK�L�5�4Xb4��K���s?V9G�����QJm��^_u�����z+�!g~I�[�}�/O�����x����|��&����ع�;�c�����`s�������׋�e��p�����{�ҝ�omu~kĄ�~_��-�߭�j �Aay}���e�n��	5я���.^U�xm@ױ�~MX��'��f�l�[�fZ��2�j?��Yt^�f|�K��^`oC�u�My��x3��=�!@*����֎+�t`�a`������OӔ8�k���,��`,�4s�Y����6�:��|j�i�i'���~���Y:9���g�*#�jS���b�/�LZ�q��j"uj�/�C�����8	����-`��B���r�="�	E���8�yQ��>��U��F�����Rή���a�{���'��#��,n�!�G�
��m1Z�x�*Ijw�f�K߭L&�Z��C]�e�#��='@�+\/t9,�:��oP�5AfE0���}�(`:|	³��I���w��?+_:�<`�J	�5v���B��~��I�$3�rV+��W�иzf�%�� `% �T�<k����*֏ޛ�K��,'��;�g8�>�3�T�仄^��Ԗ�������р�ǣ/w�����3����#��e��"�S	�v�)�����3���ڽ���;O�Y{t��4v�>����WĤ�\����Z�������:����{���y��rN��z�p�&�̀V2o��?����w���o7K����r�[��)�\~W���*�.�/q[��}`�=J8��y��ۈ�'�����zuYb��̶�_����S�mgs�{���G�S�y���q�,_c��xC�j�ˍt��<��x�C	�J��0�Ĝ���	���0?�ͽ3G�Л���� �pl����=�Q��6�	�������;h��Խ�:-^�/V������
\�$k`o�_�������ux������P;Q�d|{�$��� ?���L�lOBM)�EK�H�ψ�6%�?o�x��3�)pʥU���E��,�<.9.@�9\oU�=�i"u�/��$���v���|��~������cUv�:��}  ��+H&��hn,!4�8�ݶq=o�(��q[�z(Ӊ���(+-���1n
���й�<Fc��x.��T�����3i8E��%�������/��A0��؉��	���fp\�����0�ӝ�e2����s�ۓF�]��֒�?�I�j�/0�"��煥�j�X0m���w#�3�'x����=E㊻
i�fʴ���o����)�ʫ&��)��Vn`>�Q>`v`N1��+�0�fJ��5M�>�����:YP�|�"�@-�Dy��8%�0��sG?�9�T�/���`��:�T��l��&�:o��q8�����if�M�����A��7�u�07�e�'4���WF���vD����{Rh��Y{z�ڶ�(��7z]O��bwTΘZ����h����_���a��*8��A5¦����vV����_�K�%@��p�����u������}�����Y#�9=VvT?���OH)�2��H���G�� ����-�m�?�x�0��G���~�K�J�*�jۤ�8F��T��
T�/�n��U�����Z�/��ˮ��/beC��	ݏ���0�#h p\��K��8�!8��E1�XӰU��
����:V��@B��Q`%�wd��-���3J�w[S�Ƀ�gd��g�|�����J����<�N�y�����c����_�N�
Ȝܯ)G����i� ϰt�����巡aNmN�u�4O7Yd�n"��Ɇ���)Tƺ���bpf��	�rL�����$-��/�Dr�T���wR�%CK�>�,������,��͛���P,���//� ��1����*t�%Xɕ>"{]���KK�WҜg� ���!�.i0l��J���-��vГ��xU+�J�#)q�w?N������rk�gt�4n�����JBO���d�;g�)���m��
��(| �S�j_��h'n�{w��/Er��z^�&�)���[�n��$A�;�K
j��ᝳ�d���ȥ�2
��y�����E��PA�����R�㑮�c��e�r�DqF�q}�jK�����1�Q�4&��D�������og;�Nt/8���qR*+�ӿ�H�%ٸ�.�9K��<ǅ���O��T#�4�L4��K�B�iU���mt:Ϡ��_���9�y�z�quz�v���7P��_Dso�-����&j����p�h�r���:>�Plrc�/"����!�2�U�v]���fq(/`��u%��A�ܰ.įAc���B��j��_h��Y*�ߒ$�1(0MAO�7�u�� ��f���ç1�p��5��A�ڵ�u�٧�h׍�-��*J��A��O�x�&u�iC�n�T�I�qo�=�ʆ$.�#k�:�Vp�n�i��8=݅�� 2#�l'�+�8�m��y��Q@��˓��R�E�t`b����(�*�x������I	�Һ����Hc������̵M�ւ��}Dfp�e*�^���eG�>�n�_R����"EP�'��Z����0�n�Z�)��ů�D2����vDE>���4zY%�yQgl���a�G"���C�o"������DZ���&��%�94���^@���h�}	��P�I�
7`�n�
���RR�'ͫ`�Py�;��q/� ]-��?�K�Q����e2��{h6�A�'���lNz�*y�^���(������v55K1��/Θ	ES`D��̕�pQX�'o%/w}9���:i)�E+���?[v;L��!?�"~娗L�zL�D���B��g�8�r�lf�떡\�-��c� z�3��G����t~ �V�K�g������8W��Tw(�,����7�����K�h�����N�ٽ}7v��D�aϊ���P��v9���ᆽ�:"��7{Oy�8��pYNy�|Șrr�w�b �d^L<�P��߷��
���Q��]����Q�Yopx�h:y}�(	e�?����RmϷ����{"����J^��:�̬B��z�丙��jVT㖋�[�QI�t��`��{��dR׏�� ��Ћih��ť��u썯t;�[����-d��ۤ��C'1���<���'�����&H�uJb�N�0�J���ҨMӘJ��2�����_��p�Bn)k�;CuT�y���B��1;��p+d��2���yy�ȗQϛ���sL�-	!d�����Ti�����y�*r��/I���If=z��G�ZA����$ɭ���Ä}�	h�%(^�e�I�N�<vu%C��H%��tn��<J�e�Oє��X����uf"��W�ޅ�>�� >� X����lr	��mh��k���Z��@)pcŭ0������o\J�/�Ws��T	
: ��9φ��XCp�ʧ�m3u7{� q#���Hj���ؖc��_j�C��ÑY)�p8�����<# �x`4�-m�K� �b�Sc��H=��鱟V
����F���6�~E�4
�9{]�v��Ĵ�e�-H���e��'���r��)Қ��\4�/�Pٌ�K?P�t��[\kK4v�62DF�D#��aF�l]<7d׬���]��ݐ�$����޹4��$3�#RL��@n���]���8��uF��b~���K"�ʗ��g�;���bc�~{�)!����LDx"y�$����U.{K���L>YYC(�j&h��Afiu���),�ſ��7��Qޛ��-�D�Z��nfJ�״Hw=G��� ߇i���I�U����0G�)�;vZͫ���AB#�m�9W\I'�ڎ�}�+�+B�ia�WK �q=��ݤ��\�|��"����M��<�9�Tx�3��n]�_�����L���j �F��&��o7)���R2�$P[�7�N&n4H���$L�}\�������p�xp�
5��P]��r3љ�-�B��s�XH߼�$z�^�]�	D�6�I�ψ��.���j��0u��:z/���E,�ȉ���r?*��K�IN9�C�*�qK�s]_���8�>܆���I���<�a�֛
R߅�(�>����x�a��y8�k�
 ��L�U0ư d�����F�N{h�薂%�1o�҉ {�����*s#�{�OZp� � ��;���{Z"���l622$o� ��*?C��3� ��$�Z��[���F[LE�j��eo����)Ԧ��PV�0�\h>��1W�~�f �⢩.*'F)�{�1�d��y�dS7��ҕ���b�7�V7F�u�c�l%O)�����${�6�Ρ���&\���fݺ᧽'�f�ć趚�j�֣d���9T$��mj��WRh��6s�Ojq �3�5�Ø��@��rt��x�0�G%��3}Oqt0[�FQg �j�9���Ojا�6��Z�k�S�)A��9��KKX�ڝ�ۑ�>���e')�m	��w��l�4c-<�n0�ۛ�lG���F���yt �m{MbiUj�~�4Y�G��Q�}�2����{~
ט�/���� +7�Q��t��Tb��4�^�����)�
�*A��Ī��y�P4�fb*TTZ?��".W���I�['U�^<��%mW��ziX����/�"�M�a'n
���Q����3��ZǑ��Ac��Q�P�J_w��G����5+V=��
E�5�^����-��gQ$Gs.��#4Z�y�u6T!�'��aQwX�!G�w�=�6;��e��d�lfp�>���O�8�nd,.��J �0�|��H� �4CW�V=����_|ph�Ϙ����b'�Qzz�����U
��I���S[d�[j�d�O�ns
�v"xI?�8k����酃�"������^Y��-���Յ�E0�������+4C5�V���ő��M8*�쭼3o-���3�G�iʺ`�CZ8F<�?|rr>�i��/�B�@�� ;0n�a��Bh�*�&�o^4��86�":�^"�b�}C#�������{me�gh��F�lt�ޡ���a��1S�iD��a�q0��=壱6�['J[i��'�`$�k���s�혅�/��e�k�w�Y᫜\����HQ�@#��2�����s�C�t�l��G�t[
����~c�]L�$�ڇR��9�'�骜���7����,+:�ˊo�)aj�rgQ̷�����2xw���`Ԃ]�w�[���� ��p�xRXizE�?߲���iR��?;ƈ���dPZY�Z�����Ӻ@�_��g�3_��P��G?bYAԙ�E׾�|�2E.�?S�͌ଣ�����{����� [�9'1��w2 ����KT=�?��4y��|D,}w���`��������Di�MĀ
�8�D�=��]A���6^&��7��v�� gKg%z��p���¾y�� c��o���t�tW7�$�ٍw�]�h����q�6@�5�j\��@���-�xH 
�0/�W~�J���Iȣ���n%т�@d�
�(�i+2�"���М{��C� )I
��b����<����>B0�^-��x�,V����ůh�9��)� K�.�MXr��vʮ��V�[�[��Vs2WUt�~;�k��H�t��s;��Du����� C�z�&[;N��EA�gaR9�������U&�����hz�`�i��tV=��8	uN$L��r�!����`�u��F�+�I�
��`�Z+)	�s��;�&�[��������:�/5�[<�缦�"��Z�A��^�|�O3V�	�%����`[gۨڮ���4�����P�t�E�������K�ߪ
�'���V�"�RY���&����ËF���J���[p]�oPa{ ����]f8z���<��&t�{�%g&X���@��m==7i�6j0����h	�����U� LI	��A�)���M3�[I�*����� �{��j<t�?�~�.4� �)����\�f�$U(��y����!�I�ߧ�Qd=���߹�ڋ�Z�4E� �]6�~׷��3�V���͘yMY'�;I�w��kl��K��ζ��������>Ɛ�\ܳ>W!'N���,��&�ϸ�yG�9U�� t��Y���F�>¾#^vb���j��l
�I9<�Ƹ��l>@ ܫ<i�_ph+����
!�S}�%�r�_�[��1�z'z�.�.�Jc!ރ���/r�I0�����x�6�� �r�&>�_G[�

�re�;}���P:�Es�W��'G�m�\tA?�S�H��)��`d�� � e����B��ȜVو�G���fR�kt�/?7��
SEi�η�R�Н8��BmƮ��)�jd�w�[l*��cjߕ�:yc1���7��%1f.���rf#�FGg�ƪ��JY���r���'��&y;�W��[1S�MB�����/�ʅy��@3�����V�I��g�!�Y��TD�������lUbɟ$�I�î����3@���9��p���SvK�}���>�O��
Z�4!��C�ԉ����^�t"\)?�ܼTa�t*i���*$攆K����4, T�� ��t8��A��H�Z)����:�2v�?�\(w�K���[����V�#(�*��?�n�Z%�I�����uT�U*���P gs��n����K�ܚ|`��=Ք'�'NF�nyE)�$ ���z��{�{t.���C��-�n5?��4�s��ydoO��8O��=r�.����L!���P���y�o��^M̦kl5[
/�D��'�:�j{(Ԃ���*=C��ɯ���h#_Q�C�T�����>������B�nGp�>P��c�0�+�Б�S����� m�6�p�����AR�����Y��Ŭ���$�+�C��w��j�S��#�~���sE � �	 �n�Zj��E'o��=kp�u"}��(����Z]�#����S�I5����e�Z�:ƣ
ο����|�L��u#�Hz-S�b�C����B-'C�*Q�h[����l���{����h��*��H����� +��N��X>�2TM�?! C���|/.]*fboPZ˲U3�� �����U.zq;g
�(�ߛ���~�W°���4���l$�ɜ���ޏ�����e�L��5Wv68�'��W�f�(�پY�}{o�83OjQ긕��ú�1
���o7?y#����*�>�9�*������}p�K�^P�t� �e�N�Z�گݴ	*��/5U����~[cם͍�c9�ӳl�Eu?I�Ά�&����q��}QY�(8��'���u�qH���P|� To�3ՀIU*���f�SJ���y�����WE����t����C��èt�<ǎt�xk��D|5�um:i�5�-��٥�	Y�㌜y�d��M��;uH��!�&����{��y���5�]Ř���3)���9�#ާ�<����{��-�A�oE�	�ց2&�� ׃4 ^�2j/�?q��*((�gE��_���R��60��Z�|���l~�v���!`Va�w��Q�v$�>�O��;�8��\کvu�UKA�i��;��O �9��o���ne����ϝ�ⷔ	�k��l< ���>Y>��q�Cp�u���!�#�.)��u{�*�H��-:>�����E.���n���֛�^͒�tB��]�>������`gC�9�@mͭw�⏣���*��
ψ�TA�g��TMT�-��}�T��������9���Nu��p,��0Fuz�:���kv���t�R�Lu7mj/�.�"�G��֑��x���um�CI��fg��;6�57�[��X�07NI�������M�����7�HV��cnB\���V�t0:eFn��%o ��FJ_�^
Vp5��ht.�*�R�_>S��\g@;�zr{�b=���>t����g@�r[���d	t�)��*�>7C��֊q�+t���:f�g������$�0��}�@	�����rc±cc�L�vSD��*�	�����'�)�Q�y��9y!G�4ho*8YV��\^~eN���QҒ�/�k'�t>��E7�=R`�:4~�b�<s�^?N���Λ��t�j�c��|� �.b-�<�yi���^ʞ�I�����/���WK7��C7���#�P�H�)��PT��(�pRW��c���O�D�]�CGǫ����W�[$5��+c
i�)H��	ꭜ,��&�W>�gb�A�Bh
Ԭ�3L?af/������dJ��d���H�lu��ݏ��h.M�ES�&��%4
g];�7L�^O�N�a����Xw��Q�У���V���,��������$w��q2̸�[_��r�g-���FEK��mW��
��h\9�<������Α3�Ri�9�<�OA�+�f��L3�-?g�Ec����l����P����lX�c�F�4\���׺�V��V�u����=q�h"	���0/�FQĠ�|����9�໗�i6��F.���GarmpE�Ni��k� �[�;����涀��0WKn�H�������f_RY��cP�6�Ɋ����
���1zO����j�d�� �>y�
ڷxU����OP0Q��������Nw��Ns_��H��D�ZnA��ٶ�U8�?�;|t30�:�샲_��G=C���a�ˉ� ��y��&0���V}��l��um?R\3��sco7�ds-��r�# _6
�W�\"�Zo���5�ȁ&���xe��
��=�;�Iv��\� ��3�����CPS*�GpY�����m�Y|A�ݬLoB"y:[<��6�g���ڷ�% V��k��R/�2y�&I���W ,,�e~	�ʪ�Be��Bd��z`���\�4�Z�f#Gؒ�#�Y�s�GN E�J6�D�i}�7)أs��B*`$�aν���&7['��Kz["[�H5 W�϶u���:�V��|�P��y���,lՍ�/l��\%�C�|:����,�\��� F2��.=��=��r����Ȕv7g&5d��'M��$n�\^|4{�z��f��g������xdwB"��g�����+��e@��օ�g����%ZS��}b�/��
3xc��������Y����usH]�PN���H0x���[�]�d\�n0>��ÜDqg0 $ �-�_G�h�CA��RsL_���9��(�85�
��D�t��	S���N�ɓ��Z��5Z���>Ѥ��&�zFK��_��WM���ZLt�.��O���vb��	=�7���P��q�b�HǙ�R\��h���!�0(��A�D��I]*m�3fT4�m��C(?��U���9��vhv�,Z�d$��Bs�*���v�N�N��X[.B��(�K#j�	�k�ӵf1�ĐH��M3�ҍ����sb�a��5j�-)\�3��R�*�5�#�"�Ы,���^J�W�hmTė����5�,8��"�=�]���W3�%���UƔR�����#�m;S���$=��q���3��v�.O�8v���4����Ȭ#��L��v��W�kb��8 �������2�D�]�E�(�s^ZTK�v���J�*yϽ��$�	��j�"�UZ0ʳX7�����0���ƞ��xX�kͳ����J��獜1�A�V�y��� ����@MK�CH('���$�
��F)~��o���2��Ω�٬1#���y��EO���A�p@^_q	�ի���[�BLX!&�V�����e���-*���ɴ�Z��ʳ�أ`̿���~�� u��
�j��`�����/A�=����I��(�c ��_ �ޘHʾ�? ��e��'��=p� H��Ob���
�`��x�?� g���Q��fi�|��Ʈ��OlbAQ���sI��F)-��e���q��o1�F5�92\��ߪ�ņ���Z>@����q�;<Ĺ`�M/H�L���01$�JpkF�Fa����j4�J��N�kf���O&ۃ��tkP��P��c�=��}�T�(7&�Y[�[��54���!IE��;��&^���Gv�	��Uk�N� v�DܼzVJ��ܾՈ�I� "ە*}�������ӹ\�9Heճ6�_E�&��3�E{��G�P�TÝvt� ���7�8��i�=�M�����8	H�	R�s:���B�\)��Mn7>��yx��_��tl�^��"۔�uɎ�*�F)�dgm�#i,`��
4�
�E��GV���%	>��&�����c�_=�:�`&@%],ZyT�Y�c�5���ژ)�O���ր=��d�FS��f��W/7���3���?���ϻK!itUp�����3GBܺ��$>LHHmf�Z?�cr�Zk�����JU]�/�'��P���͆t1'��nc�rY[��I>}�*�F�#���PZ���+���qGЕf%	��{6��o|�JXȐk�pϻ���Q�1v����x ��V�
��hb-��W���+ ��x�
ј�f2��R� [��q�}��a�(K���H35�}���?v@Zt>B�L�7Q�]�H������h;6 W��=�&��|~=g�zn��������ۏ��8Lp���o´3��J�2�]ǜ�I��b�3���b�t3�8NtL#
�U���"��F]���w�m�7�@���j}��
&f�iA��4j 	'�%$�j,��CR��fQ����F<����O��Prɧ��(̡֩��F�F��(	:�WC7��j�+�N/On�u�z���*=A�\���Z�H�n*��F���N;|�/BzXI�3p��n���ܠ�\G��[�t�|�����%l�ة@F�;v�k�L(I�B��=ݷ��V6:�ẏ��ޞQG�+�p4Ʀ)�a��$�`����VAC��V+�����fQ�2�A���
���h�}w?M7��ͤY�7V�YڻJ5Z��?t�G�L�ϫ �h�uXQ���8Er�����d$�dډ�%w ���%���;����i�@�D��c�-������^]=��O��(�&k�{�����Y�D�!ڝZ��P�ʯk�6��'o����F�S��s{��]���gĵGڄO��o�oN&�!~�<_h |~��f���Mʉ��6��.�M5e,lL�^d�0��Eؐ��4۸�1;< ���j��g�C��ং�eVD�Iz���[':� 	'�]}�x��}��T�Fq�Z��ݷ��ǀ��5�w9����^���s���7����:#Bw��6`�2���qf��_�����!�p�RF�Ǹo�ʼ�=t��!M�#�ũ�9�%n�r���T��P��A���uY;9�7Я�!�d�����BT냵�rJ`���n�\-k^�����r |N���[��]������up��(��㞡�xE�x���~g�NU񟑇��"�#�)��<'4�~��Amx��:�}�_�9!�\���	�$��-		e�E�B"����^n �x1����8z��� }ΑЬtyf�ҫ�4�O;-'~<�!�PERj�8�ē�S�=��	��@E�tR�H�on�js�g�Ë�-�����X�#<�Y��9J+V:rp/L�'#����v�<���	T*骽���WM����Cݵ�������9��C�A�pik���#������}Xo�Ӎ���=ƺ���u,�_�qU�Y���[��6[�����W�܉� p��1["�|��X��>��$���fS�5���Z�p������~�������t.
�j�|���$�f��v-�x�E� sX����G�P|��X��߹�?*nV�{�c�0���W�L���d���c�z�<bm��� �uG��_!r-����(�}�pH��*N;���g���~g/��Y��*�瑞�)�hi.�؏�XJoө���#ո xga!�����=���I�#Zxp��ȼ]������h�|n��������z��p�wA����6g/W���W�oc��T��jN@�9\F���&6����Tߌ\��Dn�;����V+��77�P�se:�Ltd��?�b:�ʲ�JVlG�L�A>:����3�����Yi/�@���Ů$hY�$���r��V.��xEu�D(�?h�C&���f�l>ǑN�ێ�`+�h4A�=vo�;)j�W�Fm�Y|�H3�L�E|�('b�Ww��`0�Y[/�4��
:�r� ATx���Dc�vn�V����L$��)~��.:��������
�����m�����ҀKh�p(��8�ߞ��3�J�D��
ֹ%k��X2;|)ӻ�Fz��C�7�r�@���@PTm��{��X7
hX�ml@A���� ��)��}���BD�L6�18�4�dkS,da�����:����B������t�A�,�4�f���������;�cm�3�pc9�'���u�: �BpR|7�W���;�����Ź-��|���2\p��{;���K�oQ7`�P���!�j�V �*�rA�+����;��ZwY��ϰ�p�3Η���_ ݗ�\���V�V��������f�xT�.�^�p\}[��u}�wr�/	�r�[��"W)�Z����.��bC��{�	��v2�C���ٮ	�p�<8SP�&�f�g��L;�Qo��Z�	���&��LW�����+/�Fl�g���/���Q�V�x�eSQӗw]��g��@O~x����V�҈����_���j�(���{���irK=��Tq$l��&�n���9jf���bk��\�l2Fng;��F�*Mn�{ɶ�ҽgϕL�t�K��ݖ�U�:��PWkT��$x�=v��u�$�0��0DL2&% H��uV�%���k1�a�
�Q� g�x�'�}I��+�bw�f�rAR*qV&�=ˊ��x�X2�C$�e]o�a�h	1lfػB Z�fGT��I�L��d��N����1��h!+���Q�*���dA�?�m�[�n�hFϢ��(�c`�������6���X�Ŏ��=�89�i9��q��#��L`�Z^�/M$H��T�_J�0��'�Xv6��2��e�4ؾ
@��^C�4���D��`�
� �OK8��(�W��}�#F��M�	8eEȝ�ĥjx�n�j�P�����YY��o�����@�4鹏�Ӷ��s��`j=�V5Q_�e�.�l��=6	�{��Ք��Oc���'P��?I�(�e/�E�Iw�����i�2ǡ��w�cN�d"d��nt��i8��=�N)} �*���`JJg���fC&�'T�!�M`���JA�*�ϰ-������	��Gci{�9q���d���<y�Ls�(�<����v8�3�͓0ִ�-_vw	NQ3�AŰ�ZF����;�v��	�N���II^q��Y�����d�����ڛ�i+vK+OSJ�d׿g-S�\��k��~i�{tW,���s��#Z�U|����4̨K���^�L������P�(���zn�ݦ������:�]m ¹�ϕY[>����>,�g�2��O�\H2��S�Y�A��&2��%׃DQ����+�o�̜eJp?�ꢤxٽ
�w~����A>��Hl�����:�j�3�B�i��7-dn.}vV�Q�k����x�؏g'������x��A�!��hb��^��*�暾H�L5�&r^,'��`�gr�k�����>��p����J�T_���3��f��Q6����9�A���n�3~HE����l��#�G.�=��$����"�P���˲��h�i���tf6:��JDoW�3�j��K�X���r�WD0#~ݬ@����Xt���[=,%�lLQ��]xe-���tɩ���K���g7)$��++ʳ��7�g��m�Z�("��z�;��6�R �&�p*��~O��` �Ff��F;Qs���}�q�8��LFIo\2�� 
���Ly�e�ݐ���@�w^I�9��.���vx���M�
�B�E˸��!f.g ���=��&-�������=;6]
��1�n0m�١
8�����p��,��v�L��עo�J�n�*L�{��Cbܚ�VYI�a��Hk"�#,'E�;���"H�]�(\�8\JA���q����ک'��TX�<���ZO�c6����NXI9Z��"��NL�~Y�[/�}���7��u�yK�  5�a�.�����.t]�q�utʶ=�P���VR�s{��3��e&vk!Dk5�d�J�'�[�����C=�1m�.���W��p�s�\L��0�	~/	�e��0Պ;�T�2A�?Oڍ�WKT�N�7{ �$��=���%��rw�3���q��C�bY0I�:�HH��]���z�yy���%F�{��A�_�(X?%��ؠ�+�q�Sw"�*��C<��=�|�*Q�L��ܤ7!`8�@c�h)��P���K�!_���|X�ҕt�qw"M���e9���X�e����4Ϟ�\j� �5�)�'�2&�G�A}ו8WH�R)j%��p^t��$g_z�w���� z�pW�o�
�mt �a���2�}��(�W�2Ԓ(�\wx��z�a����x ��D�jAy)(򺱊�H _4F(P=���3.D���m��:J��Hk�� kE��Yu�O\3��4>�26�����5g�g		M���3(j��4ś��Th�"z���nd.x�!m#�5P�#^(�DvO��s_ebD��0���!k˿&K;$ ��3u�V2/�\r六�5ԇV3�۰�����t���T�����/&�Q(F"�X���#���{���Ú�0�#KU�������\�M���\4T��%-��r&�h�U	�!��x_�:Qr��߬���,��b2,�|+�P�p�	$�?���D`�Xޗ����\�'��9@/U,�-��U����$����W�b-�͟�������a�ƍ�kuN�F����A�0P|����_�'�G-��z+Fa�A���)C��m�:�-~�;@��D�}�!
H�3�M�d�E�ހ%#����~T^7A�� �vƖ�`�X�PChY#�w�_�#U��d�It>��Њ�K3��\Q��M�O�z���X��BX�>���������M���X���
lԎ�� ��t�%�\P��w�PG��W���MtFj�ćO�|�ϨN��ـ���B$�_@������c����x?P���8	>7nȴ�(��?]��� ��Ϊ���P0�O�9~䦙,��gS��^4#����O	�W*��A���~q~�g��[��`�����ȑ�H"��Ա	���f+T�d;��v�ԢT$�l��M%��`���~��r���4����i{٨�/�G�[���h�7@�&i~'�	�*����i����!����� �,a�"�zW�^z!�J,��U��8�	�p֊_E1���&�B�ȝ1��*78���X�xu��6��B��Q=�}���Lí9����P�
B���m�	3mq��m�kl���:��*��ԗ�C�\����(�
W�ZZ�����B9F��Yc���6����8�Pt0	���	v+�7�G�(�Ź��2���M������c��m�t��g�Z�(�C�6��q�?Oa�i�+����"��z���`"A!��|���+�=���+����j��V��#6��'G16�Ѡ)H��vr�]���mm�jm͛�:E�b����CL�셹��e90U>@x&�/L�n]�I)Y+�C�:W!��k R��B0F�@�w�oE�:��ˇ�w�z��ԝ"axm�� 'ںwK��zsќ�%���{���!���Ny�4,u����' ������Ԛ�]a� �l�Q�Yq�t�$HB����i.9����m4�>}�}~yټ�4�O?����S�KQ��w��U^0_�b���k�Q9Aǌ�@��s=�~��qb�z���>�Q��_ڋ��;X굘�$;[�R`6w�EZJ�9����]{��MAQ�����{)�D�~�@�_!���U+�ޗ~u��ԥ�V�*>~"6x��\�y��sq$#f���f��>�JS��g,b��a
Rt2bɇ"�f���!H�/9��\�qɡ"���2  X�ؤ�XF]}*둦<bƦ�tP���H]BC����%�%'J��}�P�P�2��6�ѻZ��Z%�LQə^��Þ�߄�9H��#�OJO]�h����q����� @�<Y^AXm�Z��eX���	�g�d\������j�%����瘪�#xf���AW�'v�	T�_!�%��YD���Q(�&@��v��˥�-�qy��[�ٞ�����N-��ܶ�$�1�q6��!U*�n�0�PD@���S3�nK�j��*�c{�+�;�e��P���e'&���b�/��<i���U{����R	������'�_�c�g�gF�|��5��YCkN�^��n��3��~m�?�n��YH���O`h>+�d7�-P2=
�?߯�r<��6jWS�"��E�* �`;xA�cb �`��*�~4����f- �����ҕS��ƣ��	�OԻ�ٮXWw�%�)��O =��gxv�c��qא�w�x���
o�7$��Ȣ�p	Nȁ��ë�'���`�(�a�<˨N�tt�6����J�x�K>��GA0�py���v5��Q�A��W�'�J:�3po,P	kn��E֑3�x�j*��(9���	ൌ,m~�s��5{�:��B�*�K״1�H ��8�1��!��Ug�MgS]e�U�-i�k-P�EDX�<-�{��xVY����ĩ9�ixm�#5[�[r�ԜT[=�c��|=�ئ?|#��,��������TUT�{ B5[�.zKM�����k�=��ʙCXw��v�C	���5��N�i	b]��3@�Kѷ��щ0���B�P���P����?��{
�?�ͦ����6s�M����䬩��nZ�"	����H�P�8�GC���g1y����ܚ�96آI��o;��[�4�2.y �tĽ�r"��6�,kuV�Vڡo<�$\�ݏ���#Ր���BUMC��訠2�����*v�
,|�L��y�}��8����gy�?o��O�r�H�ֺ{T8$��G��QlC���~E=���?ᱍ�v �-��o0��뚛�OI�Q@�m鲏���[i9� ��U9l����b�4�%��݌Z�b�[�<���{r��;�����8F:���Xy[��l��gg;tY���0��,�=�:r����p�֠���}��:kGҦ6S���1��>���?J�<�@t5�����0jl����j�r��]�MF�����Ɍ`0�����y	�Q�^�r�u.%���ωmgC�N5�����=.Jf��Mnep �F��E�i{E��HJ+��X�7:���W�pp{/ ��*��kl�YIgjk��s��������+`'kY�ID�(�Ri��0�+��:�&5�Zb���1���_fj�� {�����Œ��z�������*�Y�7�L-|�QP�L�ޓk]⇀�/[c"�wV0k���E�e�bޯ���E6̶m������!7��)�zg*T&���]���ީ��"x�FI�z�22���X>����띣��Ժ)&��R�;�D�xP�ͫ�N�u����Z�Ĳ��\B{��g~%�4�{��=���q��mcr�",]�{��؇�b������~�E�v�W���kijkw��r(v��V8����v�~��F����[��fMw�E1��G/V*]X;4bicN/y˴vOsrT�iȓ�����7���,#�S��C�����$����ר�Iue��r'�VUoXќ�'0eb�$��!YT����]wz*@�⏁��g��Y_d0)��T���#��Z�\T��9�"O� =�1�+�@��D�%��Փ�%�� �&5:p@��E@����階���ޛ�U7�j�S�8t,�T�D%�PR�~��ƕ�@~�%a.bؙ5�]�	��蛼�z
���~��!҉�5h�׋Rz���?e�c^��P�5]��U*��o$�/V��q����u��>m~��U�]�i��Ӭ+����H
�%�,v�����zF�1�}{n�-����:��N)x��t��+�4H�nL�=��m�y�a�D�� �9������;ҭ�4聬y*�J@"��=�R3�]�ؼ��b�}\����+��g��sN^�rr�i�X}�߱�7)¡EG�F���p�s��M�_?�rt�<s \�yMةg�>�PLU(F
�1��S���.I���_W��̧*d�N9Y�^�;6��L�<v�%]*��E+JO��D;�N���	��� ��cS�_����Eo������y��w�����!z�"X�'�G���S�� =r�Q�����th2sI�o �V#�T�t��!LO9���è��	���]G���q�֔�S��V&C�v�b��P�.|R��mj�h��Ƣ�a����1Mhf4�3P��4�z?������,���!Ǐ�L�+��q�W>kg���������l�8� ������-�U/�xr��E�?�ij���u����G�,MF�l�x� &��V%n�xN�r2��/�΢:��x�R���_�;y�}��]��=�J{�ف~ܟh3z���ew	��|G?��S���,P��"���'0)y�#z�8p�1�nI�O�<飮S�H3�₻�J;�����Vje#5����ˌ�B��m���ֆ�
��S ��]y	&b��-�F�X~��(�u(�j�����m_�"�H5Z��k�9+{K�����A?�ڈY}�x�/l�w|�xJl�%��Y�W/3�W�8pĪ`���DN51�w]7C莳�e�J iq�L� �˕`i���>���Dv���hD�!ZPeU\�S��؊dU�:GGp�hr���P�Mh�YC �b���X섚d=fn9�])R��gs��Sw��\LpJʔ�T�󎠛��m[I-#����^��c�h^vy�R�j��V,G���P�����y�%��tp{��
Y��[4�		�N?�ޤu�N�/m�6pE iE�(���T5���J��v�8�f�|��Fs�ag|�N�d��ii:)d�fc���<X7�nu3K�CnE?Сy
%`�;6��ս���R�ί�Er���<�L���-��׳�R��L�ʋ���g���q�����D	��9��D��?�V�D-�U�^pO'd�K�5���ݎ+v�m+�~R��-� �1�ͯ�=�i�8��9�.�ar{0��H�~q�U�X�cfGa=$�vQ�.�1��>��x��M���L�?��Vl���&�4�*.�-L;�������U��x��P�KO?0��,��&��\Q��߻��D1�r�y������Z�^���G$@��,��[6�$9�a�?5b:%XQ�;RX*4O7�2�m��K���Y��A�c���dS��^Hnȭo`�et�T�9�:ޑ���N�����X,�%	ڞ��b���������)S��r] џT#�4��
\l��!�������/a�FLn3j���y�D�١ĸ$;�4Z0�@=ć�b�"_x=gD^��KNd�>n���G3s.��<���U������,�1m�����|,FY��Y��f�"�&��9Q�¡K�����dB�E��E&�	���W����Zc�I7�Kn���ofU���u%�9v5r��X��gg	GjT+jHK�sKܶ�v�^���&xW����3���8��D����	��Q�d�^�߂�
���~��ȋ͏���!@T����f8Q�wXN���� �Bv��s�y���htf�v[�lO����ϒ����S����`�鸡��0�>[�!^����go�&rZ�ɴ(E,:Qɟ5�����M&!;����e��c%G?R�ۘpY/�A��v�ü XlO��6:𽽟[���R�imDN�r�J.e0�,v�F׊1-y���0��ooZLeő���_��b����Ee��#�l�F�4���<D���y�6����4)�#��
7�>�o �H��Y�CuR��c����jZZ\����E"�b�6o����ְ>2��!Ǣ����PZ-A��C��՝C'�7��Xp�����x��b��ي�FEI��GP�/���#�U�3߁�_}gPh�H�m�U�{��j���N@�hRP���^gQI_����`��Q�p�]�&ph��x����S1��̗���wW���7k��t�*�,�ı]���A!k������+�|8Є�E>_����W���;����v��8��v7��.��T��&]����9X��ѵ	�=|�Q��!���ܛK���[�rtŽu2w�kj�kn�Ҿ��֞ZDG�si��G�́�
%�tY�'6��x�y���v��������ꏭ�7Hr�4��yԼ/�X$��?1#}� ���P9&W�⏏���_1y��������7֕=��V�o�\�������/)A�e�W��� 
�&!�̒�q��T:�<����	W$��o�� ?������������a�*n�r(�9dj�3�~����f�Z�q���_F�GǾ	���0r,WE��?؊c���l�3#�
��}�p\���tg/O�y��O�}Ü��i��'L��g:(��k�&�A�Rܳ/m�%}us��Ғ8~�]�?��nɦ�4�7�si���ױv�IX����M�H�S.���&%gb)AM�K����Ld�Wo�Q�|���3H\���u6?:/a���kaG���`X��ƞpQ�����@�eP�Sb٭�+���^��xcϫ���r>7x�	O�JH'R@��t:z�����0G�Vl+�T�W�o"��C�0J3T=�#4������4�+{PI��Ң��9Z�x�(wT������o[k�mE����"�]�L;J�F��c���M:c�v��J��'���}�W,@�,�9�$�*6�Q�&�$�f�Y�Ş���}Q�쨸��co�o���`X���$�#3�����>.B8$Ƨ2�`�J����P�U��yxޣ�W��C���&׬y��cK2�L�p�/d�-~ {��ы�����OH��o�DV/��3��ݴ=��FI��x]�<<���$W����1���D�_�o�R?�����_[4}G�0|���c+���i������ϟqwWr~F�ڢ�ޝ�������3�0�V���s���Γ,�p� *��N�@t���K��(r�@v-���6B���Ey.�g��|�7"%Z?���%��Cf?ɜ�1���[��nh�VK�@�� tkjOy|��������Z*���
�|փ�l��>�m���]���a�-�=�
UNY��G��,�/���(�4�Mǉ����ZP�0]�1=�cA-���Y2�B��A.�МB2��c���~+"������|Y[?.�})[�#��@3�E���Ɗ�G���`� �.ME��=]�J���6�XVi!�[�d\$*<�����e����3,`�ֳ����� ��./���ʖ�f�/7�"l�(�]D>?S���?�c��t�	�i
~-nÖ�Re�xj��q���D�GmD6�%�c0��vf�-f������B,�>�)�keE� �Ј�$ڀ�3ntѬ��d�����vS��l�h'��B]k�R���R�Þۨ�,�2����XS>%�}�3�q�Bfh��'��|��j���:!�XB�� �T��(EӶ�o*���#�)�bi�3�?oL���_�S�",Tq漼���awU\�.��E/�������K��pʬ��1�Rh1&�e��s���.J���ԯg�M�W�zKׇ|�}F�n��)WO"�7dsu�����\Z�.[.�ɴf�xӲUo4}��Pă��s�ϒ��h�tQԌ���$e�g�e[Ah�F6�ުXMi��s��#@��4'_��Jx/`:�(oz�J�:	k+f���Ř$���U�*z��ƌep�a~�~.�#!�_���U!��^�=���Fsr=�eX.�83W[�$HDs�ը��$���?'��_���ݏʽXԏ���ŧ,���jB�2�p?A�ӥ�B��SP��^u��J/��4�pI�E��_7�%��=�������}lf\���@�e��`�}{҅������@�1��c@���q�=�U�D��e����JӠ�w�E1v�E�(��l�0�V:���1�>f8LA����m��iLP��ʓ !m��ї��V�5$m�b�z-˞�h�����8r�l�����
�i���B� ����G۶��R�4LWYn6�lB�v`6���c�R|Y�����B¬`n��(����V-zށ}Q  f�����r�K=![�NoM�S۠��*�X굂��f���<�D�6��zt�=F�և��D��?
��yv�!,"��d��QB��2�V�(&C�X�N�)r�^v$�y�}&��+��<<�9D�~Vsk�,�R�#��0&�w#gV�00;�A���B:�[ܙ!�ƪ���k�J�E���.���z]+D�48i��h#����9���ES-�U�wB��%<Z˒q�Z�d��@��%UV�iNA�������Y.h��J��1�o <Dʈ�uz/�CX%����(n��z��ķ{VsK����h�8F���Z�ژ�F7��������Y6�^�r1��TY. t��e*YL��+Mi�VC�H�EÓL����f����P�Z|e�U���ožiB�����9��#��*�+P��=�mt7%]����Q8����C�����ƑƔ��k ����L��f����8_������ŪO�l"+j�H��]�fu�̕�s���Z�6�;��m��C�PeU3�eb�D-�HcFz*�/.�Kv�U�s��I	�5�s4��k�h�%),����ظ���xڎS�g�X��������q]k�l��� ��t�9JY�o|����h��)3I����x�c�-�W9*�t��!KLF���ם�x�{b�l����.<(m�WI ����>=���v��,S,�̳�!My�~�����UE����Kή��������j�b"�k�B�Q_#MM�ZÞ�=�Ⱦpc��p!2Eڈ�{�<ވ�lzXF��ډ�\	��9|�vqə8�]g� ���;\�F"��|�!�/=�����=�B�e��M9�q��U�{W,�+$�n�6v� �@�B��O���/9$���cQ����ߕ��J��Җ�]�����P��e�5*�㒡�4�N]�4�p,�����p	%�^�+�����	Czhn_�W���Ӧ�P�+\o(X�w�B��x)����=Ĭ��<2/#�ƫi�"�*�]P�P/"����ʐSB懊O�1�v�V(�V���P�M01�})�ҚPm>`�pA\+L���ϲwB�~6$�LG��x7=6�&�M&�FH$<!���c6}4o>��#�
����\m�"!��,�4�������r��2U�vp-LI�'�P9�(��D?�%�8H�o{af�.̊���?e��r� B�q��w؀e:0��;x�o�����=�X͠�� H�Cw�S�dx���FG��6��5{�ӄ�?�! F�F�"�[���*rǖ�\��� ��>ѾǊ7�ߒj��]�:�2�H���Po��S+~C�+�^�?�K�2�'�]��A)#��cL�i&��ǵaeVE��ڬw��;!��y��Y��fpV�ǜ�}]=s0 ?�� )�4إ�C"8�e!옫�K��2K�dݸ.���s;�|�<K�|'̱�[�
�5d��q�P�Y�^F�j���E^�[���CduO8fc;�%�� ǉ�:�q�l�9�l��E���+f�=�"D�q�Xر�o������U�!15#�%n����Taj�a9�6�e���(p�3͘��Q\�۩A��,�6�g~d����T�\ �e�V����%y�u�PzbȲ�!ذ氮o�0I"&��7ћ)��"�A#`�����RF�G�DαG鑒aw��/�q�:��PQk}T*��a��RYɄng!�T�);���uК�z��;t�(|�rи���jٚ�����W�.��gL�H���83m�����Φ�_ ]���b�m���nX��D=�˖�lTm�D}nwQ���b�?^�CG3��&�Ի��h�G�2*�`m�3������R�7����a�9܅"�g����g�I��#\V��H��z������I��$�sC�y��y���fbwK�gu)����Y��d��n�4geX����g��롉ѧ�����E�ǉ���쀏YFp �U4^�+�$��>`�ZW� �_ƫlD���۔�I�*y3R����'>'+6#T����Uݕ�����2�r�F%���傥���Ώ���Ѷcf�|�ɳ��,Oja�V�AlQ�0/
���S�k�J�9/��X���ͼ��?ךZ�r7ݮݔ1���K�EWOՊ����yz4�n�T� ��c��oSF�w6U�H ݪd_K|�Âc���5��RCe��������O3�£��K%��SU~}#mim�����ե�ڂ�7:T1\5]�ȥ |�m�w>�$D�&S�']��0t�l-S�l7�l3C��Rމ(ږ�F����0�~ݸf?n���.zx�~�ý�ku����-+A�,�^�㚧�!6�m]ZZ���G�SoV�Ir�%�f�+��h����*z0�x��Ih�Д�,O�8�ʹq\s#Ia��a�|Ѩ�ݰf�X3�&�:�+8N�[i?�u�n][�����F�l/�'I_�KĽ]O�P��,c����9=R��Wݘ��f�,/ʣ�K��RH���O�%�����vM}���Ŭ*�]�ܖ��Q�r� ���/���.�D�\�I�QE���\u�a�{9YP"o�C���$�GSEdB!0"�N�T'��m9c��]R���xۢ��u�w�R��۬ɒ~񰹴����\�vdD�׷���O��t ����n�;}����D_a|X�1N��Ŋ�a ��,�[���vU�r9���"�U�g�V]��O�
�zL�9�uǔ�0�=	��m��I�Wm����D`eK���> ���l?��+oC[&��/	R51g�HR�����O�Kl��c2��-m��#��"ˁC�����:��j\'�P J��LX�̨,2(��+)_�=���a��,�����/;��`X]R�O7��R�g�m/ ��yt��)�i�ϾoZ�1$�LfNF8(����x��	�����.������7@u��,<Ѥ��3��5hbBP1N�0-u�FpZ:"Έ�v����)��b��>�Ԫ��	��TK0qhPܑέs��7�Ζ��$ �x���3��H(���N���>($�R��4
7�?�q��I)�y`Ȍ<��!Ȉ��Uur Θ�Z��
��jנTڼ�T(r��	[�/�p}�7�1�	Fgq4��N�]!O�颱��kT������@4S�m�8�e�e��B"����X($O�F$^"����f�g�P��7��:Xg�~�==Φ|&!�cQ8�je"���-@��ğBGd�'�\@S�L��܎7Hb�+*p*b�#�Bv����*���?�־r�~��ح> >U�d��-߳xO�����&pc��<�$6����h�̂���l�o�+�	~�v��q��/��d5z�>��<4��������
�A�*����|�9Ҽ��I)S�y��N�̈́��`��'�+ ���f�lF����em���O.i�1��5e�w�:E@�t���"�E�DX� ad��Y=1R�P�����/�G�4�8vøT������W���T�'0V��g��̸C��N	�@>3�'{�b����x���==6�˿B$=���Ŗ����	[�MA(FX�������br�{��p�?2@���A�=�X^�� �cڥ��q8
���_�De=�9���~)0JW.�C_�y$T/G� �A�T�&' [h�5&1��Y�@�\��ѝ�cYv��g�|У�5�BeN�n�B�q��52��^�@�xߙП�Hrw�g�幍�ϲ�
Z[��4��s����jT���X��|�O�,Т����-�'b�x�F��e�l�Q��<��[�	8�m_�i�z����eaJf߇\�iJ����m�d�Q�Ղ����}��S�H@[��f#�	���tGnr����x���OϷ���y�	G���f �A������s�c���A���6���p���z?���(u�R?��L��T���8���iLk�6�]~�� (8T����snN������	�p�� &M�ۖ�h�zk�º��D����Ͳl�i�
}L�"�k���BrBF� A�h׸�k�H��
(��a3Q^8��\�����4�ڃ����a����7g"�����2��+�J<Xvc:�ù1��n���%�'m<���h{�T��%�U�;�lz%g��ό[+QܾZ��Mt��$�x���t!
̵U�b1�U���g]���#�P;�Wa��λq�����O�� x�mQ��:�;��_��["=���!J�,��#����p�ғ�\��V+=��d$��{���f�bG�Tj��=4+���������T]�cX�H��؃��L5�vHF���dͦ�7x�..u��3d]Zd�� �l~U�*w��'���ؔ<ǘ�e�n|8:�{aDd��{XNj�������C#�ᄼ<�������3�x�h�����!��u�|�\�u!�/��xE��^ˑeng	���;"�Bp�_�s��̀'{���{*��͊�-Zg��C��]L���X/O(Gs7�8�7���o�-��s&�30\�W�,"� )���sn�xE$���]\�[G�7㓧s�XH��o"����V�,�������Xp�.��倍�Ng�[��>��(Cs+���K(��'��,��<���e�J��YWq��2,����r��cZ�g�8'{f�4-�Ǽ~u�,�c/R4��+�0h�2��*�H��iP5냟�R���J�{1��^{��+��Q�2����Xk|��VH�<Þ��Z��;a(m�QrV� ���#��)�j���o��?�ݹ/�����QR6#T��j��ׁ��z�$�ϖ�AEn}���M��9�i�y�$�_�r`�3��
R=+MR����Ժ������>�ɉ����4f���e7�h�d�z�b��eg�}�?��ţr�y8����s���d?�����ժ�'�ˤA/�> c?�N� �O%R/�/c���9H[>�Y�����Gd�#㧠��D�&x9Vz�W,cvU�b��v����se..�������J[�V�%�{1��2u�Q���=���Ø�X
��<�ۘ��]n��QR�e8s-\W��^X	4HC_f��"�%���
�9�|U
�H��"�Z�ҴK��+Yυi��n�N-�xL��o����y�\X��3([rw��Y;� ��/�����rP�lTzɷ�^fCW<B���.�R��}�,���������LC����S?�d^��5~�F��i�urQǐ��Y�Ҁ&WR�����f�$%�������{�l�o5�"�,/xl̵,C�9w7�R8�8͘T��pXN�����(�tRP��y<�>e� P֪
�N����p��Cq7��n�~8d�ϡ�'��l`F�(�b��Um��kL�9Z_
�w�^'6*=��s�.�2�)в�D1ӭ�A��JF��r�Rn�{��Nǩ#f}5��Խ��c��Owk/��'�ók���=��$:�	�Ń�+&&��	||c�=E�Q<��=���^K�@�	�l]<V��w��ǔz�k����S���Vǥmq��7���ͩ�����.����p�s�`�m~
[�g�@�\���y4�#;frʑhc��V��Tw.HɽN	�P���i��M��J(>s����Z�`S�*a�0Tx���jZ+D#2Х�tMJ)�g�[��^.���m�,����w�^S�� [��p}O�>Cww�o���Ґ������;����:�w$��Ղ�-
 ���T�6y�:=1#-������p�<֝4��6��F�p_}9�����(�5��E�/W��W@t�VQ��!B*~�^ս��R�,���#���ֿ|��+TԎ��.��Y	����cS�9����e1��v`�����X��������}�RM�Gt��3����� �߱��D�b���*�2z����ϙ�"p��{�tIb�'\�&��LW(~���$]��������a����m�����O#��<t�p/��X?��4��ń��+*l�E��d�	�%5�R ���=����4�<����xs�x�� ύ`�{���~`\K<d��cߧ]�M�yy>��FسX�gR��d���7rC�����	��Q�����)�b�/>�u���������C�7A9�S|��)Ր�`K0r���8v�2�X3?�!�V�,[n��2@���Y���w N�J�Ǣ���S?��{� @�b�R�/���l�m������*NWv���FU�	�i�F̫�z��ii$Á�eGr���^����B!�Ӷ�aɂ�YI=`����' ��TY$9�ʧ�<���fd�p g�bz��5B��S^����R#��?�����;���U��v����S��G>�e=��3��D0���Ĥ��'x��d�#{�"j�b��|d'`�������e����6�'`$V������8>�I��ϖ�m�V.�6$��JY�����.E��Jm����[5�Rw��!9s�w�O֋�@������ip^�0A���D�c��7�� �/�M�?�?<�ж��%�8�����7
|�!1@���
h#��G3�լD��m^p`W*��? ���G��V�6G��L�֑��^�-���`�ښ�Ym6��&du;�}��f�����n|>~�z�_S��<�6Rŀ|H�������9[X�l�/Y�M��3{Ï����`CݝO��.P<̴1eXɔ�y>tu9Jn�i=�ʊ�/�ӯe�LEǀ���1*�qęa��[Fmt�[ݤ��-rW�s����2�g]�B�M暑l4��R�7W������?�2\�%�輳h�^��#�	EY/�<���,G���a����~�1	��6�dO�<'+��܀J��&_�{��x�&e��*�k���O��a���|��%��I� � �������Ӹ����PPpe7���yj�y�+�� G��$M��ϼ#�X�s�Kϓ���;6Y�˱iO�@�	��� �#-	-+6"��-r�Nې�Q��/���*+���wp�H�~��Se�B�?y�յ6�WUe�'��ۂ�jk�m�p����SZҍ��{6���7X5�v�)s�9��Ж6�.��!�=o��G:*e>"��R�����_3O*v��~&���%;������z�cAtlj��L�&xg�H�f�+smDۅ(��<h�,��+X
�z���=3�Մ�6��Cò���R`�v�dB���|�'+$�*�u����UC�Gmք}>� �hq��mK����O]��ٛ���[����f�cg@<��j��`\i�g�YZ� ��e�i(-J����m']fLN! P��� ����|P��h=+u荠�g�L��i{�`��:$��N�F�}�e1~�1G'��؛��ӱ5��n:`;���e)��^=j"wx%��k����Ҵ���q򈘹$hZ�PH}��7P�N;gB	�����k3�k�b�(���?A��I�1PbO>Dp��10Wu���F���t�<�߅��Ė�/�2�΍���`�|�o~76������ߞ?�"
�.L�]�<��a�AB�:����.L��I����'km��'޳��gr ��g5xZ^�n�����vIθ;�B;�?���"L���:��T7�����9W��5eA�C�0QP���8�*ƏH�at���م�	�Jo�3�ZwMj��ߔң� U$\��+�ͬ5���,C<)>-���V_�i�7^���Z�T��d��{u����5$��B�,�+��D����鏕��=]�«�����c<uJv�����/��{<UT!sĆZ- �����ñ�&�"���;�(P���QK�2C�q������Wv`4c*�xF,����4l��܌XG��U��v5��+_O��Q�&����Ǡ]?�n��v�΂����@��Yq���>��W��JQ���Ly\�E�A�j/�L�
W�����lHnŚ��K�cr5�r�U��wK+$��J�$�����v������,#�l����[�5'C0��Z�54*!G~��m�ظ ���SR�[Y"�Hcd�sW1Wa;�z��2%��*�\�������#0p�AF�i+����BM���"V[�L�LFs4��.�|V�A���	т��i^m�0�I]��$I�B(X1�#�,�w���#-���I7o���r7բ�]X
M��O:�i�q�鞄ԯ�t�� �J^c���_�p(��b����e����6��0.	b����<Ws��;�U���x�|�8�N�٫���>���M�i�lC�T���M;��r��J����ya�<As�s��R�$O��̽S�<��lPx�R¥gJj�2d�#�ę�:3&;��� ��"�!Ĉ�[ϵ�`�Bf��X�Ed�����5ު�^K�Lr�r���lO͵��F���( H�ꯗ.ͧ��É�[y��4�Hp��R+�:��4L������	�H���{�M�Y�odz"���h�omTAdzHr�p�ڛ�qBˉ��_��� �f��V')���-?V�Ŝ�͔;	z�O>�/B��$x�^������]Br$/<��O�`����Ng}�BPh3��
/z�����Q����W� :X��a��>dV��t|��g�e��1��m�|��hơ�ēA�|�wm�\��[�����¯�
��-i���6��.	�"䮍�7pH�}�k��I��ܩ9������ǧ�ӽ%�[�]:�賭�DJڸ���u��LS��'o=d�Lޗx�� �,�RA産�W�C>ߏU���z�*1�;���n�A�JW�ip6��Z3�^�f�#N������}.+L�����D�2�6��/k������ՖOy�JB#%�vO�[J6� 6�@�m��w8���	g�_�4���^��'Ƹ3�?�}�yJ��i���]�@��#g�P�=�9�q}#��.Z9�Q^�n��!��p�$	B�O����M
�GQ�+��0J�gCb��`.8krͼ_��@�uiY�8�j�DB�}��jI�7"U�Mwp��a��5���`��?���̜��P
|�wv(�l�e��Zy�E�������c�i�;-c�Z�K��'�)��;f(H$ �G�r@'�zȺɒ�|w}y^
�4�^ʓ��&�j�$�&�UD�����|&ҵ�IאH����ZUvM��ZZo��Q��;	�x�S����[@ZuAj�s�Ƶ�w�s�3�wѰ�"GV�h`���A&��Dk������BQ4؟����ԇ��D�=߯#$_�*ZJ���T}�ّ�:5FV�=zA.��D��@��[�kO���g��������_^<uSf�Wd�u4�ֹ���_��&��u4�ZI߽�l&T�u��W�Uպ��}q����<�\Oe��=�EMBQqzʣ�v7��V�5�_i)>�)'Ĉ3$��Ý#��,�z��%L6:�qq=\b�_�'�X�����]���T+�e���X0C��FZ��Z,� U��Js˩�5�-�,�n&�:����T852G<�d�g��D���}��C��`w���D�E2#���I�2�E����c�igh��l����+����G/���,��iŋt�U͠��^|�~��E,y��Ӆ��D�7ec��qE=�7뉸�g^�8w�G��h	9�u'ZY�􏇕e6����0��kpx���g�mh��Tg]�&�+�*7N3u�0�,�I���Vء��e�eX��΢D�Y�I�̹݆3�M�[����p6�u��&�u��0W �8��s1�/x<TF���N��܄�#����Ƃ���FP�$K��wѰ
��>ꤴ� ��|x����o�y~r��+��� ���B��i�/�{PY��`A��>�+'����ѭ�׺���H�����4�1����jd�ݸ&��_�R�g
��ܰ�wC:�ݬ��j��
tʖ����$�ʌ�q`�<�(�ӽ�or�)1��Pn^��2�yw�$Z.{ L�r�M�;B>~S���Oa��rkͲx\�7 �4 .��'ض胫X�o���]QQ#�~7o�﷡xg��C��g^����h2�Be��`�=m�jN�[w����y�2��F���VH\@PR�eV��w�Ž\��Ud/547�y���g�򩣇�M%zm`%ujƠ�x0��[�z�����g"$�i��X��!�Ud���Q��;{�.^ǱK_Rv��ZW���k<�%��u�מ��,�S���uk��$G��1p��=��0��M|r j/�=�ޔ����^%	�
D_P�4f̔����ց�[)�4�	�Lg!Y�R��G �=��&��A�0��Hv���8RE�M�F�"'�
^^���8���NMzV(�bc`#�%F��.��~ο��w j3��_mA���{'����Ѣ�>b|`=u:F���b}�)%������Ψr$�29����[�:��!�w�L� �tJ�~,Ɠ�<ZG�0j��Ӹ�'��~�·���DQ,���BI���8r�+b@�c�_�≛$�r�����꠽��I��[���0�L$q�䪊�y#��4O�r�
 ����D���@E�����{���G���G�j~Qd���� Q����J}��yJXf��M�pߑDa�4��%�J���:�}#zŴZN<1�����x������  �8$v/_��_��}�-�ҏ�H2�}���Uv
Ǻv6Ca�5�as�:�[��H\˙�s�&�@�<��U�k�>1��I\Ε���io���^��e�n���������ɗA��|�9�2�]�;f�9�9�8"RZW�$������+0<~/�YR���3����X)]\��BN���	��z"e�-g�zW�tS2�fr��Tz�?H|�'�[H�!�щ�^��m�d�P& {hIP.�� �b� �gnD�8�G���lܵ��}YF����P�)��͎�oBiԜQt���*h���lʺ�ݚ��7u���pNI�p�,�|ⓥ8�5uS+���D4?�~>k�T�@^w.�R��FR^��H�q��D�R�4@ �x��Y��n��v�H\�g$8�$>�u��"�
�j�z�_�G"e�����3��}X�qټsj���3Ll!��TX&�ߕ>��T��� �=�߄_����e1�n�Ƣ��-<x`6ݶu<�����B���Hr��h�q]B�B����+86��r��+a��;�*J*�#|HHQ\����`�/��R��H��n@���#zt-�>=%��a	p� �_�i`��+�Y�1������&mUZ���p�Q�/�&}���6n��tά�?,а~ߙ-�w�S����ƕP�)��6��j�@�9�r_!�\��Q�c+3��z�>t �H��!Pz�k��3�ΊQ� ��ֱ�d@t�fH]�p>�0�G/8����u�n]�+`�5It�T�r��' $D��]f�
�Q���V�N�aXF�J�����	�Ѝ��[ۨ�(��.��cW��A1�%���~+�I�����I��Ttt>u����ZN��~C\$�x�6:����n�j/���O�*؏�Ls����z�W�p0zs�$G�(fg,�4�?LfE�¾����8��������gB	Ew��]=�x"���5�r��> =��Ư#5�f�I��<��<�q��
��堒�]䳋�F?���3X�:!���8qCn jfit�߽$g�D_��o�NS#�屉�_%�".������5K�y�Ж'R�m��	�#��@�&_P8�!�[p
������@��[�)���������3�k[�w�1�I��ȥɊ�W���������� ����e���c G�����ܠ�:�Jz�BbA�{�imY��3�E�h�td!x�4$�G徛�� \�3��y�u�	9����JkSYD�>���k�k�$5�m̈́��2MJ����Ag�c�������m���.�W�5C9�28s�?jI58E�7�<'�A�u|���c�]w��RRFa�F��&�4���/n�^��BAلrf�t�q/o,jy&�dd���G�Bh�NS7cJ>�n
&#�(����1�y�⿝�23�Ѻ��x&��i�
z#$V������H��$�	��W�W�_�8!�G�7�,ض��d®��tT𸧖��L�a�:��]�,��֐1;o�e��`�ez��4��F;��:������!�MA�AWͷ�v�ŭ}7&"�Xqu��wIW�����ͅb�k!����i]����^7���(�>�9L{����}>~�+�'9c�M��r�%@0i�Sr R��@�=x�Kg����C��r�|��B��CZf%�s�G'�C.�^	h�!��|j�cS����ҵ�M_*/����ʯ����=�,�nP)$�'^j1mD�E��z�*��Z�x����HG���}ܛ�N�DmY�Pq{�� �r \��I���~		�3X�`&��
��^H��K�+ԙ���x�0���P�y��pP,��;O"6M�ȃ�F�64rLj���@��ua���#��s$�f���4Q�{��-t���e����/Ccѡͦ�; �}x������P0cY!KE�YPH�_+7 4܂�tt����{�^�4&^��z �9U�c%�U�^mcI����[:�RD�Ƙ�\+i�0`�;@ �=�KH)�k�&?��@x(���ҝ�+�ޔ�c:���ޢx�V����u�d-Hl��z���Ϗ@?�x�ŭ�����[�1�8팽�9�֛j�Oټh�G�0wW�;����e襼��d)�]��������mF!8�cE���cRKۇZ�:�ԔC�e�s�^�k�@��o������I��B��k јҴ�$B�3ħ������Ŧ@��VL8"�NRe�,��q��M�5�{DycY�NU}.�J'����Ӫ+�J�&��lV8����y��,d�w�VіH��O:%�nZ7(��Q�5Z�%�����r]-��w��p�m�V���V�F�D�!B�e��y��S��2S��'���Fݘ�gs�&�8�*��-�:�V{c%�3-ES��<�jN���t$���tH�Tl%�Bu��A�����R�����W�Q���HԊ��)�H����c5EB��#߀~Y�6��_u�s��x&�﷗w�Os�\(5�li��D�;�BbK*/{�iF�bzy���Z k_)��t &s���f;ٶ��c	tm�-�L��^��S������"5G��1R C�x)?����w�N��������<ڕ���?���e,r� ��ӵc�N�=��:B� F-8�V-֛�:4��/]��Æ����JQI��_����΂�89<�1m"-��lR��P��^в6U�?�x�ݓ[�[O�p͚�T��"��],|Q���
��Tj�Q�����)'!^��԰�Ĭ���*/��d��C6��m�D�z9�]0��:�|����X�C���Ca�Pt�9	4���-�x���`����Zb6F $�	H$l�D����{D�WnS!��Ƹ��3�`��T���Ns�e�wO�S���'�u6�ۘ�[��f����1�kI|�5+�OS�4��-鿱��?xn��j&�����,�=�P�'�<�/1cU�]�WbQx�G2�^��t3j�h�f;��j��p��eccζ8}��V$�m��6�"�(��;[a��1<@��v�P'�`������zY\��j��e?|��+�+{�Te��j��ı�r*�ū�ɰ��:�|������5Si��>n��
#SO�ޔ�NW+�cK]�.D^vg1eO��Nsz�k:>@R?pZ�$�PD��>jߎ0hW���U)
(�>�/}�//�B������ݓ�)��3��U�g0��d�W�w�co}��w����i��PRڦ��'}���E�VS!S\)�	;2۩�H1��"�� |Z�&D�z�.���omLj�~%#ݿ��{�a��dԎ�Eۈ紲�R��lA\^�AwL��������ŭ� ���ro]W���qح=D���j6�����	eR��v��6<�}�!��KJ��\����-c���om�5��HG�
u���xxA���y���U��.RYV��c�����vsQ�Z�#�B��n�/�8� ��2�b����}@&aى��Y��Z�Vo��F7^q]����X�:��fj��vw�=��(��0X�Ђ	ɕG�p�L-!n�_�8!�R!���U'�Uw��L��-��J��E�	�cNy����u�`�-*�>$ܳN��W�����?o����Ӛ�ڽ�\���n�W�$7Uᇉ:F�X8�O����F�#}%����y�+8���U��'`��1c�qV�{��]0� ��
sz�EטYq|_M����$�1�B����� ־�!��D*��4F��dP\a^����=-R�|1~M�u��Og��"�/f�.w�DV�N����I�b��n�r��ʗ؉��L\�h����ܚ)��A������)π�������('lƲ�z�_.���x&��}^�\�5�F[���Έ�8PTK����ި�D��Lw� �VԹ0�Y|�����0dz��s��߸P���P�ũD�	`�����D�+�qȪ˭0���͠�^�r�����}6�J�-��A�*d�2D��	���܁ߧ��1�>Γe�U�⢁E'��{���z�W�u�c}��`�3S�_� �~`^/aE�WԾ��H����L�8:�ʾ��q圯3��F/��E�.H�����d7���aƔ��RlWG���>�?,�����W�����/M���+�e6_��Q�?��*ˮ����ȶ�N��+'��7�#�-����I�C�������Q!���u"���7D;�,�xJk7�ɍ�e�ω��)�z[/�>$���՝D�(j L�7��O3�xp����A��VT��6�����zv�"N��.��������E8�M��4�]!��B^�֕W����R	nK�I��k����c��!�^;��fki�'Ϫz���8G��
쏼4�����AhD�N��F�lcq*>�Z�g�[���+��ߕ��L��{q!h��pi�����o���U��O��I����b�zHO�(T��#̊ f	s�"1�q6	t��a����>@�!��_q���i��_��(6��x]L�)������^�IJ���ld�sN%�'3z�3	O\�J�S	�X���T#38��a�nI3�h�
�� ������H+�X�o�
�m�(��l=�x�ɠk��}Ƕ�7P�(����}DH��=q䉊�v���X� XO��sc�CV��/jB;vyz���M�ND�+��/{���;'O�K#%|�C6ٸ"Gr��}�]�1ٟ=z�A*��>�Ox{i���iW�$�u�L��ui,q�X���8M�?*=��/b��A����D���07_^�K#���Uj���������S��s��E���o�L�@ie��8A�&�cJ3��'�ԇ-�8������?ODm���	k�@njm1 *O�s����չ�K[�"�1� ���9����ϵ=��d���TK�y����;�`
4���!��ĺT���}W��)��`�s۶^�z��%~�����V��Ăj<�a�3�:��5v���gT����"��#��C��N�b��|$�����'�j\6Ș�܌�w��KX'�qȠ)kƯ�=���w,Nο7�Ʃ�q��̟QXC?%$A��;q4�l�r�_q�B>ޭ�`����DM�猙�yb;���\ ��LHl�8U �=B$��Q���L���c�>.RZ� ��q-��рM.f����^E��H͏ӥ9?�"�d�]�����s���OKW��H�,�g�������p���`�|�v��2[M�[�eM��dh&�e��H�
'¿[� �27���,K���v�7Q;�0���~�eUJ�fe�P�-����$pk���)�)bri4��s���8K��U�99�d�P6y�{��{�Z<�;�e�ԙ�ۈ���S|Y|�mm��b�`�j� '���^
6Պ�]��h!��L���qʅJ���3�x1���&�/Ž%ǈU��BpaI#�'�6r]�(މzڧW?��ϩ}�����	\� F�8�{ܵ!gUE�Uc�w�t�ic�;b���X@�_4M�N����8�N�Ȟ-&n�Pp�nf��z"�V Q^W����>���*�!��t��S�� �-Rм���9�2�
W����8d-��F�_�Q���yi.q��1Ղ��g����Rp:n?4�$Y�+J���-��'�Y�̻#ץzFZNh�~ �P�U���2�Kz�(�=I��~!t�7�����CH �����,�e�Fa_�L`�$�m�D���IH�q"e�{b��8Ue��0�������lE����jo3=y�e�OT(���ce��œ
�?-�n�Y�sɖ����2閽G�(�2�|T&��N��S�c�Ǽ�:�p�6�����;��>'�A���z�aUBI2ڥ�\ �W�n��zk���[5a<6!�+�P?[z�q���%m�w�AT���'��Y��f���닢��B���B��)��s�����+���L�a�n���#3چ�Ea��Άo��Vp�p����ǰPY
��x�����������C'FP�v� ����
vtK���E}�|��(��/[�򑂧�P�^3b
�҉7�f0#�qe�Q^s����}�:�.P"�\fQ( D
��F�Q��@Һ��^�A6c�H��K��>�a̻ɳ�"�1���^�1�{ ���}�)�� hl��[z!IA��7�k��[�����H���1���V��C�jl�����7d�Pm�~���=����J5�4qv�����W�~E�#;��s7t�gL��%�W�"����I&<c��R���r�Y�c�/m��S8��8�i���x��X�E_�Z��ΞJ�Ѽ�I�#�E��V�ƌ�&���9bލ1��Y�H�</j蔝H�;r��;̤=�I0�T�N���Z���Lb����A[�xer�5�]Z�M����Y��w���bN�}�6�pѱ�XfK�����F	�"sl3�ٹ��o	�QO���QX`Xl�`�*�>�S���PI!���3�76ǝ�e��+d�K�^%e Gx����>D��wvbE��Cx��-L(���<[���(Y����~�T���{�P���U�C�2Θa
�\���`%b��B��v$D�T@$q��� �P��v����T�G�ɭ�@ZX��#�W����&78�à����@(Q1���r���ӏ�Y�����h�{�k�)E��Ǿ�J���9;B(�בl���A9� �%H�3�R���[k,�V�Q�����¨�'�k{)l%�n��":k�؟-����^ .�H���J$���������Y����UL��`��b�gD�Sҹ-<"m�ǝ��Ī솓}������2�i�4"�}��όb�G��x�?�|��BF&�ͱ�p��&>IGƭ"}eԘ���N,%Id����ϧ1J�,�+|kj�]���C�pn��f�]<]\�"�n	����/�r���7����|�G�,	C#�x!��4[��-�kM0@��N���6cp�3�0��ܩ6%�Ki�8���ܥ~���2�����j���26�>v�)թ��sp���| �s]�j���z��|I�o��xO`���q���p�x��-s�8���:.7�
T�rZT�5��QВ6Kv�	5��Kp ��%2�,@`�k�Ǽ��<D�ۥvAKu��J��<5�.|n�I�e�{�ڏ��3�G�B��%�-4����7�M��֚9^�b�a����%�|Ѻ���Ԅ�~LR�.�Q����qj��Y�sP�ܔ���\º��iMW�Lh���,p4��FE3��>&nh�i�hSk��W^h��)-��H2����4���r�`!�0�<�$Z��b��E����B*�C��.�
AXwZ��c��P0NƼ.zg@ �Ě��hΌmf�V>���J�������)�?�F��5,�$�*9�m�j �)��z�F�����UQI�u��r��ώR�R5�Vl<�ػ�^�F����k:p��\��l���1��j-������~<,�1�#�e.u%�r[��5i�G���m�8�rݸ���M�"+�A��Ts3`1�w^����+�^�2�,iJ��[�a�S�������@�M�ߗ�@������=i�K�GG�jG�8���I͒�"��b�������8e���z4n�P+&w�ǁm�� J������!�����j���h������۱��P%���Wp�ؙ"��?�,ж�q�z�:�:��)ť�g2r�*���\���+��`CH�7�X��׋�n19�I�bU�����$����D��b �M��d�{�H������LU�vH��梁�'(�1�r/WL<*P.��ώ{���!�����pc$R��Lv�0�c����}d���Dp�U�'��� �2-%T<:�5���1��yk����mk|=����]���¸����<#{�R{.(�P��YҸ��,_�@���v#t8&-V�%6���׻(�^��e�JO"XǴow��D�0l���=x�`>�u{��f9�?k�����ы��v�8��o�I�&eNW}6NO�c����^<)�5=<��"5t"%k(�蚲�Dm�B�<�,�1Cx�!�G�I�<R3G��n���r���h�:m�b:����i^(�׊(m�i ��9���<����o �"5(5�>������h4��{˾W��<����=�F���q�E3��h	�\�F�\��o!K_�eD�{J�o�lR�&�\[w�j�����ȳ$��H-��J�6�1��w����v�5���_����w ��"U�>��kl �'�n`(����%��ۍo��%����j"J��K�����	~��lPR��MJ�/m�9��ֺ�9ؓ�)t}��u��ҭ�U4TPgU5���X��_X�n�/�y��,ӛ�P��¹����������j�b�>�P¯|/�&���<�f�e�Qb}�ï�X�{S�ZE�q��8��,�H��Vx;�d�'���Ͳc�iX�K����.���K����F.�>��3�0�L1+\MG#t{���wU��]�!��� '�/^��HH�*�+��s|)�v�7�[Z�Ϥ�~��X���ܢ0ڹ�Q�������c=�3�D�+-�e��8�T�F�Nٛ�6����|	�}���Ã�
^L��\F�Oy�d=��K��߀�
噋i T?�T$̉Ԥ])]������!�I����T���!����,HV{�O�ŹD-Z���8mk@ h��a(2�_�'Dʰa�3��2�1�W�.Q��CXMa�Z���i���.���p�Dh53d����b�Jgz&�}��p����<�P
�nn�5���ϝ@:n�<W�'�\�%:�~��m���l�����=Vf������D���<߻r����qY�(?�:y	�Dor��Ө��K�}C ՞�zVJ]��:���
͆	�h�sg�:�#��`��,K���5$ˋ�q�~0�t-�1|8���J��_
��?Pz�3!�Y�|��"G�8FR>E5�3CE�J [�jܝ��f�sG1�'���q�ԉ˚�X����R��u�:�G4��a�JA��R=���k� �O9(�fp��QF�߷�ӗ�2�O��wb6� ڸ){̑(�S�	q��=��#��.�r��j�V��E�1T�p}f�O�u����~����$xH���zY�цg�<�j���5��<�>j�E(�/bt�<���n�L��%�:��VZ�F���$A��� ��e��=�z��w�����*�Ǯ��k��1�H���!B��R������������ii��9"��X�,��>�%�c��tr���yFD��85�S+����ű_bp��ޑ[#x	.{�\58ެ��t�6�/�](3���MkB��Z�������QF��?�q^�7��:�D��������H���@��)w8N%��ผ�B�c�Ԅ���m�V�C��)se>7���.��Y�%6�}F=^ZU���I5&�"����[�;��}HQ�9�zD�U���wK��9%��Z�_�x�f��߅z�NM,O�gJ���p������
��`h����,h��$��7�X��^񨑷���8o>��R�C�J��ݐ�^���oa����)��_*ُ���!��୭�P]�ڛ^�����Z�ź�Bp��g�on��QO��)5�Κ6�W����Iİs϶�݈3]L�{����f�_�x�qQ���#��.�k���3`V�o����d�����Nfڿ	���`�U:4��	rp\4Ʃ��,��reo�u�<�	r�ɚ5�N�xR�>��$�Bѽ�Ӊ`L-��oD/��\����A���í$�L�{�S�J�V#U��O�C搥l�{����pwe��x"���AH�X���G:�1-=/�ܔ��C�1�v?St�7-�F��*�H1���L	���I�#�#�٤�;�,3� �y9���n�@� 3����NF���릅!j�wr����]?�He������lE�	D]h�����$�PtbE��G��_���ʣ���;�
v&p�O�^1c������Cψ.�uy��G������ �Uʍ#3��vb R��RU�%ś�>2q��1����l�=5	e\�\敖XږM��~��<�E9k9�S�����;���SWĮ9O{�ϚPQE���h�"�˒/m�V�ִ����*��Q�Z_�6��$��Lq�	��~��\D���a��x&��ţ�
0����U�<ߕ|��n6"��\<���*h�j��U*��,��pR������\��+�W9��Z�e���^�Q�w^%a�-��̓X��5��g�@t�@��NR�k������ ۸���U���r
�d����i�7�z�Z��^tϡL��4�xR5ev�D��[��^�缥��$��:�����us�ާKâ��t�~M��&OI��9a�Y�d�l�dV�a��4�7�y��ӥ�T�o����{B�ҋ�_�ʜU��k�,+�?𮑛U�i�L����3�/|�D$y.]"���z
G��λoy�)���\l��A�x���{�\0���D.�4������y���Xc]A��݈U�!�U�O�� < PLK��� �%��T�������ꚷV[i`%�N~�L�r(�;���§�_�4_��b�/>b�Q�!;��W�_��W:2'ǧ|����:���ӓ|1F\����Hw$��<Jnw��Yxe�M0W���x#��B��II��V�xt����F���p{��>#�ȃ@��*�u�s� ���5�H���n�&]��槤�{1�X-uҞ��i?�3R�)�ĕD���[#��s§͎�i�{ב��+��K�������̫k�Ǐ[%����`(����J�$����bёJ��xLU���E�R��r�YL�/+�U����>P^���*BN���D d�6�궦Ã�`쐊�s�QUx���,�R+��5$x	��Hh	*Ǔn[<+���S4P"�B��vbkތ���o�i��[B�&z7�KLm��Yk��!��Q�A:���9�Z�w�ـ��Y܍��7�����E�D��;� mH����N�^ɹCa�^):.��~�N�mx�|5a};���1H.pY��i�L���au��I��v���!�Mk7��a�� y���w{htm`H��<�6�J+�����H�,�J_����V3���%�^k��L񈊈��V���d�5h�&�ya�d
_�Q,��F��u�Kķ%��Xma�p��vw���
��v_�$�xQ��K7yV�X_-�Z%�,DJ��!rڳ�$��E���\h��`��3�=�� y������rőԂ#<�_XQ��ͅ��C�x�F 2����6\���u"��M�־]k^_r��������G�[�H���,��Ͳ��&g�@�Z`Y(�K�C]~R�q�D����Dq�� ���*ڂ�gJ� �? ����ؔ"��0dy]��_2�o��$�����Hd�13�J���I�c��d�xW���R3�0W}��I��Ϣ�������^K7��ÿ
϶d���	�[
y�k��vo����D��N�[�u�A�?j?�[Y�ȴ]����9������v��}c�Q�0.2z
*�}uj"g���!0�э��Y������i݁�W�K�(J�q�>�X>�f'�Q��o�g�LX�2g6g��}E�E�V���-��urC"kc1yq!��8������wo�3;6�}b9+��{%�
��ݚ�v�Df��������j�Ŗ8�;��"��b�k<���z�c�t��>�����{��@(�[�s��<�!�K�*G��6����l�,^����fx4�u�$qa8�Hzq4:�����m�������;)��`��	�·D���_�Rl�F������1������6�/�C�4� �ơ�e�f�����}�j�e&>�,ńH+��,%E�Ҳ*�i�
�.,�`�l���H|�
q�ܱ��:��Yk��|Q�K!&aX�l�@��n�y��{��%��X@p�S�q?�q�xb��|�/E��Wf`X�:/atؙ�tm��͖O·�S���<kή�Q/��fG��T��#�j$�\A:z�ާ�D�ӂG�X�ɶD�#����R�se�1b/�_p*:R?6�z��z�$�Ut�5�?�~���Dj�����J���ʵv�p�u�.�Cʽ`�g�N>y��5�� Q�����D�Xo�L������6a�~�.k6�]�sA�b�-�f`jCxς#hڴ��%�O9�,����?Q�����}?�(H����Hf���.��F���Y|MZ�w�TKӇ�.񈒵��	Bz�R&)�BDv��pê�H<`�;pu�w(�&C�v�����t,^	~#�h���G�G����'��uԉ7�C��}�U��cUd�1��xR�#��|=&5�A�%\~�G�/t�=A�KV�S�1Z������7� ��q7�
��/�h@���-�ed$_kSa�r_�����=C29�-�sL�1���v�˃oTt����ϱ�����N���I�� ��H���?8��6ݥ�vd��f�^�@��YT6l%it�B�%(�	�m��Η~�>�5�4�ؼ8�'f��� ���}i��at�E<#3���4�8.z��y۰E%�Ci�ڎ�jggE�������1�0�?&�~Si�޼�1��%b W��'�@K�O6�X;�An獮tg�_"��϶DO���-�V��.�vU`<�{֕c0R�``�4\+xy⮀�6r#p5|I��SZ�l��l^��$N؝��6B� {�Ǵ8���s�
�1��D%�{ 4�)ߎ��b7|��5���V*��C�z�?��G��QZ{f\�5I΄#��	i�����w����o�?�`���q��5�ę�.O8�� ����ʄG���8(�%��](������F���~_���juH63ց����m��<,��!~�Z3���>8?�:�?��D��m#3b�绑|�ʢ�-JS!�V��숪_&ɂ�}�E���F�Cʫ`+���e7k�x�'B]iK֠�u������
ABZ��j�/��6�A_�'K�BSQ�˾��?6��un�0�:�`�Uf��L�yĢ�h߼����� Y[x�|x���c �VJ�;��~�B�ֹt������p�qK������&��m�u���7t�g#�H���^�]�3����p�Q��j�EW6P(iq���q��ܖV=�@tq�����z�d�Rôΐ�&�<P�Ml�¦9���P�<Z�Ј8V;O��"aH75bP��i�r�ӕ~���t�ɴ����o�m�����[g��)��J��L�����F�H)��9`˥>�:���_ υ�-[�Ł[��+, �3d�_�����"!��'�U�a~u����៨�v����j�uG�)p����Y�b�y�ρ���ě�C;y��T����G�y�q���=�aAi:�MT���� t�
d]�~F���k� pN��Pw���Z�7Nq2s�>�#���T��F��u���s4-p-��,@����yዙ��o��fO�B����9������:T'��E��R����g�]�v��6O�FnL$W%�$�.���?W+3��C�*��B�=u��sk�Jm�N<R:�R=�'"�����:Ŧ��kD�>�����u�ʙ,S�%U�M�q*�P����Wd������3k����{�Q'�N�M��)e�4��
���'AO.{M��oĹ&k��/��4��'`ع5a��k:�T�^T����߱�-��<�\MKzKx�.����s�Z6z�-RdV���ኒ���s��jw�P��o� ο��C�i��J��9��8�3��tY���V6��^3	�3��h��P��\'0,T�ME���x(�!*�1���ݸ��q
�+a�,����dꋉ�~��_����+=��4�B�0�jZ��\�!��U���|�=��������=�	���Cd@�1�Y�U��r`���
�'�������\��]ljG����q�(lȘ��Ʊ�0iD�E��7}2Yչ���df�Y ���*�n��0d�c�O&H���v��1�5�$��&�-��oZ��"х&�L�`Jnkp�L�Dtr�7r���]@<�P��Γ�a�j����*��4�B�{+|g��p-��W�CN�ƺ��PW�[�M}���: X�O6AO~wu��hw u��˖t{��DH�YU�R���h����FYTe���Khk���&��ѱYHJqM��T�
n̜I�zX�)A/�̘ӝ��<Po����NM�/];*�c����s�l�ng)yMT����W���ezτƜ����4@rt�)�c��*��8+�FO��,Gv��(ù�+��d���}�2���EE$���XL3$��1��yKJA��V��ㄐ).�Ĝy�XNk������wn�<�������?~��m��zd��3�.N��jO�bR��Ǧs�벑��Ffʹk(�ɰ|�9p�EE��9K[�Dv�YaP6E�T�����XT ����m���KT� �>�;�8�W�VpoS���!���tP?I�L�����rs2�f!hXnr��iP�@.��+ �i���SL�"�A�� ^�&�?�<���BS`��/Ʋ�luz��C�ȼj!=@a�����?�����O��Axh���_hx��8%�0�X	W���q����=YA��Pj%��/=�N�<��e�Ǧa2���� �óc"f&	=;�B7:��E;�	7�Z���,�C�u�$D����|�.�o4�����]K�e�˓sr�fv����h�y��y�=�u�י��4����\��\��C��1j�7�i��u؂���Tc܁���Y���}()�\"��0K]h��,{ *��9��@s�*��z�n��Yv�?ʬf��Uǂh���{=V�b�r$�,��R�(l3!E�p�6N|�6�|����~�4$V��wSaFl���g�������_n�>*���������{��v��9��TAt2؏�6�!��mI4	D{ש����x�J�U��2�Ǫ��{\� ?ȹ�u٣)*���7�Fb�&@�fM�=B"�c����5^��v��WG}_�������k�łΦ��m瘙7�L�"P�1�f��$�9($jl�oK�6�|Ą}dۏ�iw&KVs�P�'M��B�W��_\A�O��5�%!3v�_h9M�(��u���I �~�S�U��$���׋>�G����ţ]�m��k���k��̨M�s`�����{ewɖ��9=� -���`F)�1������!�Iˡ[t��چt��)�Izu���\��!�l��Ga�W��,�&P�e��9T8��V�{N�
hԣ��GJ͹��T��P�.p���4s�7�|���^��og-a�F�餰�,�9�TS����QX��9L������_�)
+w���g��O��s�\߸���|��
+�M�Z7:g�!ԯڑWYۖ�s'b���孂$Ⱦe�K�e�B|�������0f{�<��wdi��B��G�o����û�^�ȭ���]K��E�pWg6�̺U�/j�m��h���q����!��J2�R`�'9���c5|�S���MDQbx�[��S�6�}|���g"��6����/���D�c��.�ut�b���U�[Jn��I&P?U����h�� �;3��lHT:��-�uގ�,��M
�9o�L���JT�����\'�ϋ�F��9��[r�=�ؙ5n[��16#*7H��K�&,V�E��8$?��
�`$)Z.�����2�D�x��ic	�-$��_paĩ��x�9EM�	�J�����XlY.��X�)�ϸ}�c!"&�=����F��[s�=֟3�� Um(ڋ��Ov��]�?g'����k_�ǜ��bGon\Y�x�����V�����ŀJL�D���&�3fh�9�G��L�9��>��UJ�$S��o�U��H�v��j�j�����������5�9ɝ����c��Uh)k`�?�צ۷�O�����SK{)ގ��k��i�m���*p����tKJ�g���
�˸��X����ɍG�A*,9;������
�m|�=�g��l�|��E6��T�oK�f���9�b]HSHPct�����Ǆ��e��W���f�����)�1���b�2�b��ztE��"Ղy2*rv� �o�KC�Ԁ���o"yW�os_�m��f�XR@���G� D�oT+��g�H�Dp.trG;��Y5���?z��a�
��1l���1זº�A����]��{������,]�m��iH�j��4�����9Q��"do�1]jM����n�{QƔ�m���C Fu�l�8���f���v�\�{df�=�H�,K��ٲ���k\�me����&T�Mxֵx8�#��N�B����k��m}�U�6�`���A���0�Y+x;�+Y}T�b1���SߺOe!�2�U��I�Ș��u9�[Y�])�߾���N}	�j��6o6��L�����=�'y}5,[BvЊ��ӆ#!�ob�Zxh&���҂�u3���oʸ�����U8��Dl� [9���x���gfl��0%b�AM"y��<k_�xο ���
�9(\.��_\)�y_h��"����"�����&mvg��4��i��/�:Pc|	��UXѐ�:��hpv;�YX�T}i^��O��~z
�G��	�M�6X�,���y,R��&���N		���{2�1q[K/��-�F.;/&�n�?�Y�ĕo^:vs��ـ1A��\���vR��J�[��`瓊ιsM�8y˖qW` Wƹp{]�Tw��:D����K�X�J��Б����O��sEŸ��`���Z�Hи[�8.¶[��K�Ρ/����IJ�d�k�̀$jof{:�L:���Cҽ�}��n�x=a�'M�z�uB��A�0SJ8�TdU�ɼ4�#�.��H��G2�x���������o�θ���gL�J�%�;�7����8��%��z�)�H]>wy��)��HP��T9�~`ь"M�o�a�B�|�;��~�u?������φ�9m��Lk�	{�z�1f� ���YT�sLzB���l�T&�$��L	�{	V��F��h��d�~pw�U���5[Մ�`
N</�n����30�F���#EutQސu�	<9~
:����v���Kˀx�F%���U��#mc���k��'�f7�w~}����t�z����n��m-& �߯&#�1�Vw�A B�؋(��n"��ЁI��B>V�����ILfϬⒷ�OC1�pC�p1�y��_�'� >�ׁ;Җ�!���P�5����q�XT�*�i�����Z1sJL��]{��0�.d���l�t�2�܅�,Z�	�Q}{!RL�aoyx��id��{��ͯ����i�;�J �!y���)��D���8�c�ߛ�v����O�����=�����0��9S�)X�"��)�U����}�=><}�J4kĺ��[A��x��^�C'�Ƿ�&�YS�Q�q{H�EH��o�	�2e�z�3��N��m"���$�돻����ڶ}�1�f^�k�[�6�ѩw�{��w�wQ�'�Vݹ�N8TX٩����b�[���p4~��V{����x$kI���|���=C�� �,=��������;�?Sub�+[¿�0�H��Ƈo�i �$��e�`؇;����!+ٺz����;v�VjPD[5��t=���X���L�[���Z&~��;lRul��@���KӀ.�vq���*C��&����zS骡�)���)m����53���kȒ'�Smy����� M��&���E�m���ӑE��E�q���'U��h�!�o�2U��|��o�>�$��c3n:zp^��YK�$���`sW$Xȥ��Y:�禚��t"_��+n��9�\������a�r<���g�P������]T?��\V�ykt$��-Ƌ�F���L���:�k>��m�F��(��	����Ƕ�_�vb6^N�ᤛ�f�gWN��49��VJ�]���@��<���Z�h�J�|�ȇ��>4T�������p�؂��N���%r\���`.�����QNL�@�F�KC}�+S�f���2�0����,*X<�d� q}v{��V�d�-u��!���j��� ���Q굉������W����VymCj���׍����������9>��6��ySh5s70]�:H�)x�T���~D0����!�m4����Y.�4��'q�1�r�6�o��qx�p����L"�{z[�9P}���S�3����Y��4����[�ɢ%����U-�5�˹xi���].s�
�6��5�?��:��/�����4�Q�<z �z]����!</�Fh>R���5��� ��s��S
���=5m�h�	ڌ��넓�ܻ���$*~��S���G۳���[=�.S�`�o㿛��"��uI�9�:�T1CR�c�b���?r�8����{��.ȫZ[n6�U�~�u�W��d��uȞ^尹�]��Ժ��HM�
��.�U��D�ǰ�q��B���0�#Lr$'�T�����������*��j�����h7�<����O� �^1>l7�8�����&c��V�$�g��9��7��$D�9`�x:�tE�:tF��ÒUƊ R�@�!ȿ���P/q1&	j�)����Z�ę)�"�J�<���A_����4����rT��ү�,"���'����,�u�:x��r�:�vO!����1�qܣ��bHV6k;�������a%l4eNM}g�y	bxB^)/ԋ�$A��)j��T#��>�-9���H���5e�r�je�ٴ�\���= �RF�z.��`�>�X�9*K9W�y˝��-��Ǭ�F�~�O"���ػ���){!���IT�+$����w�����!�j��0��}��Q-P��c��0�VCV2am�'�\"ø�t���3��bw�L�!fҼ�蛽i�{\�� *s��q�{K۽�Zbw�>H��'��a��r��L��97&O��=�@y�_�����Ñ��#,I�w��6���2���_����
n's���Z"j�[L�v77�w%ws3I%Ű�m%f����֒��
|��F�X������DV�~�tN�l��/��h�dן���F�N�/S�m�@�/�/����8Pd:q�cz:Z�|�e�Q-�Q�{�|=��Dy��bB����y
t'�����I�(u�:US�����-�D��B.�}	g@��Ae�'�My�g���!���a�^��o����a�����)i��1���Ӂ{�+���O0�*(�)_���O�Q,��mq�l-�������P��7P!�i8\����2ư���$L��?��տ���K��c����� ��x�h��k&7��yq�\Ѧ�5DK5B?��<8�@�򱨬�[�����ǘn+��]�5��+#�l��H����?Ta�������Ъ����R�����H�&FY �vu8�d�p�w]42��U�!4�P��Ҳ5(_d�M�_>Nm�7��h�jY�z���k����7\��B"~s3����Gr/ĳ��7s�˲��	ڢ۱���t#�+��.u�5)���8���   ��h��ev�m�'sD���2���;=',��* \W<�)��껝PU����\�W�����c��m�����Oĵ�[ڗ��T�L�������[��"��̶x}v7*�S��(���7֥/��]ja��j"M�͑�ƅ��� ƔPR��Y8��<}
������� @:����e4���Ҳ�fC�u�Hy��Z�-!7m��[k�=3�����e[�� ��Brr���_G�Y�!F�~|��]7�]�[�:�mɊ����v9�_Z	J�x�-�M������#ɼ,#5���x�W��|O���e����%�QR��'\k5���L�$��҇;��G��yh�?4�I�6�����ho
����&-��B6˓��:��Β����Ut��O:��f��p�s���M�1�_��R�o�=4zn�wGJ²�Y̝�/㸸���dW���򓎔FxC��z;ք�ew���Ƀ�m�v�)5�TL7���,��&+�d)�uOlFE��j:�Hu��G�+b�����E ^w{��z����Q���|4��~�󴔮����@B��A�?���!�����g��blc�h7]F���Iƞ���@�4z��0c���^h�H=z�3�>.[�}�ζk��C-9e�.�Wn�ω�8'����?�S�|k�_�곂��Mq��r5�W[�"�G��������Jo%Eua=�$��y�QZ�k������eo����M3��l��۠�c���&��և�#Q�\7��=u
'��c���*N��{��!�%ͫ�bU���ɛ�\�
ckD����V��v�Ⱥ�Ɓ�(*_]���p{��ޥ���f�zT�؈U�U7r�k�<��l��S�����N����Џ��R��ʜ9f#�G�*�Jέ-`v�K�\�'��	�X�L]�� �݉�Z�(8���4r����k.剟p�s�8�مĵ����I(8�Z��'�1�����UT�R��'���I�	���W�v���p��h�kK�͚qѢ�q+�?�������;Vw����]��"�W�����-<ҷVE��-�a�F�:��p7D R6���(���=L��;8=h��@����Z��rV�6ph���W7f�D�h=U_x�K	}�vb!��p��ꪔ�G,�84�Q>0�6Z�0˖�]�B�ilʏ/2�U�OJ��T '\y|M���;��7Z�X"G������HL o/ lL-���ֶj��׶!�+dM��X��ڠN�|�i�����.U�G��2���ױ>)_���n�[�\��]�m��5�E�܌��� -��$��� ��,� �qj*�<�_�0ǉ�4�gڹ�{A\�&������fy�|����+RB)���G�pM~v����/�oːn}zэ+Z�d;dbӓ;�Qr�juƔ�K����)��H)��^]ހP���$�l��&��	�{i�J��Y��'A|~J�]R��A���F8Ti�'Ԧ�r���΍@�HտR����ů�6��lQ�quY�"���S|���n�}79�Ir�GQ�q]ˍ~���X���+	q�!<	S�M�	��-�����)X<��{za��]���t�V8`}+�C���QW˹p*2R&Ey�{J%;��V?�,An��1�6�vg�0�2L��zj��ib��j�1����;$rx�3��h�`���������7���?Ss�)�����-o�	�J����&J=��h�O佇Ǒկ
��3��W���K���p�r��Rx��^Vݷ�ᮇ�!�%Ҩ/�8"��?��J ��t��8C�(iү���~ւ����Y ����� jyL�A��sn>��yc�����;�!���Rj��%�l5+��J�ޚ������
��▄�+mo��y惔���5�G���x��M�_�+��փXS�^BD�hxm�� �N�cW�T`��30�\B�� ���v�7��K�P�j�	w�q�����r����|qò҉�r)'�
����-(NKչ�m�dT�]�w�P��uGr�����<�o%0�W��~��Ã�h$c���9�����z�y���J��'���yjd)�E)�T�l1�"<��c�Wچᅭ�<��8O����?�5��D^�J�!9�I�����|�a1
^[�jR5�E0;4����#�`��J`��t<a|tO@�d �@E�S��ϒ]e�u��\�}��D1�������=@@���?��Ȟ���s��eK����|I�_l݋q�/#�iqq�g�����GG�m���������Z�+A��}S�mD��fF�uĈd!�ɐ.e=�bt)� �vV���A�:۰���Y�V �d�<�esS�f�m���$��{��S��}_
0{l��C�XDL��~���;��~yr�CS	]%V/(�c�C�j����2���X�@L�TA�����nM1�~�F���c=L����?.F���}�+��h�*�k	/t�:s��j	��@����7�t@Z�0+�G�֣I6&߳�/����gC-� ��,��V�K��$��{%�wM�1b}�Q��d\��z��ضMXE�kV��L��E��Ir������5��z�غs*�l��N1��F�- c�˚T�֐#�&e~]�.@���*S>ëFŝ�wx�e��������r
]?~�]ː�HlC�ӈZf�;���s�P�rΰ����i�&������h����w~;�A#g�Z�E�{ILh�M�ܬc4��_�	��A��MQܖSR�B�ڲ3s�Ŋ�6�����"]$��ť�#�����I�j�!�����I��p�j����=s�Ň��"<A��e�?��~7�U@ �f�l��(-��H����t�`Z�i|2���s6��3ރ��0N3�e~�z���Jq�c�q��Lƌ������De�^^�I���wWױ՘�����g 7t�׳��Aߨ8�t8�NO�P�Q�*�3F?���^TS�T�Y]ת3��_�H�ځ,B�	0Bwh�b`�@O�tҍY�^��f�C7��˜�ߙHo�� �_�Q���#.���L|(9����G�������z)�"2Uc_��C�ZU�o�:v]
���D��jJg0�vQԒ Qr�/�~���:�����x�{�;� �b��w	�X��o�=��Żo�i (Iϖ́��j��	#(�)��Ѐ���J��~���-��l"m3��Ìhd��V4a�����簆Pfԏo�`���C����<��	AKb�EN���Y{�G	$�n�����zQ�l�T�0��n�����9P�M%��Wt꼳h�V�uG�`���wE.�w�Y���{\�B�9���
������Y������j`��#�-/�hj�m�����zE�� 	�GҤ.1�b� h�а�􂄲���=�Z>�uh�L'�֩y\�k��V4o.�Z��� ��w��L������׻��Έ����T{��S
���CO�Ng㛾��V{�a(4{U4�Jv&�e���`�C��iD�
�!��t;n;Ǳ�v���Mk�͒d��K�T��[l�bu�ێ}~t;��?�~�[֐������$�������r���M�KKc>}�>{�3�0���|��ƏNn�%���N��t��#tv�&;hj�0'"n��~[e&q�3��싟�6A�WM�5�%JP7"�B��(��"��Z+��^n�Rӡ,\����� ��x���Á����c�����H�-�0�l϶M�v3jY����*~�*�>_p�K�2P�����[c����.�]9ٛ�	����j⿾���)�x xyF���s����Y���|c�X���t-��M��e�J<Tr�?k���u=֙�"�\�uY��t%�Ne��#�/k�ws��!��p�Pxb�!N֥1����X�l%}1F��ՃcƑ8�.�=Ô�"�$43>vA���k}q�x4�r+����aI�&q�B��(���(�����/c��xs�d�9��î~��4�L���ű���[JP)w+���]����,�܍�-�D]d��f�. ��7
/X�&�?s5ߺ�?���G��H�.(�K�`�?�{,���)��vD.�H<�R*��ƴo��朷=���=�����W�]�N鈴�RD����E�����L�q��&�$N��Ӛ�EZ����<��"wZ�[�_�6A}3;�5�.T}+���g(��J,�%�^���*RW��HsC�σ������tCD(Y��;l9�D�O�"�[E���)�w��]��F�0xQp�e���Zo�
���y����6w�;T~�Z�$9�������5�.ϫA���Nmz|����2$vQ�T�BЅ������x��\67Q:��rvy<���ո�5��:��'�� R]�mî��H	 �"�����!�)��?���~+(.^�5]+6$cL-$"\b@�C�\���B��ӌ�6��U�iM�gw��,��� ��l:b�#ņ����V��[�����W�	>�/�ۉ�]�.q7��mh,s*H�Z�|1u�,�� �'R�����E�F����r�H!���~J5��"Hs��A��?�q=��R�>NEG�����)Ɲ���p@�a%�!��(S!�S�l�9$.k��1��k�.��,�rp�o�!2ꐜB!18�<�E��4�,���y���ڜd_�B1��Ce�F9+K�m�:������Q
��j޾�2	�I��ڈ���F��ϥc�'�^e)瓽	r�a��%�ʷF�Xg7#D�C��w	�~��p�/e�fT��l3C��#Aφ�K��P��+�@�d�NvA�-�RJ�M_����PM#ʵ�iC����^�+������o�]K}�YsR+LV�d��x��5&r4���	�j�H��t��l���=�1�h-���A�J�鯜=u�>��N� s*V).|r�ۧ�C{��MU�*ysKb�de�����"�G��Q�)�YXa�q�PԨ��T��L�>��67�� 6U ])޸�������)��E��X���+�Æ��{�]��[�[T���x�����(�_���# �Y���sE�oG�Ybպ�0��I^
��P�`�����$9F��J�l�ƻGƍT&zcb�Ov��aT;����`�GW�b@���&s��&��&'�s��j`]������(NN�_���,�@�g�3������m�[ �������(g9i��!�rϏJ�!I�+8i��gDR�ꌏ�ѥ��]�%�y�l*��}Ń���{zZ�����0�K���$�QP�f�c�χ:P;�'��.��׭�:9��jG���� v�F����f�d,0�ĉ��ܢ`��3yu��ZZo�ڟG�}[�Zm�l%��Ir�t﹄X���A� @_<k�3��O?A�,N\��AC��<��іj�8��?/,�0���[q�����2ܡ�P>�DHi�>3(������6T4_QT9�i�IM,·�fix�1��Ċ�
!���ƕb��z�`��&ԙ����;@��q�5}A�Ǫ�"e���1��\ft�1M6� .�ǉ�w�N�'��)�v��G��_u�io�?�y�	Mm�D�xzM�C����Y�M��yE�#Z�!=�WX���L'b( Ti������^,M�N�GA�b��2���Sy��N1���Gxȼ��܁�ޭR|����X����ယ�;�(��V�JՔ� v���%y^��&�rط���^}q&Jq�I>��X&t�K_~"|w��PHn�㦫��g��c���H}�)��ٝ�� t���4���	ar]OH�0:@DT1�Qx/����>���S�G��=U�<�1�m�/�ۗ��_�Ո�C��<֍�K��a� |��2|�5#|JKn�Da���hx���'j��A�A9�tg�-��bŀ8�8'dH�e����͛V��4��E�	���Y�'���w�3�X�~��V�w�v�� ���KSϫJ_�M�_lH����g�:+fm��2��g|����uC8����^�7�e���ryQk'H�Nد���P(�1�(֍!�)��Мe��]@O����HF3ÜZcOÏǻ�kB|��� ���U~��*��q��%3��`��/�c��
��k=j?� ���c2�4��j��2�u����Gcf�}Q�^v�~���ݞ70�;o"��)�,달�ο<��'d};h��֋=�a����47�$R9]�y���a/�����ctM����5�{�h�l��W��Ej�DX^�:H� �֎N�|χi�K�އ����1�(�M>�|D���=%�
6�iE�Y��~�#��O8���x���4\3ї��X�b	�̮x}g�C]�r�%pl�1V;�7�m��ٶ���C�(x��PG�7�;�`�L*�\�29�]�}��&(d؂�[�'�hpѵ��[1i����
 ;��/47#��9�9�����2d�����w��m�ir��6�}�xgg�VOc(�p�s���hZ�:�]oG`�|�յ���Jĥ�˒��#�C5�P���`�d�e' ��$�
������߮7f����S83��`���V�e��oL+P�,��.l�Q\�5�$�(D�F١��2�(��7�'�;����%�7��`�C\V�Fjb����J���L�n�$���qi����(����3���l񕑓�=WD�<���90O
sܟh��|�cr�7����<�S䚢�1�C�H���	|A��J��h��%JfGs�P��U	�;�JY����Q�����d:@1�'��;q�-���+��xo;9�5�G�/ه.Pѧ��@ihB��#��_]���}㴿���K,�]� cn��iп�/��O&��
�;-����,���Ĩ�"�)ڂ��Ƅ�3�x���[�9��_�ڄk�j�`�����iC�'���!��)͚�K��N�ق�U�޵�Y�Um_�������IS��C�E�֜�M�x�!�%� ����K���Sp�K��W�A�	�'yo�X����M&}��]�N'Y�܁72��X��1��-��K�EBi����h��Y��r-����'��8?��l��w�m�3Yrһ��kMF��h��h�����g~��j��Ҵ.\-~	]�������A#�{>Er�<��g����%O��\�?��"Ax5>f�`���M��u�+���gǃ�0ݲn
�xn���uЂu��X�l�,f�s��d^��D�;�.gX�[���!�4Al���]�#����Z���'Ι���~h��_�Md��GϧZ�������Qn{ ����"~ê`�p�ԗ��g��3� ��ū3^�B2W��?�=����Sj���Րz���A�SEFA=�m�E����� ������3݆r��&�s#w8�܃G���w*8w��G�'^w#"|�>�����Z�K��W�Y�-�-<�!�MU�A*P)����%�m�����O�&�H��M	�Ѣ�m�����>�v�x�Z�%��q&��2�s?v�i�t}h��0�$���x���������)�ß���F�y|�!E�1�%�7�)�t�X�����Quq����j�O+��!���"b9w��DM<f���µ�q���m�3�hT����g�e���,.DA8#���s�N���}�[�K�[;RY�7�F�uHL�4�i�\�Fk�֛G���	-��
�G:y��lw"��$������ ~���%	C���^c+�`T>+�D
��xz�Ƹ��(M�e�e���+C(�VO�0; ���I��>%"Jy_�Ɗ1��w` ��W�����d�v�/��Ҷv 96�E�F��*�E�կ�\�)a��9~A;�.t�<T��f�p��dȐj'y�vk�EX�玱�[���n@�_6�d_0�`�k��U_h!��9�Ba�~[e8�=�g��G7�B��=����O�Ȫ�N���q$�	��v�/��}d���������4m���C|�S�/�Vսn�y>��q@�F�s����j����&�k���:Q4X=���B�!���֕�)�������F��{�b��$B�g}C��(���t$���i�aV�A�[s�&�90f�̍�7�Q*q �Q����?l��ZoF�S�J���rH�Ö^r���u!AC6�y�t�M�~��_�Y�-�uW���?��,S���8P��~�b����x�(/T�=��̪v� �����@���gR	�Ce5	�����l~(�����+��p�G��T�kmw�����ü���3��Q8 "}ݩd�*%!�r�/������Z�����g?�A�^�Ot�L��84��K�v�
�"9�c���9,��<���A�.�-��)�8��+��/l��D �Hy9�@�[��u������,�3Tמ5������qfs�̒*��v���~3�V')/@��q��Yg�g��\�c忏�	k#]H�� �+:y���	������21�bT��Y�F0�l��Ye�o��aj��d^,�c����,�"w\n�s���]U���%<�'x<9����V���L��7kcrQ���ƜM���Ԙk�Ѐ��4+��P,�����.�c�8��#0x��Cjn���'IآHH�
�C�R3'o��}ŧ�d(��L8�x^F$>��D࡜D� ��[�(p���?��}ŝ������� Yn�H{QR{��nP�Z����l���i�p���dƸ<�'�����Cɟߘw)��;M� ���{:��;C|E�����,��"�0Vn�3DMS���gj)�g���L���{j[�Hn�sA�h�;�SYwp�	l�R�h��M+E� �����N������7ů���3���s�s���?�IS31�ۛ K�K��4�Ń�%,�{��W��g�r셟��-'ue��vP���`8D�Q���J�r%�@_�68��#��=�*���ɍ[?�7&��/U���4t<��5��sc�tE��S��ma]}�M(�u��N��㟪������w[{�^�ՊT�D[�͂ƅ�p���R�Y����<�b18P�
	��p��=����[~y����{�ٟeR�sjCO�3�x<�4����1���#u.ӠO�=I��}R?���*{"p-Y��L#���������|D�|�����%I��7��h�)�zE��1IVz|3�ru�𺃩w�Q���G���t��8��[G�U��(��a��m�2�V�5;W�x���urU�!)7D�w�z4:qɀ��vK-&�mU	�K�W����)
	ᐂ�������n?E��/cND���V����jC���&z���[*5�Z����Q�zM�e��M)�9*a��Py�P	�[&��dǈ1��bHyK�'_+afy���vH�{���p��������UpdI��8���H�WQL�����)��ڑ��$�)!,��}t]~�s�ܕ�c��~�F\���J�Ձ\��%PG8K}���5����𬕻���coz���1~� ��,iZba;�։+���3u�w'h^�+lO1�ԅ��	��ٍ{�%�Ц�+�,N0Akh����'������=*0�C� ����� GJ�����j� i�˷����@D�l���/P���X�#�>��0���D~����(��|���
����n���a	�J�GBHw#ݛQ�B����u�j($���g�_5��=�r�����/`����ʈn�H-��΂7�Vx��G�o�W����S���L@;@/n.x�
d�etԓ��.��c��	G�~e����ޅ|�����X�%��T� �wH���qb}�v8�����`���u�N6*��K��|
0����EDoc�H��@鶣~�^GJG����#�X�
�,o(�t���7i�lp�}����=��*qM�G�?��Ͻ��>i)y��pk�FT8�/�x��\0����;�pR��}+�t�4ʊ��SGh��t_C�]L���H���X�@0+Z�]�#$(��<��@��jp��`L���u�8⁔��(P�	k_�+� _�/m$�[K��[������v���[܄Z]`�Z����R5�~j`�]���= l�ɑ���J{
[��]?֙{ׁ�"��y^��	x�w��x�$�Kȧ�m����I���b�</Jr���J�$�3cD��Y�+g՞��J�FN�b��.�W��X���66
�9�]��fs�AO��\���m�+�)4�{_i3�@So.�g��{�����=�ReX��A<,[.0�~�nO^�oˠ�|�����hN⿫��=�B��l�o��Ӑ���Qm�$#��1����>Dۮ=��9���nS.LB��iz�y�z���-0Z�O��+R�ܒ�R��#����?��TCo����I��|��;��I�a���bo��{!1C�<��A���)~�M�k�!�٨���y�si���g�T�(�w:��@7�2�p ~,�:��:M�P9�&�e>�?�˹�� ����
u9C?���6�麻"EDk���N�@��ٺx�c'�Ы^����î�FF`��`��g9�X:8���t�U��E0��$ T���	�?�v��FA
�.��=�T���+nh��st���w���ֆI�Sr���A|v�V��g5�D����M�@R�����/�P-�¾�]$�%Φ��K8L��@�J䤎1:iKY�̉�L�=V^$\�c�*C��G���]�
1)�o�l�Ac����+��V}�돣/��gD�o-���%�#�3��8z�a*��r��"�e�T��b(��u�P&D�˲�g39RC�C8�ߎ]���WW��k���%��'��^n`�@O^�Յ�t����lW���:��~�=Hc術����m�ײk�t�Ԁ���h�,��<d�L-N�(O��ϐ��9Q��q��%�4V�ڏ�0ypD/5�qf�(�Z�F�-�V��w��E7y�X�yO0�~4&�!�/{!V德�PPq�r��s91SY��u�`�J���O�MK3��@�+"h�a�^^�MWa	Km��ʖXr�)�v��:b��� �AN��q�fq�I��g�Y�������n�v�*���qY	E��cf7kٱ�I�*D�z)kߎ�0�@�*H҇���=�������Ɨ2�[�oUcl�}E�qN�2@R�~hs9��o��+�p]aо`�N���[6s��-��ź�C:W6�����E!=����p��s��uhd��b� _o\���놎 Wa~6�mݠ��voFqć߱��ՌV�E�k�i�.X�9k��q#=�W��+�xDX�L��A�#�B�#�p�I� �#U��s�}A�v�W�ݹf��T���j�Gb�HK}� 8����W���P�����a<��>�ؤ����7�p_{L�m��3L�E��v�g�ʁ�b
�ΆJ��^�ߧ��9�C�/����V%���=G����re 9�����v~Mg~˟���!:6x�,��c�y��1�1̛�(�_,�'�}C��(N���G,��%q��6U�Bz̾����Aw�$8]��f���K!�@���t)c�ة���&����>�O���_{^���گ.�&)
����N�c�c ҿ�*mF�}[�$����AL�m�>�uG���*<>��6?l�0nӴ�ɜD��Ǐ�o�
���Be�Q�w��� r{�4��S���`��0��^t4�������]�fI,@�P'gmM#�����=/�����ʔ�@��p���$��+=�� ��j�v��6��f����4��*�=M�x)x�C����=���]"�6�xZ�B��`}J��V<kvN2��cH�����R?,R�Z@���z����D��Q���QU���e ���9.rd�3Tq�;S~�H�߄h�G@����Q�-�(\�0�e� ����#c�;N��j������T���ײ��I���cM�0J��9�]�|�5#�x���Џ���\�[��E8N�ox�k!hF�#�M!8��	�Ľ߹�٬���P�_J�cEȞ��ĻB�uE������4����b���dM�X�~���Н�2AܣnuS?R
�x'6]���R�V^; �	��c�x����-�v�c���i��<b��7�4�e"G��c��n� ��x;�'�R���L�����c�Ƅ8)a��ΪA�=d�{6n?���>��wK���,Y�Ĭ������4n
X�L8Q)�A�^�c�N;��Q�&�4�k�՝;8�+q_-A:�b�{�7Z�i�����E�d�U����$d�N��#�"s*uN�I��hIN�e6�Vf�h�%�O
>��%�]0��"�f/��)��&To��TI�,u��jĠ֢*��Z2Gk�4�fA�h���&�B[�㓭٫i�j~�����+���\�&a�٩�͈1��I[e�ڔ�G�����VTNk��dɌ�V����D��$�J11?��:���`z	�/l�L�i|a���Yx+�7��d���P�V_ͩ`���4���:ț���f�y�v��ٙ&�Y��tf���7�gư��Ң�v?.��-��;h������lp��l�B��ǁɟ|^�G��[Y�������zL}!��3Fr:d���"�E�J+=�B,�K�����%�-���{N�m�����p-ί�"!�fߜ��|��"���i�sJ�B���*nҺ��;�$��)�dӋ7d�I�O�M���������
%������9��
�nq�=�&"��+.��_P�����K>�)��0ͷ������e�Po��,[�ԗb7�Q��US�~����C{�F��>�3��M�KU˹p������/���� 6�z����j�n8��Ӈ��qU��E��p@�sF�
n���$Gl�-�>3�����-|h��?�U;�c\�Yc��Apur4�Uz�uȾ���ԭ��&|�� ���IH��GB1 Yv*'6�&�>��֊��.�Ar�G�颲� �y��M�� p���D~�8j�c26g䲻^[�XX�91�\N��H�]��Qʏ�o|��ԭ��ج�ƒ&����4zĚ�Ni0ʘ��o)�f���y[�Ex `{9�c��S"�Տ��i�.^�<�Z,?�$bZ/	��z��(7+L�n�1(V�f�s,C����ؕzO��Y��f�Lu�xp�$~Y��'PP` �v9��Ĳ�:�Hzu�N��F���(��l��e��2UX�xZ�j���%���R�]�L�
��ޜ_��Y��_�Q�2Y��o�۬�S��mS�f����P�_�zV�e�(K,
�P���.�Π_Lp�ʹ��i�0ކq0�������P�F�ԗ�Zp5k�����a����Bg��hbH�ݛ�5z�a�2�Qg�ڡ���>�4y�aX�#~DDZɫt�q��6]���K;V��z�ԋ�/��U���͍gu <���[;f�?FѯI S��!mA^5���	�^V������6f�)�XY�7@�C�6vD堕Gs����1�t׋&G�B�WU~����+�J1G8j�GP\,���f�x��ՙ�ҍ`b��(�z��f���Dl|(��jm���{%T�ԉ�&�ߨ?�	bE�D��c�k�Y��Ί��oKJ;���5��ɥ0�����K�V��yo�S�Bd����r	�S\T򛹕lmܭ��gL��i+핯5U�!ר[ìkT�~�Q] ��B���Z��2�_筊�~�J"@��8����mJ����Z�����H0�j�1o@�Y8���8���p+ɯ��s�#2!%��'�`����11�Y��uU�>*r}o�$�uN����C�?�JL�C�L�W��)S�cϢ$��m��@d���h5 8��0��y�N&��=
M8A�$a�R����b�ڐ��R���T`;�;��d���~���51�9ʕ*xW��0k����ZcǁS�~�։m:��.Tg�E]�;'��O��;�P38�`�g
����E��0,:�雛n2���ֲ���nU���)�Q�gv�iM�g�����0FNe"�V}@kǸh��~J����E���==D�V�7��.��K��Ieg�ͻ���&ѕ����w�@5WP2�ʏ�^w�P�����Jᓔb�����[s{��X��2Y(��|`�r�ש=tm�T`�Cϐ>��@˙�R��)^�vb�Kk��AF�U7cG�i���9.�������kL��,V��>��oF_��䖈�������6S�ronkђ�T��ݣ�V��W���SWEȷH�D��R��}s����CW�라�֝Q>1#����]1�cϫ�>t6d`�p2�0���^�����=[��0�
��4��ت�׻�j�<��S5AD!��\���i�m
�-]����>&��Y~(��Hr�z�B�n�&��δ�3-,��i,3�,��H(ѕ�3��}.����%��c���V�1�)� �S�g1����~�g��D���h!'~Z�j�t�]K���?�Rw�	|#O���2¬��p$P�g��u�s�M5"c���Dy3��h�8��T�Il�d�]f�u�	M�^�΄&��n���]���uMt�S� ��iV��l0ia�-3K�����*�{�P�'��s�&� �Qq�v$V��d�J�m�������x���Ge����P@3�|GB����%��Ƞ��a��K3frl�J��0ms��M��L,r�!� g�ړpucAGb�4�SH�,��¶L=S�*���,��Gr�?G7���:C���z�l��8�&���j:o@bŐx&'O0�Z��֧l�?,`����]p��l,�$���^ap�t��e#���U�����XP� O!5�?���74M�+�&/�`�6j�K$��p����\x����rվ+�h��'����IF����t�ZD�=��z�&��fk���p�YH@7Q1.��$�`ud�LYjW��/� �����<�k��h�x���/ۀCyF?Q���/cV��X�BH^��+y��'jȌ��A� ��=v�!/�,�h��$8��R��dvCl�g ��/c�s��"֨������K�	��E���|^���/s��J4#���=����@D?����b��#�&�A�^�ŔQ@e����N���61�g�>Ea�߉Y�tE�[�e��;�&SM�}!f^ =�g!��Z���O�x�٨A7FV�����n���Rwj՟�<6�w@�G'Mf���h�����؝>��_�&�^��mʶ���'�TQ^��sT%��G����\ ��}	�@��4fao��B�ӜC�SNN�l�[Υ�T�!���~�����$�Xu�Lj��ԣ�֦�?l�:�$�����5��4Qm��U�)ɬ�KE�p��/e��%��wӆ ���w�M�Jf�˛�. $��Ʈ� �b�IIN�T��/e �k�ށ�F�¶�PM%Υ�j�[��JN]��S����4�g����dl5)P�H
���;��^�ЗUC���lD�����#F�Qb�[�A�cv�I0q��u��j`Qnң�hT	��}e���˜��R5�@ Ϭ٦SQE1N��1����]d�m̩PkD�!aH�$l�������^5��%I�O�\iX��9�GT���
ta�F}�z�$����W�=C>���`�[�Ȅ��1�j���~P5�_�ޱ�E�e��e#��I$Y7R��\�:
\���m��+{�� C��,�U�3�{��9<P�H�n���C*Y<�M�g��K.J��ҷ�.�2���$��dq��Esb�D8Hu{�kbF-�H9b�R�<����32��p<�]*�s!Z� �GB>�-�1s���>�IO������Zbd���4019��	[2�Y9��<�n2�g��l�B�te#9��.Cyat���J�0� ডs�qdظ�)5o��I�v?Q��7��*��cz�s$U@�R�������^o����E��й�cB@J�?�ԮO�Y��a;�t��A��)���^��)L�u��(>{��N.-y��>0]
O�g?�5�����|�o�c@kΐ�3��jl��:7�N��XSMSlW�cI8���U�;)#j82����Jj#2r7%_�"jQ����Bv咂!\�E��5�ID�%%s��k'`�xS �T��(N_Pє���5�*���y�0�qm>*�E�8���U�F��~}j�����J���q�)r�]����؟B�P^�~�d��
�"�� �l�dlp�My/���.H��*�W���\��U�25,���l��C,��mA�@�l��6$ �^��Ψ�N �!�<�4�û�_�k��N�+Iv�bNP�W��Q�6,��M��4���́�
 �sx)
��F�\/�/
�|,��O�S4��� �+�˲S���,�`�C���a����_vml�gY���4�0��#�W�e�ǄR�)�g���<���:ٌb�������╨N��6Ɠ�
D��)TuPz51p�b�YK��)9��\�Kb��{���":]OoDqH�U�r���{,���]��?�#݃���6���t*AU�J��+P�^:_�B��Ơ{��7�)+����Vg.����+:��Dn�z)�iBN�/�d��W�@i��O�m0Ad�����"����J�5�S���K! �gBf,0&��-�}�C��7��Q��
�ay��������}�v�8�2�}~�0�9�Fdk�O�O�"؊P���e�����`��u�D5�d��\�ʿ���b�m��� �z_�%Ie�(ϟHQ����w��8F�srψ�I��"�4��y��l��2g>e�:�!�~�������%п[,�L���:�%��{�C�>J�|&�L���wv��i9�hc�wj5�}O�/��ԯ���0ЙW�9�3 G㫔bz�+��KI�okX�4��u_������a���ƨ-���"��Ԥ��##W�)��+�q�捙�?4���v�+�v�eFAh�A���Aö�9��� cw��]Ѝ��U��š6� �9�:�S�B.��t�c��3%1�h�3w�Ʀ� !�g��|F�p\�[=�nݟ|W6I�89'�k����R�LT����a��<�Z/LPeJy}���L)�D�E[WB?[S�d7l%�(�rҘµ<��+���,���>�X�\3�2]����p^����^��^Q�}J��#)���8Ό�>_Γp�8}�]������繬�J��2l!��~�"��k"C��,}0Ǆ�P,K��z��y�S�+	hs�H�����	����ΰ���P������$�pxä|� ���7;e�jAo�3YZh�� �ܺ�j�=fɋ�%����>�Y�[Ϝ;d���g���#K�	�9�cS�SuԎ9�i�E�#� �RR�&�st�	�.l�:�9�xǈ����D���csr��jd����l�q]9��O�9�t��k��qO������pd���1�SMR�C U��+D 0��a���`�Ë��YL���ҧ,9��d#�,�cX���\c�1FW(��E)�M^"�0��Vg�]��S.$��snK�� ?�`�MF�khBzS��[63s&�3|���;��
�8��+�ص���(�1�1�����Ň����	%�ʲ����R���v�W-&e�1�aF���c���2^���Y1�U�~���첟Sn�[}�i�I�<�mA���B�(��3#AV��y�ˀk����S�i���\L���4'�jE�Z�d�����QkeE�>�� �iR0�Ah^���+��B����F�,�(��-5�w
#�\:hcs�\f�W఍�͞��N#rd\���Z��PEa� -dӺ�j����[�X��/>�G'�s���tܵ����@�4+xQX�c����x�8�}�Nċ?�Ũ�#.��0�)� �P�%�����o�B��}�M�hU��o���Rzས���)�9H��~wC=5���?O[=-�H�nX�Ѯ�ɱ(O'�z�و��FY��g����
]ID����=r�Y:vB��Ef��"�mWI�ꞿ<ߜ�3�q��㦻�d�׸&�/hN�ɴ��E踴 ��.\�ϔ�V��ܟ���d@����!�bV��4>�^������6�^�b���ay����bbϠ��">�dO�f��78�K.��yﱐ��DZ��K��S������E��$%�ے��$5?\M*�Kga3�g��k��e۶m8�bDW�,LyN1�/́Z8�/��Fbꂑ�}Z;�������_����BˀŁ������2_:쿭��6��D�^�,��;�.�4rYG�k��fLM
B|�)�n)�wm?���va2�ɽ��T����6���;Ai���۱'qڻ��} �������Q�i�=\q��ò'�_$����_mg���^=�v"����)p����;����ܥ�̖��1P����B�]&7�<f�h����G:PN����1�2,*hM�
�l@\���XA��Kgs��sg�gñUY��렳���U#г��ZG�R�b�Zǝ�LwQ(��D���xh.��||9�����Hì�/)�{���&N�!�6��'�X<�FGTи��m�bv���Gm�{���5��65�F�J������-z�,U/���c=d3+d�o{��Z��Sd���D�(C5'�g�cm&7i���X��U
�J��A��6�elP/v��2��'_q-l;�Ğ���L�&�䙫~�cv��g���� H,&���nG�ܜ�ب[�6�>V>~��Ӡ�&qX��E���i�m��L��x����T9)��?P�;w}#��'�]�q��l�����G~u���+i�n�4�A�}]L��p!?6YƱ3�����Q��~ET68�S�7�,�~o%�06-*�rF��8�f�o��c��p������^D�;���2|��L�u3-kF��*��D��]W1<�j�/�vĥ��-)/���'�̉�ͭ�F�ǽ���G�'�tbf��?SyP��kFV8U�:ny���gyk,�۶���~���������?�Z�]G�+]:l�U���vt����ڣ?;n5E)�U���:��d]���������tN�Pɩ�t�SP�2Ll���:�T��s	���H��7�y>�S�Ɉ"�x!�p�i� �"%��0o��k�"�egdl[�9V��e�/�H&�h�.�È�G��U��r,C��t �&��2U!����6́<>k����䫏��N�a(�t�U&tr�pn���2Gp�����JR���6 H�y%MJ����l�{��xp�_ o��h(�Q����,��������'-�@]0%�	1f/���Z��ѣ������?�ͧ��	,�P���:�p����Sl�������Rb`�#9�:b �8ar nuD�+��{���.�G��6)S
���G��<��h!FW�^~�~-˲ 6�$XEԖKΈ�s^q�]� m^�Cz�l�sl!CP�b�c.�aE����Q�e/z%V���Z�+f]G�b%Y�D�]+\���D�	Ԕ��&��UG��?��>��d���KKK���m"�$+��[r�J�S�Ʌ��@jl�+"A:��q�׭�s����Th���x�r/�h��4� ��R�=��c�Fk��>Z��&�;�	�# M���Qy5��ŎԖR�؎�M
�E� *���S�zI���* ��M�H��%�8�#���kR+�[t�RY�V�=�f+�<�]�x�	��e����(.L�q[���2��4�/�k�XE/�g�K�O-��i�+��*��P�?����&_4�P�[�6`�H6�U�Q��'�M�{��O����¹�dw'�?���Ib�D��&>7Z���HL�<�L�ѿ����ޠ�\>�=+>����$5�Eb��%�.u�2���=����[�̈�Wٕ�r.f���:�}s�����iZ�D{E|܏��y���'������/��)be=}��2�$K�S6��!�ֲ[(hn6 T�%4'��������m�xG�]�(&|H>iw�������N��n��w����h���u�{`��0�Ϊ�i]��o���6��U���;(N�������!�Gr%��4������Aww�`bP���b����t-
8^�L"u����8�R¥�x	�DIX��Ś�׏1p�g}�����G�)�#K�װf�è��g�;�Ϲ<^�����\��I�-��������"���Q�Wڅ�X}0�����E��|G�lwM�7S�׉��%��+s[�k�3��K�ܛ������gV����{���6i�]��u�`��[��ͪ+p}�{������+�<���5�|��3G.hk$�ҥ��&�<�C5�i� �}(��4�O���zG>������oB:أ�o�$���pseH^<NI��ն��R�stWݲ�I�yP�d 펙-��f^�����x��( �$�nXk�t�O��5��Y��4�}a�1��!5��;���~⭒QezT�񱡆��h�+2�Mi9Z�Lp	��Y��܂���jv:X=&����%��b��x}�l�O}����������&�ll��C�����PPm�v�hnaN�L$s��]G%� Ϲ@���F�E�/��W
�y���C�;�0��H�,ƌ�,�֩3B(�JW�p��oe��Vic!�"��<ȵ�h�[��,�;p�q{2O��j÷k�P��1��
֥]}��U��� O�h#�&v.�r��fz_��U8��1�{Kg��T1����8�l�y�����̬�V=U���qb�<D�z&X�@��cMv�|s��0c����O���@���qLg4�AZ���LY��0q�QrQ�k�l���^a~��RTBo��y��ǂ������w|�OU74�k�/�l[q��*����O-�*�2>W�)n�[�o�1��<���~�	��A�)�i�4)��\�?1���秓HdK,�j4��˽��7�D��cRE�dD ��vģ���U��W�-��1J�6�f B9_��ɤ�vȅӲ'%21�{ns�YE��Y���:��>{�$ڷ�O��M���ʮ?eM�ՠ�R�g�Y�/�/co�*�������h�ze,Ǒ3�hI��3}�}�b>��6VK��Y�G{&`=뷧:](� S�������k���@Z(��-3�8Ȅ�\qc�\�]�@�-6�mݹ��;�d�<�A(/��C/|
9нI�F�Ԇ�a�̚�b�#m̺�;�v(���~�+O2���7Ba{jK܌ Ȅ���b�Γ�qk�û��̉>�Sq���E�ԓ\ �ј��߭\��O0�VDɪ6�p��:��mlȿ�
@8�����m ܼ���J0�V�V�I�m�i�r'��!xU ;�+�58��-�M��J����:�ش"=M1{"h�f�`�ܿqV�'���%�x���T1֫?末V���.�Tn��R�>�wEggu����=3��F��·������=�P=��2�,h=��I`����BÑ;*�0q32�-���c�Z�į��#۽�K���Y�������+&l����b>6:�-hv�pݾwE�l_�����f�o�A�v�ĤN�ʻin���/�{��AI��|#�S��0詟�e�]XʋN��E3�_QkLx^�(V1�8���,��ѲE���-���Yj)��SK*����Z&݉��s@��K�t����qCx��i2k�� Lv$��p`�09�f�����3��P��N���k���Z`� ٱk�]U��N|�l��?.�h$�2{�%�~	��U@�-d����@!g��/�^)��(���uؼ� 4ʛQ�W �Ķ���I�O2l[D`�h�o��ף����%�?ĵ?Ҕ쏧y7dn$��s�4�J���C��[��?��e��d�n��EQ.8���c�Ѿ��؁��=�J�3I�����zP�g[т�i�{т�U����x�uS�C�A��w�v��c��H��FE�z.eT9�$��P����uZ�Gr�K�Az�B�d�A	�J�jAl_|�(��OWF�c"��!b���� w��h�oL�����5<��>-� �bF�_�
3��{�Z+�`�%XRu5I0%vB����^� �Q��>l�m���p��E��m�̈́���%\KҴ=>H�^vJp�Ծ��0�}�R$���8G,u���,���B��o��_�5oP�o9L��O���Q��R�-3�К��r�n÷
���T�gB�J�Ӯ��KL�e�����r1�Ţ�D�ٺM�>���k�z���3�|/�RA���z���̘L���,Lx� c*c�Ov��3WF�V��ФT��R�<i����Y��-���	Ŋh"��B��6FX1<��}�Ki�^���%��N@Ǟ٭zX��iQ����˓О�0�
���g���:M��~��|����.L�	Xz�m
D�	���c��:�1޷��|75�A�2��������9_*y੍s��i"x�Ƃ[��,
3d�U-��#�&�� E�������a�yyyN	=q��}��&�sw}!H�<i�v&��?mւ��u���5r����O܅.A�@���Xg���M7�`���CRru��˴J�JS 袘���2��	jZF̀�4�ˋHIz��-m�"��n�k�c%B<_z����	�mߒN �5C�V�O�dZ�ӗC��
,�j����2o�ך�v8�LQG�ug�V��9�Mr�_�˷�'o60�(�]S+�m��N�k�~�ڧ��=�[���Z�ۀ)Y	���\�]��Qd�,#�ALS���V��&��({=�&�����moQ�H�YU���(7<G#m��L	�4čx�y1�P�����'e��!H��9p�,����η��`=`8Y�\�1���<b$��pk>op��^���g�$�HV#��Nb[����s��l&��� �C\��u�\�-o�?ۗ�v�9�y8�89�o����%eЀ=SRt���z���;i:���d|�4hA���'���]m�(Gp�h���?�#tP����6�d�W�ԡF�_Z���k6Q�)sa���+꧴�A�D�&[i���D��q�.U�S�U�]�&��ω�70����ɬ�ѩ�z�oFAq jh5Ԕ��v}{)�W��\�\u�J��v�l��R1�Q鲼�n��n�B�m��4�ß�: ]v�7?[~gQ�#�x�W�f�f	Id�8�($p+@Ԭ���,��n2_��ˑaA}�f�Sh7��n��M.)�|��̷bf�c�E.��L׍�v��������	V��_�q+������?�k��a���K�Lӂ��� �A�����wc�2*���d�վXQ�J��6Tš?;�����uRj; }�7�� ~�{{�l<~�&#��xT���%a 5J�!c��@����+xr�r���B\�I�ٴf=1i��
 ���}��江 �R��%Dp���zZ�J��&����~~��ҵ4�."�Z���]j���qk8`N��vmU&9�b�s^��9b�[T�H�$Z��� �X�U%�l'�[���z�>����gS�4�E�g߃���cm����J�&�w"#B�݂��Pտ�QT5��o�m!O769B�[�<��7ڕ�Vu�g3�%��[�1�^Uम`�~Ma�K�`8�XJ�v2Z�$T��s%n\��$� �	1�����Q�����p���Q������	�]�`#1ha�k��nlZ6�,����ñ�R(CT~�_�% ���1��#��?��荆n�g+��j)G��/_؏ơ޲ek�����"��h�bu���!���S���8�ܠ'DW�\ޑ-N?qJ�rߩC�X�h)#m�H�!x9fI��4D���������	��W0(Jp��� l���ذ}/k�k��Z[0���P���J�]�7}��b�(U~Vd]�|��AvJ�e/�v��?�$�����q��22�K����%vd@��>F[��]r����>*��-�ʧÈ���	l���|e����0���t���zo�{Mb*�t�`�*ƅ��"���%�Y-��y�Q�� @\�6��F�B΢���L�~a:* s�j�sORG��!�p�-�+;ԤZg��h9ږ]K�ൢ��S6�rrsq����+W����Pv�,�)�'C��L�9|;A��=�d���yy�l��"�E�P�ֈ	�6����L��LRՉͬ2�����{�w���o��obl*����zJ����O���Şx���Zs4��0oX�FH�Zu��^��g;-���E��3t�V�N��f�,����cy6|��tk��40k%�:p���>���|���T�.�.`+���Lo�.�Q�����*��yJ��	?���H��#>I&)�F��˽��̯�A�gԱ���� 22q6��2K��!�W���hzĎ������gTz�v OeЍ��i+__�3�GB ��2��(3�@3��0�3�)�}�=��J��U�7���hO��ȈK�cg�4�j%���x�FFrR	x�oGw��13�y'�D]�E�D�5���[���UMb����q�&yڵš2������9P���������=���+l��X�6R�8�7¸�^�^���-�hez	,U�9T^�Sr�F��!.�����r�$�a�ѪN�W�qC[��9�f����t��{N�Xn�m��1D�2z٣$������͠)���S��ӂ\��V���K�p��h\!�G` �::Y2�=��v\�i��5:����+N�K��p�'�)a�1�X��^EA(+A�C��-�3'����ж)j��#|&r OH�f�oC��H�2G:|q��������7���N2����QThV�W����<������},��̲\��r�G���:4�ۨ��9
�R�#:���੫���CJ4x8���>W���,'y~�N��g�E�3�*eo[E�ڻ��&4�Ww`_���v�*`�$&2�=	���}���n0w7sx6�6�3.א�L��%�V����m`N`tWc��?�d�;k]C������)4�$��Dp�0r��ȜXlR�1%_�ލk4Tu����� _� 3���,T$�d�U����s%���e~�*{G]�!ԓ5L
��|r}����,��{��Y�
���1���W�z��ЦN�~��u����L����쫊π��?G�{��F�Q��T�6�/f����Lǳ^����ߍz�G����*V��������X��SG��D�=��OB�T��9[�\O���jU�lJ+-^��5u޹f�}����n-���r,-A��/+��^�X�s�t����P��]d���]��y���ZP�z�fk39w�}������>U�M�R`I��~D� ��j�
�I�^|T�A����A�u<�؇�
P���
Ѽp����ހ�U���s���	k���d���ϥ�y��Kߒ��*L\@�z	_l�^���'u�8`���h�	��J3���<���\V�%_�_��w�AG�۴���������9t(���ԨE��jKʥ�;Eua������C�p��Y�����ɳ�� �-�i	�e�||��s2f7H�yӬ7b��|���4# q^�����V?ݜ�w�5�h?X��̺;/�8��R�	�M����	2���/*.�wc0Tz^v��x+a8�
�
2K�Y��("6�"���d����&p� �(l�#������\%�Շ�4'3���%G�˨��:��6r��.�!�],��j��:*�x]X�X�)I3��h/��`�/n��;�e<>\`���}��7�N/�B:��z[��c�on��zup`�f��^��=�y�N�Ц�M!t^���rق<��$Iգw_#��/�Jv��݋��Z���/�SR`m۫�e5�/c�Ί���m��
HB�e�>m�E��i�_��ͨ�A���fk���b�!�r������gM��9;�Џ��Դ����ԧ��T(�Ź��|B_���T�Pm��R��/��;�"j�G�\
�;�V�^���6�<i�Gt�@�G˄��ưk��V*ʄV�T0�ځ(�X��|�x��QɆ�k��H��-��!h#L�[$�M�6*!םX�g4��N��4Z#̉�Y��nR��wg�:�eE��V>��)
P�u)�y��ϟ�!��A��2�98�3|ު�JH�#���Ϩ|�敟�+XB�P����J(J����e��3�1��+�"���՟n�Wy�&MM����c��j������]X<�o�*bs��mg�B�.��ݟ"c����Cz�՛�A��s@���'s���'\0G��2*�Jey�9;�(Û^#
'/�ҒG�i.l?�l�홟vƛm6x�(�q��p���n2Sg��n��ʍ�wl\B��$?8F�>6{���qJ]\���w���8��I�$�=u���V��~IY�g_�L�����$cP�c��D��x���K/�["���X�k	��H��x���3�z�Y�Y�ƾ�#��Gh[�5|�*��݋�c؜�����QL8��Ћ&u�vV���W�c��Tړ� ��Ȼ��.�Fw�c���m��-�˅�J��l���)��-ت^ik��^���d}cgӺwp���O"��D�5Y�����7F�[J{Mڿ����0f ��c7��&����,�+�rw=�>��V����"52��_]n�FD���]�����e�P�@�\j�٦c�d=`[�*U ۲�2�T?�hf�j��gM��
ۛ>(*��u�?]=�v]�|��w�5�qTu���_���*��~R#�)��j�}�7���oGoB�~���?�]��˓;�9��t�e8���M�Y�7[�%��XjleRHt�ga�m��gH���^�FS�?߰������۫������	�������?Nu�Z&��sҕ)s�}�8����V�ߨ!���W��X��ou��[��c�ߜ�e`u.FِP���ё������yW4^��;�9@�!����4:fB�JtKѼrҎ�*:e�����##6;��w Y�]��V�'^�}�@kH�ٯCX� \�4JH㩆��v-xP��0��*#)&vşi�ٖp7�7ϑ����Q���+rQ�6��{��ykr��!��K�J}�-X�vTU}���Y0'��g��F��=���M�X~�����w&`XGI4��~�M�{��cpDK�Feu,*Ø�p���"�<0a���W3s��<8�>ͣ�����)��mLò��z�ހ*�S��^Q<�yQ�$��C���y��[.+]��{bL��ɯ�x(Aa����1t&�rI��L�yڢxX����8��'�yg�����fv,;/꘩ƈJ˶�PJ�E.T�1��I���N�k,�c"J�va�T��u�"X�A���^�^��Nxl��U�L.2�:���6�o�8�1"O��)��Qd%f}��,���yՒ�u��A����$^5��ZkfR!��a�Ǉj�R�=t�^~7�t��K(L�&8��w�"܇�,�?7ϪQV�5���g��}E��ԊYI�)��Ppl5��6:L�~�!nۧz�i�Y�
�^Ixr
����J��o��L�"�6M�:"�=bV�Wz�����[�\�'X�6��g�43q�}�ayJfs���I�HR8�>8$�EF�v��X���b�`��������b���ӽ�	z��8i�U����J+Ǹ$ס�h\L��Eq&i�;=�W�W�ٳ+�=f�L�I�	��_��O*� ���v�}/�&L�D+�����g�f���F��uvС�2!��#�9m���,�eV�ϻ�9�?�D���,?P����?�d���*�!%�G}4�x��L��N�~��ȍ��u:��ء)��; �(.� �;:�.U�!�i�臝H���͂u|mK�6
^(4X:gga�z&s����t�F���
@���ȓ�w-1:�qp��)\����4)b���>�߾����T���g�N����Z~�����'#{�D���cjn�h���1cfpJ_�>���Id�����@�ӟe�.�۫BY�y��>��8�)�g�G褽*X��)�H��8�z���"l�/(��ፑ�V,=~%�Ʃx@R�9E��v�B���nb��G9�]�5Ƒ��1U`h��@Y�
'жm���|W7��ꤶ��7�G��<}��z�%�"%��N�C�$�q~"����$��(�gJ�L���3��!��2Q��/u�D�gWi-�uv�1������w)��R�NK���ȃ�<��k�r�$Z����BE�I\�m�^�YB��S'�ui�p?q�ֳ����2�*�2�p�̱�!,$�U7�N/^4n#��¾("=��Ű-	U���l��rM�y���SM!����y8ש���=kV���pp��R�cr�`���'=+��&+&yE��"���"
�!��!RI:ŭ$- �H(���	�O���9]T��ì"�J���'̔�����kiZ-�V�D�4��AZ��x����=��
f��F����#q�j������#�c}���k��a�8���Z��|��(bi�#��[�(��qT��Zo�v�HF������Wr�i�骘�y��h�R� 40¤�ժ�L���]�濝�珝j���e�2�J��d_�������@��ll�CKo'�F � ����!J�|S��*��ĩ�F%�q���ԏ�x�hBGbg�pP���}�u�* ����cAԡT�O}-�^��G��3�d�\��������
��H4�ڳF0�]+��ܶ��o�%��Dl"������ ��Pd�v������0&Wv��KP"�/�Wd����Z���H�pv ߎ.�SIyy~͊�Щb�Ӕ���̶�V����+%���$��l���Bo�/�< ���V����-�fbfbڝJ�[l1;�P-d���!2�"�ĝ����ߤm<q���	�xL�&&�#��ل���S�*ӲB/r�m2m��n��ZM�8�P�:(b����-K�PW��A[>��#���vm�4�?}ڳ���N�8&�+I^��8q���9����D���7Ct�,)����'N����ͭ�x��E�kƟD_7��6g�L;�%�R�mi��@m�E�^go��/O"���q��,*�{�i��:^ӿ�F�W$>��X:��s�\#��ʬ�s(��|�����2����,|�jD@�r���9ř��	�u��3s���^�uOcݪ��:Ψ|4se����f�\���c�G�W~qz�֢ըϾQ�I@��JZPt��-��;�w��ق��	.��v�������f9��B#���7V���ؾM@aZ���9���m+K��,����a��S�(�Xh�1���O�yT'�|X������S����f=�I��}`�������$sw~�gqH#�]�7ES�?lZF�'��y��"O��vg`��5�X��h�S &.Y+��8dMm�|�Ī	%l�@.o���(&խ��L�ܬ��x���L�&T�Wk7��D�y�=�5��%qr�NGl���"6	�6�ڡ.�����f���y2�Ik��v@�DV�}�l�f�~��X/P�3Z�RݘPá0}��S� F���bTFaP�\2���퓂JB���E���%�d,�.9U�Sv`3;i�犲{/�7Ʉ^1�:��OZ<���DG4R^���qo�����qN�N�Γ]�`�m44�!�5�o�E(�	S!n����:k��ϬL���fj�V��q��]�u��L/,t�8��Zr��3뒤�M�g�΃��rO���?Ӷ�s�90�d�1Z��g��`C����yHR���[�ө�{���ռ`�A�q��p�u���x�8�l~�t��yi�ttพx\��kB8��0)d4�QA:SUtB������&@|���tpc�e���Lמc�C�;G��7*!t;�"�ho�僳��[�������ܼi��]��A����/@ѧl&L}u�Ng�y�\2GK&Oj>o#x�hЉڝ>sl��R���J�,}�Z�~z�[Tz�0e��G�'�g�~;� 7fH��..��9Xr��iv��U%Ŭ�ʧ`�i�,��=��o�12w��!H9nq>�u/��L��~���b�?���O�(G6u��S3g���-^2���<�ڥM!�6%�m.炍u�/&�a+��&��p�C�t�	��Y��N�CtT�}X�t@�/����ŭnoڮz�k$����RpM�������tәr
'\N�{�򌹔�#�}��T2�΍H��~�u��T��=�W����|��\|j�W3��U��sc|M�H�]Xn�H�b�d��V��oH��#�����U`�F):nL�9|���An�DKR��|����N�%#�?���'�e���������S}���=�'bfV���5�L<ix/7�&�}�����&5k7���[����[ݗ��%�*q�:���I1�܏,��'\p��h�-dA����+w��ۗ�>�b�t�@�/��A+H�-1
�wS��|�}�@���zY3��\�ٜA��/�Z������.��"܆z��K�����
̳�`Z�~�\J�`�7����[�P}��ׯ�تL�n��~A�a�»%��e+Hώ@��Y�����ze�}؛�nܨ7+4�e/����QE�q���^`��o���7�}�)6i�C��`Pe?����j;��}vf���^;���r����z�^r���n�Vp}܌���6
���H��â?����q�t��ӂVb�4��b�B~r�(����ߺ��?O�(�MH�S,�z�s"�{7�ͱ�bf3���P�C)疣Ԙt���l�־JO��o��#�ڛ���-�w?���a	<�uX0��J�*��˶Xʁ͐J>p�_�c6�c����>GJ�F����R����*C�V2���x�����U'�̽5i(~���3ԃ2I��!r�3!���P�.�Eo�SBd������0��]�v�������F'�S�it?��E?�)�#
�0p���'�ܒ�/m��zM��P�uS�\��
�}u�I�	�`���,�.c�俓˿�eܬ��ԗ�j�:hQ��C<7Q������}�d L�q@J��,)�ӄɟ�8;PV�H�u^�/�~��
����W�nƈ�l��&��3����7LHq㦳#�[:�m��c��1:�l��eK�x�mh�Cm^o�J"��x�T,�V@?�Y�?�N���G�QJ�zrw�MD�Y��G"��;߼s_��W�~nJ=���^���y���y� zٛ��x�e��?ȓڌ�<.�2��B[�v���He��)>�zЫ5�^���5ܧ>V�����F(x�	ma��L��X/xP�=�F=Ee�`�\�(��D�nsH2R��#���C�������ې^%	6�M��X�֠���/��B�8/�PLw�Gm���$�j5�qF�:Ά����K�c�Sd.��W�&��|:�X=K��U�2�AΉ��55�^�9V���fI��kHr,����E}�%za���Z�A��4�Z�&����j������Pҕ��g-���
ܷ)8a&c��:�܎R�tK����������*.�Zﰩ=P�.�pß��P�qo�"�# EU[).ȱ4�����<��������1��PZ)��_���y�W�?nUŃ�o��m}D�6	U��?7�ęH��d	�O����������P������"r�bX�Z=g
�*p��K��n���C����bЎ.��wY����C��!#�&`��Y+�vEݘ'E�ˁU�Z���pnMj�Q�����O_���<��0��>��0ыZ��\��/m�L�6��Ԁ�ե�!n����?����zA΀�+J�n����ƽ�6:ai����K��|�T����5�W��Eę �	}S�K`���ŕ�s�`�w�(����/��#&�w꠭�T��ۙ#�x]�c'�,�a0�>�Q�Ǆ6�O�� v �cT8c`�л���(��b� ��Z��eC0?�ҋ渇z���p�u��K�� �/Tf���H������e�,�
���m-k�M,ޟ����r@r�_���v0�X��hDc�;�1�"�ĸxh��ʭ�Pg�7��O��	Q��������j%��f@���+αZ�!���r�:�:s���V����������pI<��X��3�;OrϮ���P.X�p���6�a`��`f;r˧��������G����u��'MG�����sf(S^�sU�
١����Q��Ew{�)A?���t���ED�$��RL[�E�����r�΀�4l7`�H�pϝ4v֯AV��s���FY��_?�x�#��� ����ݬ��%o�b��W�Ѹg�a A=���D�]U fG���
�<	�&6�w�	�v��d��Ŭf�o48뙄�O1���i�t~z���/���$����v�M�t��"~
Z��s�\�]����$"9Q��TG� �B6�aO�*��\����
�*Z~��ݮ�Nn�ލ}B�o�G;����ղ5�?Z���Bi��i��_<�p��a���S�K�^x�[����/��v�T'�aM������S������ݩoQ�|AF��i0�=I����ͅ+N�2e�{ߛ�z'j|g}'s!���T}vP'޲������8��זvj�9R"�&Á���b �Y�O�˒CX��_}��s�!���~��v6��W�O�J9���,�f�i=[�z3��,MUWL�:��՛%����H?�#���U"xÉ�Bc�X��~���ǆ��m�Oކ��9'6�1tz>!���8]���KI�X���d�
{�Y6�L�����-�HG��l��3!�g V��rXA��ȧ5H��7�?)=�gU����f��"����8��|N�vb˱ ^~��*��=�I�$:�&�S'��ԃ�pJޒ�w
���o���Ռ���4���*�h����._j���Zs��ӶQ�҇��G�����{7=�ɕ�zv��$�:�a: `��A5w����r��ܮ"n�#^��@��a��o#�۲8�D�����z�f����w�w���s�$o����!�0qd�>���+�a[�P�+����/[�C޳�,��K8�2����͛I�6M��s{��?�������^5�*Hʂ���h�%�a�Q��ճ�v�hMI>GO�ݹG4\�2:���F���gV��?��ަ��`yэE����61M`�1W�F��x�ު:d}�<���b�����<��/g@y߁)!z��$�U��'��H�إ�Ĝ9%�C-r�ވ�S��m5(�_,�k
2�0\�(��M�)��cr�m�̦3g���ڻj�"�34���;v���N+�IH1�x������i��Y��,�ǘ_]�G3h|�l��R%Z�r��G�F��t��&5��P����A_6�|�	�� �?�\�t7�J�"Iq}0��X�����q���E'P��b�:&xG
�=��V���2+�1��,�& �=E&Dt��$s��Z�T�7��N^��@)�Qo��#���
�H`[����Q3��@��������$L��]�J' m�:�Sد�
���$��R���� ;�����^*�X#�	}�G�Q5B���2/����q$b�M#�ڼ�y��O-�}q�O
	��
(�M�W�F�dhx�����2���:��SZ�kԬiP�0�`"-~v�[75���_r��f��7y�ڼ����9�ă�u���x�bt���.U �"!X0�I��[Y E�wX��4�`%�ο�~;6;F��s�}��{0?����
����O�M�]|N�98��DДE2��C�&��ܮ}Ƞb��w����e�ChY�^��`X�M}������y��>�"Au瞰������>���&m�����W����/�b�SWh��+� ?��M��w+�����P�_�ʓI�����o��X�b#V"�������HLiݶ)~ޚ �t_$m�=��a����3��fo�����Y �e���H�4�]��sH��{�s��n��
a#N𬞄J�q��h����N�%=v��fL�e>����R���9{ո`�b䭎��M���.a�3ވ�=!j��%�t[��.��J�hu��@�W�ڶ�3�4b�$�A��� 4���vn�z0䬆`�;U������gH-�jvw�lfV$ߥLo�+&�+����Y]����%0q�/̜n�*-D��c�o��c^Wm(43�f�m�SJ�[M�(9?<�գq�;ɑ,�P�[�EɌ�5\Ac�J��0J7{�Ҋ�7v1�Y{��������xr
2iӆ����O���A�ѡ��:5��0x����݃I�4�e��
#�gɧ�;ȣk=�'s��Y)����:��q�����޲�68�"q3�?M3��_��#fA(�W3|���Ȼ"��`&�XL�4I�������+S8c{By^DXӯ/(�̠���9����	�ǲs,����i��L��gm��-E,ޞ�(.�R��,����Q%�4�l�����$�An(:�v4�▀�Բ��������5Afb���x����&��v߂���,�"G�?FdK�W�/�x�ITB|˷:n3�ș�+�z��zl�j�B���3q�a� ��(Ö���<��IS\� =�5Q�q��`L��'!V�����b��:5���f�3�b�lj��o�Z�0$�[����ZU虗o���kX�{�,�7�֜X\n o��qmV�j�k=s�,�Qޔ�)'��I�~ϫY�=I�����{���G��ɐ����X;�Xfoc����v��0���oV]A��aW�q�*ġ�r��:����9�𫩣�,�Ɨ_��TF^�>��"%Z"o�D-�h��T����O~u�?S��Q�`��'G����M��^h�5Hu6��9,���ܞ�%�����ox��z��-�ߵ���N8����\�-�O�Aa�A�tQ< h��,�g��چ� �Cr�~��R��6<f�h�B3>'ٻn�3�'ܼ,g[3��f��>[�!�b��F���ЕX/˱K�m�O/����G �J��K �kth���6��qN�r��_��T'��x��IjV'��UOB���N�{�h�Tmt�^����8����ֱ�!�5���Ɋ.H�踶�Ȋ���
�����:�����a}.<��b���bA�"��u'7��gCx�j�s��N
�;6~�����Kz�J�cZ��~%���G)Ȳ�p�/�gBՈ�Y�1��p�IA�"�o��f�9a�U�b��%���N"��j�G �y�$Čg�ܝ����l^$�C�a����<-�����=W�f�XY��>�Y�QE�j��VP*ӑAwqCɀh���w��~��f����ˍ`T��qPj����������临��̥�p���G&ˎ�j�B��ሼ��I?z[�4RA!L�7\\p�d+�Kނ
�$.��;C쯜#U ��սPRp�+v�u8D�4���$�����&� �۾��d���;]�J�>�e�������0����%��X5��R��I�يS [u��G��b����)C��"�1�@Ɨ<!�˙����N~�6<h�͜���2����ͺ�����@b�L���-fy��0\���<<X�!t�HHd8nTùX��*�8e���,�u�*�4�Mb^%��$X�$)�J�B�̵c׮Y�Z�$��(�p�喳��4�4T���55��;y��3��-ʃ:�$�$�����ô�ӣWĪ�R�`�B��Ϯ(d�G����R�ǃ��Py�v��X��4n�����t���8[���V+qد�m)�1��*������61ӿ�N=L�\=z�&H&���t{�C�:� `+�� ����/�2B�P��c�}��y�a����;,�m��lm�[4�L�PȀ��5���"(�,₧�rq�2"����o�x�t�����L�JB�F��uMK1_�Z���
����l�g�O|8;�=\6n@`�k^ZW3� ��)�^XOJ/�9m�Ā5�{����4�)	d�\��5�}��l����Z���iaϷ�(fG�Ik�_V��^��~��R2	gHt�0~�y�ƌ�9���q����;�֊��C8�Zy�q�v��ѕL4>��#��RBc��<	o噖Ӡ�)m���l�a@�~���:'�B~�U����w5�Cj�]"�<8�=���K;��~���RI����z���i���� ��&�p�f�:��V���m_p	��W�4��ը 4��o��@f���ʃ�����8��{�Gj�Mk��c8;�d��X�h����s+Qy���`�H��E67��ܰV|Wҳzp_���& �b�0�F�2����"�&&�*	^)=ꅪ��t}��x�C��.�PX���߮&��׸@F�)O	1p%�Ͳ�nsnƈ��a%�9���ܴl��a����X��8�:�Ĕ��:_�F��?U�0��j�v�XX�Y�R bo����'���ծ�5�dۡ����t���2ÅV!>F��ˋx�W�>������ �`\+[���U��gz�{�a�)U"܎�LI��T�O��]L��v!��'A���=�)�U���	��<:1��˔�i��q}*��j�H��ذ�I|���l �����iJ \�Rg��zK�}S��W�I��WiS��,s�J��v^C%�+�?��P�Y��|D�c��h=��ֺ�?r ��n�_����E�G���K����ɻ��V�lV^��幵��cO�^{3� "��sE�P�^��6v5ZRX�"�?iӪE@��������c�f{A���Ss86��h0�!��.ʮ�Y�Z�E��ׂ�L�-�6+�~���҇i����� e�x��s�6`��Gj5�>N�f�(\"�<�cd��XT�Q��L|��{�}d�����f�������V�"2Z�7ظezlj����0��8��h�5��q�1�hz�s�g���>���B%��Y_��v�#�	�D��a��U"���,C������:�C�U �=>"{f�.
$�rJk�4O"�ϧG�Y,SJ�}57�w|�En�F��/�ˍt��5��Z��+���%.ٻ��(�0���]����Ψ
 G��Wv���:��e�p׾�{��%+�����"՞i���V.!R�O��%klB�[�8�&�y(����xD`�쾲�_�9a��פ��B�;�)��w���d� ?���I㋂|�=K�ւ����kV��\��wf�F�_=���qUߟ�u�w*9�Kû�=��{׌�Zs ��^P�n�c3���T�<y%~�0�TU�f��i�g�aج�0H/j3�B��¢���,������Иh?�ꈗ)�����JX��[����c�
����+�9洷T8����h��˖5��⪸�b���珥�lϯG���k���H�b�:.��w��_��CMul�"�5����}㘄QԂ������PN�ݧ�.Vc�APt��'6ؘ�Z�='��\h�1í�t\�f��|<z�m+J���x��ֽB�M��k ����7��͘�K\'_ �@�k��"TpH��J�ȩCׄ����n��B��Ϝ<�ߍ��$f�3ö4��Ӥh�������o�)~�+����춺g>��L�:���U.��>�FC-U��QC(�H�gܮ�<�LVZ���qe��򐘙����WU9��/,76R��ӑ�}ˡ�B��׎��d�J�)���x���fzQ� ss_�^�|��9`�R�����a�67.7ԦT�q���U���w%k��U��n�=����l���P�-7?`%�5苦����6�I�O���֨�(�=���������,�aj|�������$B��L]n��+��ǒDrO�e��1���,2�h���;OÊ6��{��bv��ED�
>Ҋ�ԨWj���P�S�*�
�3���XQ�2s���&������;� ���v��0�Xq���l��7M�)���am�M;�J�rss:5��g�r1u%m�N�S�_;�ߒ�>��.�yU�!�&��{�zp.)��f�������|��"U�dB�1c�P�7�i���1)?,�g���),������:�@Q@ji'A���������/Ѭ��,�7��ϡ%��a>�N���}uV*V��F�H����}w�o��7Y:���XA��%�75Do��.;��ɋzWc-#���bOn��W�/h�2l�q@�tiJ����}L)DV��O�Y 3&������7د9��/8!(7������iW�9��E��>�5����p���7���;?����p�$��*yb;���i��[q����#��p#�WX� S'�u_��r@�q$,��:�sec8t�,��0P��g�:a"m�l~Z�r�2�r �cE����)��	��S�#yK�1E���|�]Z�!�����VQxړ#��_l1�,� �>�)�.�pG'#�
��y��LDɞP�7��ٝu`�8j��H��+���W���RB�u%p�&_�ȺU�c�w� �JJ�~�}�_��a�s��R�e��.B(�������o/�r�@#��ݓ`�}8�İ�m���5k��$��n1�{|r��f�v��"H�#3a2�t!R2X�4)^i�R�Q�%޷�u}�oy|t��H�_��D�4c��L㏊�~9�O��![��I�:�'���Mz�/2Œ͋b�T�_��cv�,'���
RR+gCN�3���_����d0,�I��"�~|��߿n?;����G
�1�ذ�%,ն���;W�-į.mu_�::���f�ܣ��كs�1;*�jv5�|���7�_Dx�{��N�FW��Y�:pji	�e0Ⱥ�<���*��mGV'm��E��Bp�_ҝ�H���L����	"�l�q�j�q�Ӻ���t����Xk��`O���By8�[(��A���:'�����W���6|U۲������e�1E��U�%J�����o�_���q&eM��F(;��)U�_�Əۍm,��^6���;'r�ѡm>c �G�l���_�&}��G�x��v/7����H饦��_�\Sz+���{�~}�f/��c�?�ib�4H�b��k�읓EKP���̓-��"X�AT3F����9ǰ�)�C����S�m!��O�5[�[ޗ5���Hro���a�>��x�~���ỳ��NQ�΍\ۈ�q��b���OUa��is�1������խFC-�� �n����4�u͝�9/�!�$zq1el&�d��J�5�3ּ�\��R���mz��*��OS��T?�����Z�UR��*!o�Q�!v1�K�;�3�k��nC��1�ѝ�"T�p�h��kQ�rA.>����i3*�Z)�4��$�J��RJ\�g��M�7t�U��A�n��l�$A�;��p������`z�RWu���d�Z���ĶS��@̅P8��0�Cdj�G�'�0��v��>�Gh���<Ba�y@�)��Z��Ј�璭���<#�;u�G0iqXqN�I��ʾ��c\�2Uhx�/�S��S�a����5<ga&4�0�N�)���`�}����J�Ͻ��.�*
�_�اX��S��kq�������Q*Ł�%�ס�wL�B ��rS ���p37��δ&�t�2��!�[�|`�h�MA55$�yh,<�2Z?�;^z|ǟMA��XK�	7߽dF�,B݇kY�)�`{�����h�6�V����� q�w �K�����j��9���3����F=����<簼���\�$�AA�ؼ���>ggP������$�]3� �5x���dk�Xb���z��n�=K��;�׶����'݂����)mR�LD���"a�橍�!/�ư���c83�V�	R���JV�Gf�5@����۟}̚;�������4�����&���͓j�=�5�K��liI�횳2]��� 5E����w����`2z����I�9T��yY��b�����2�����+���C����`s�z��5���/���uh�Ķ�
�̱9׀e��:�A��@p�H��Fv���� U2�A{�Q�I�T�F7n�ݓ�A!x���w���塁mq�S2���9��l�&�3�b�ƒ;ekM��8�o�����[4�e;����g5���
����	M&�>������cԮ�b>�����D�/Gd#�qO8Ѩ�c�9�(��`�̇��嘡�n�֩p�¨�U����1ː�
������������=�[o�K�B�myK~�� �:�c��՟��'y�s3�@T	<��L"d|��s�@C�p��sP��H,�%�d�֡�	�0@��R�GՈ��J���������~p�T[|}E���ժ&=�7���Ȟ�aT��Q�Щ�Ruj��'l�T����v͆��M��fOba&�"=��t}��H&8Y���n B��0���o0�{k�Y���t灄���B2����Y��
�0P@�-j������9�N}��1iFAL��I�]�'o�e���ȯ�:�'Onq/!���,,.W~�h�\7hm[�ҋ	OZf=�z��*���~e���G�#��|$�M���U\A(���ؗ��&�Xb�"�n���ǫ��F�C sn�é���'37���4���zxY*���X=i4pKiQ�� ��?/�V#����y�����B��*��&�X׾�0�$�>��J�=̀eW����'��ќW�e��.]''x�Y�]�5C��ke�1Y��o�xm�[���7UW��df���B�Y�@�Hj\�2&�����0㮚"�E�GU'G&��=>�0��$���ٝ���x�#������evr���;��U����P�u�M�⿈�n�D�?��_�/J�3��'W[��k���>��^r�gZ�j�$�\XP�8#��@�	4S[��ZH¡_&w� )����|����b������bKњh1��9`��?Ԥ}8��y�i����>��{�H��ǭ�q�L���o�j�*6a�hr��/��=n�\�L}�<����gT�@P�#���u�YgLk�<��*�T$pk�M��՞��xt@������Q���[��f��#�ܕ�2%�&�>�]��g��ߥˊ�KO�Ѵx�zq�����ϝyЌ��W��֍cX��س@O��:WD����*�)U�(�/3!�8ȍ䓌�J�3}q�*���[���G���&���o��4w���me*xd�S��W|?�	]K� ��('��~**�񕯦e酞��vCR�!l���Oh�rk�De�����m��Z�OJc 3�fB2��ݔY�{���d(Q��2aV�8rc�`'k69a;C ے�4@�<+rG�)h�B�a�!C0�@�JPڷW �TW��.o2kZvऐa
�lXwY�ps[~�,���po��-i���sޣ�a�u���4?��V����R�|m>�D�9r�Ɨ4��T�גek�rb�#��Oq�a���&~�g���rv9M#�sVX�.:����p����L{v�$�s�ܠq�=�����,�����:u�$�b��������x�:����Z�k��K�bX1$��6JB�⯲��\izB�<-K�P�}��7r�Q�d��S�����l��Ɂ�Nw��j�SS@�Y��f9��M8rA���0�^˻	��w��΍�BKx�n�$綍~A"Q�:�=��~��M��M�T%�.�;��Pj*�E/����6FMC�4$K1�)��]x|y�Is#P*����r�ۥS��So��$���Sp��x'pD�%zq@�E���ba�t��"7��������H�;����h�-pً�o�{ ���T�y�y�|�\���b&^F��1�5�4&O�<�fPX��z#�Rc�UW}Kj1���L�Nv~z����$�� �Rq,�ξS�Ȍ��+�� �����Q�^$�a���vz��P�@�[`P�C���LY�Զ�1bJ����j>�Zk/�:嵊���9y}6���ZY��Ѹۼ8�ܬq~�kc�-W}g�Cuڲ�KX�%�"8�&N��Es=I��yeĩ����t�6|�Mg��TW�ƨ�Tq�Y�`lo�a���9� v�;�n��!���s5��qK���,I9�y"1��S�
_���V��`,s� �;��֦��/*�I\�h+�2;��{\�0����+;G��T?W�)�Y}��v��n���H�2	�啚'~��5dpH�k���v�?���n	#Ϫѽ>c�+���E��<'7c�����d��������L��<Cz��J��3tq��kY����ΕȊ AW��j]�������MZ/]�^�z��V�p2���������7۱�S�*��T�P���p:�o)���Ύ��]C �>Wl�Qu��M�j2�D���wjv����J�XoX��2/���P�U��h,Jm��+/*��P��� zR@�r��J�(��}7J�I_�Qu9A�x�Z��
8	M���F��a/R;Z���E$���у3�`N����z��+�5�l���]��iF�ɥ��%��9�#[�`O0��H���Զ7��_u��.�cQs�%���Y6���Q�X���h�nL]��puF�����)�V&�!�z�$�:V1�Bn�/�.��Z�U�9�N�o��3,Gps�4A�F1cϯ=��l�@� ���W���X��0�Sz��,hR���bq>��Ę)E;`)���3Iw��\�8�?��G�	�15�"�x��(U��M���1�\x�d���1kN~Jl������|x����L�$�{�:`7ʅ����<Z�{��L�Ru��K�8��$��s����0��/��/yr^,��݇�*M�����E~�Ϭf+�Xw:�z1� 	K/�K��R�-4x���U�:�D�IҬ��>n��pֽ�!����b�D�v����P1�h��MlC���.��a���'�hok��>�5������JE/��g�r��zr@�n�xX�@��=�'�P���P�K]3N��u��W:��*�� 垁�͚߰��7�>�;ؾ�=�>F�Y�fLr�=M%/⎻�q�m#�>�J��SW3��pE�P���M֔`V� ��)�����P�f���P��L�9L0���I�YYVX(7��,�0A�bs��HIG�VD��
�J6��k���ʎ�
+n�f�2X�(%�B��d�n:��@�YA�<eG��~��2@,9忟�;�j��Q*H�#��ӕ����4|�S�D+���k-��Q��m�{-�($���ZFr��-v����y�)����$������ܙ�3�sq�W�S�An�ͨP�a � 3�a� �U�e���7@9��!
=E	�gnDї��ģ���~��ЯpH�˴ls�5n��3�&�T��>k��{�n�(K/�o�"*���S0����u��*-n�"d�#�QW�̈́w.B>YW�Y�`^CqM�c�����}|�я�ă�;8;z˽n�QzQ�UP�Z�^��ۚ�N|�JC��}7<|p+r� �����0'�(g�� ~��:���{��������Z�t0�8��^���.�<�: Ha��G��s�61�Q�c�\.�)�3'�+�8��s*;��1�tY��7(��6�mR�'�"w��%9�=��2k�M���۾IX��sC��UZ����2{G�=�Ւ���0�ڧhW�:y�ź�d.�j��cMT�<�ݼ�� ����R�AL�����	vv6�[<o�P�/E��c�uJ*�F�o, �o�7�bh��N�8��܀2l���􆘇���Q�⋧Q:��\ˇ���-��F�?ޝa&M��.��K�K�O=T���\x�P��u<�&r�͝��@�E��g`�w�sn�U\�0%^Nj\���ࣘ�� �~.��;����6�H���F��B�JF,��K����-�&��-�~�NP��~<K�3þ-%"�&����
��A���y�� g��˹�C����N9���9mX�`��U�������W8��91�?���V9��߰���Ex;�c3�/`����5�y����W��+_L�\t+Bn�j�X]�2�b���8pE�M΃h!���V�7�5���c�ү��@�[j�__~[�O�v��[lc�(�|�LN:|5A�$M���\�S�x%#�CвP�PN�)Y�6�0�mGd�ە���elm`7I�b�����<�G���(�1Z���>�b�z�]J��WT80�~�f�w��ŉ��%�l�˺YM���࿨_�e#��}�S��7��C��K��%	�)��i�[U�܍�A3	x�R�z=��D�5��r���0�؝9�Rh|�`�W��?b毺Ǿ����[
\tZK�m�Fz̩&K�^�#L����n�Wd:��������3�$���ښ ��+M� kŅ^��-��U��z6Ԙ��U��rvz���$�t⊀���VY����&k�?	u-~��_19V+�b�xЧv� [ul, pB
(H��C��9��.��?�arv��JV/����b4Sl�����b�b��%0�@�!�	��KTa�N�Nt�;�Z.-���Ǆa0�8�E��07�O�p&ハw�I%�����|�שie2�x1���Z㴛��}a{8�kB�{�f�U*s���!��\Д�3r�쬐����_g�@V
P���ͱ��ms����їY�R�5��������s��YUɮQS"Ig!�ZAO�O�����:.)�|+��z�}8y�K9I�௔��@���}�� )SHb�[��(텟����V��cU�� �?N�F�����a���l�dc=L �A�/[�:��\e5����S���6�+��ݝ�<q�E|'��Ǝޛ�������TAvH:���RJ�bH��{TlA_yr��X��ʥ/C��s�C�e�du�7V,kPY����F�n�����,�MY���Yp>D�D4qg�oVZZ�7W�50M�ކȣ[b*@�|Y�gm�`s����U������[��_-��ٸ���^���q�4��l�����uc�����P��#�E���¯絼�:�eß �)*=�@�&��vt�;�"+����B0�0=��'����9?�K�%3t��<&@X��ՇF��	@1�{�މ��� ��ʩ5�x����v�V_|�ie�I�r�7��g#�i��÷k�[H�1 ���rĠE��z��"��t��g�F�S�a�|I~�����#ǎ湐���Y�Ѧ��r��m�s�X����X-b$9μ�3^v�웭��YY32��%�Ao�d���q���$�.rK�m���5V��B��j* Ӡg�N�1�)9��X4f��nU�qĮPZ�S��8Ki��%֢]{�;�}�G"K��(�a��}Hx*�Q�]�V�C�6���r^�z�,as[�Yg��BC2m`��@��/z�St_�g ��)K��GSv�:a�9��.1_�1eB�.-�.�$�k~����cc�t#���t����=�&�s_Й)ȡv�%�[ٗ"e#�ѣ˩O]�t�
^/�m����͂�ø�Nr3��p��94H���?��+�Em�UH͹g�8/����J��I`�0g,;�m]})�B?R��	�PS>��Ѣ�����^��#޵��ռ��B
��f�5 �=Ta�Ｄj3���{ҧ���BRE6?�ƿ�����c �h}�.���[jk�/����z���D}{�q�*� Tʓnk�jY���`��~��wQ1�i�=���^ ���w�Oy��
�[��l��Q��5�X����Q��)"��V�0�ȵpr���Ӿ�{t��wf1�rI�=���n!`�l���g�Lns<��:P��p�H"�,��`�+=�wKa��X͵���6�+b�!"� q�9�
��|�<^ľּ羦��k�/z���I΁$ �@��ބtdU��!.l\���oBu�<�i"kH�Ja<�w�>�x�x��~1{x�j\�����*��k�$w{�ۏ[T�L�DB�ͮ�Ε2`��{�$I�}���)����'��n�0��ym'"@�qЗU���A�y��e���vT�j;OS��4��|�jnmBUN�\��v�����(�V�V'~B���px,ȭ�({t
�䦏rj��W-1��s�§���È����x��v+��/N�\ |b��TоiG)��6��a�*#3�J��Gm�b�~��������TQ���*����V�ϿŘt:r��֗�5@��$^^^��o��K�B3��!���'�!���f���#�ǃ?\��J�暠��E�Z,���N����5][��;*���D�Kks#,P���2\2��K-�]M9_���I؏���T������p�
ᖅ�[A��q( �p.����D�v��!SP���}���]�����h+ͷ�U��ch
�	'���r��lkƞ��W/�݁����B�ɋ��Kc�Q���q�_ �����՗��-�����B�)𭋽��:(�.�\��68}'�! ��٢�Kp:����J�^��fZ��O3m&H �����  '5�J��q�j�<b�UI4my�)�4�z�=�=s-��jv�=�L�N4��]�G,�(�-$�`�$ F+�
���5�Q:M�(%�h [D�<.N.�gj��P��I���;���@�'���C.�p'.�c�6��c1V���[.n��{UeZˣ������d����g<�
��� ��� ]�~_��+w5/��J�I�%qU#�5�K?9�x�R|�e�/_���٬�۽��<,���YLz��iS���tΡ� �-Ncz�Gs������Śj���X���tx��8����H]��Ќ %�]�k�޲�/֘/F2�hJ^�[7�P������oD����Z��_�Kv"bT�.:���J �	l��oM�p<K��[ov='����*up�If�ht3��S���7&��e{��*�������x���bT?����+�6�c�@���@����[�ӥ�2���)�ʢ=��d�MW�
I=��Ki�z�
h�bJ+�����i:��Tܜ��_b�����eK�� ��Y֓?t��ڜ��pw��8��U��v�'[_���l�`��1�.PX�/@^D9Z{S|#^�T�[��@b%��;�Ir���4͠��^�k�������?=��I_q~�@��*^���Oƶ5��׋?xU�V*��H�76�#���PЎQ������%t���m,�닭�q>"��f��} j���a��"�?aP�����Io������h�- 7�ސ��r3q�A��J&c���Ӓb�|�;��sir��;-������@�� ;)P�z��>1�E��TD��5"��d�!
V/N?G��K�/����:}Jy�nH�yz߱�%��ߞ�J�MK8�΀����o�[3����~{d��q|߸^urk�hﲳ�^����������O����W����\A4zX�TUL
{Yl?��	�?\L6@�M�N����4kxvry3�pKE�@`��
]Ej,�w�׬�-e#��~��.c{b��0���l�sV4���Ѵ㓁�]�퍖(t��G�#3;�ּE�q�z���l0R��أ��f�r��ŭ�/�t��kX��b߸c����i8�d�5h��7������-�b<np�����t���J��-[�	��}�~�j�s����tWٴe�x�mG�|�_ߋ�@3|�)�Y�Cz�aE�l O3�i�,�W����U'�B�7֚ؑj�uW�jY����p���¶��n`��"N�\����2�kΖ��<����e	F΢��" ���P�}��QM�LJ���~���bϰL�/�dIo�1���&���R<X:g�>�n�ZS�<5��Kb���._:�#©k�]��*oI�[ `2�y
փQto泓���x$%���4ip>��`���fqt J��G�<<T6�?����H�W�?�Ą�\���j�Gݍ'-��ʹI�m�%�e[7�^�4�a����&�o:Pi:c�0�t���:�W2&���󦁦_�5�5!
�)���eV���G��9d��~�ah2��`�D]��t/�i����o_d���Ö\jI�e}�G6v�7�e�"�s^�&���?H�}��qz	H�׺Uz��<��F��Ą�خJ�o7�Y�zԉ��	�o��	*�L�O|>���GL&N<y��N�+�F���@	~�
�M��	f5��,rF�mXU�s�����ta�o�ފ�v�j����k�me#�8����U�5��S'�p~�ĀS��
�j^�ޢ��OB
o��%ܰ�9�	 ̤����h�h�	�[AC`=�BUE�{o^B�(�:Ǻ����%<��7���)�"@q�D����H �����do4��>�P�O�M<��0���"��[�(����X�π�O։9%}-M��q2FH�8=�@pZ��x�U�$B��	��4�_�QZ}n����P�0~�j\���0��8�Ì������C<Z�B�ŖC��ꥅ��L��,˛�!�N��Q�_��k"�� �8X�)��$ hI������n�[�G���õ�S�D�����}D>�i1����zٕ�]�����86���^${��A�]��WH����Qj�g2�W���a	�Z�lm]�U�s҇Rs���j+Ԁ��(���d@�#���� h���>N���V�l��(�?<��X^�䝞���D�*�RNU-��m����dH�lͲ��<V�4T��!'��'U����o&���02$NW��v�uO�up�P]�T�*]��fn��7�V�2��[L8��)w1�&�BS�}��W(��=��b"��#6��	���{4z��d��sèp�p-�;ܼ�ڔ�ѻ�\=�]�5=�I'�+�<��LS�;8W�� \�MA���c�Y��<�k���&8�vg@�)���v߮T	�,�T��&�_0.&�	�y�I����+�Sy�7Sh���srx)#M�5����U��aE��ʞ��݇`^�h�I���L}�O����v�kUB3���~�w�#����"S�s&��S����ݲ-ΰ(��Ka�Z���J�<߰9�he�rfkbg�B��IO�4�N�1/ɥ��^�Vϭ�d5q���eaޱV-��O�u�ґ��EÓ��]�_� J���$m9�ד���HD��k
4;�����1F�ٰ+QR�4�) �a�:�����Dn�R$�M#�JC��؆^ś{r�5�fgD���S������c��X�W@'����B�R���u_!���0����\A	o�KLF��6+iD���471��!��/Ar�4p	L���&�gA�S,_���i_~xl�C�sy譍�Gl ��!��5�����&�n�_����X�y�ꜧ�*��O:5F���Ns6���zgJ&��e�$]�qa�yv�e�o�Ʃz__��=`�w���u��c�u�m�v�[.Dp�0�0�$�
{�<d��w_vm���pRk�?��vȪ�ʕ��Ŭ[B�b���u��"r�a;g�m�\��v�k�՛��:9A�h�7!�x��K$�w�]op_S��]|*�jyf���R�˃��U��n�x"���qO��7_�La����܌7�ŠN���پQ�_�0m�~�T��jt�؞��?Z9�scj�s�i��L:��65!��b���g�޼K�NY�����A�t�QӘ2rs��wG��d
m���T2k-m>BA��,�X~,/H��'4����<g���׬�Ւʋi�l�\�	���饖>Y��W�^o��B!�;�+�"{�v��U�` z�5+`:�D���QO������('��8�ݓ��fR���]����&�t�ŁE���n�.3>��ӯ�ml��}��1o��p|�[.�L�
ݝ���i�&��&�\S�^�В���@%}���>A�c+�oJ=t�Qu��3��Ȫ�Q� '��^�Lgi>U�m��	�{��W	-�}e9n$ci;:��9T�ِb��%b�W�7�5�T�T\yPuV_y��GhVjP��}���7tm��W�q���CW֖�zi�K �s?R*�ŷ+*��@:(4����oX�����n]g���^.�"�km̩��\H��Zy<������ZkfS�E`=B�*���������#=��4�Y��JF[
\F#�OŴ΂����Ҹ��+�VG1��#��MP5�I|L���)@Pه�����7�-Ȟc�_�V)��W�J�G�^�����'P��d�;�av��D��ܙhK��Y��H���l7|SO�6����z=���K�u^�'x�̚��2�b�U����0b[O�f�(�q�z77���3ݰ�j��LĪ�|L���"��=&�b�1)P��S�4�[�i��yX1�5w��ޡ&-IM�?n��n���)s��D�>��qK����733����k�E��H7�u���xC��څGX]��~^T��P2n�˿���fU��Q���m���ڱG�i	'E�r�|��p?d�v<�=/>f3��3�Y"p�TQuu�/� ��Q�+���z��O��H��`�8���H3���+�"^8�a���SL�������r`W�@���!T��xqH�=����C�ܯ6�#�=�l�0�Ĩ�=V����6�͹�ۋ�����T�.p�e�����9����5�<�jS�b�hF,�X���4�O��ћ�[��rm���KПж����_����q���� �:�u���I�&g����&���G��Kh����D��Q�]�<��������Vg�����cT�ؓ�k��GK孾��r�[Ia����+�K��,}q�n;0�	SnX
@��Y��/U����TM�x�zG��hki��!�Z;�޹�H���.�\�.9�2����@
i�7��x� a0K�%P����V�.ߐ�1H�祓��e>m�2�=s>&G�&]*U(,��G[�|��d{����{�������l|-@3�B�8����Qا�w�</��j����!��K�s�o1YQ�f���-pECE{�Zc�X <S��Y ��%
��iҫ0�Q�RL�.h���R�&KR��(�' ��}K	�]�-O�EP�I$�㙠V~�9����|;� t���̹2�6j�jq����Q����_j[�4`g��	�,%�!|ޚS�;��,K�ъ4�r�)���C���[5��z���H͞���뤘�[��=����!;g�Ff'r�b4p3P4�Ǳ����C�x��1�'�Ϫ�(��N�uw �y��w֯(�:w�pS4��$�Ǧ�z����x���jsiqi9{\���C�PM��z�I�S[��Z⪇�A��l\SP�a�"ဋZ��Q��a)�І$�He�I��� r3�o�/���I����˻�P��i�'���~0<�F�3�JڰUʝ���8��	���!��u
 ^�p{�.��,T�=�N��@����k�ﬢ�i(z9Sօ鬫L# ^I^s��m�c��QSX�Ӽ�[rx�j�wz�|ĂUl��cgF���&)�U_���Fh�{K��E�S!nΦ��[[hB.|'�}�7*�U+�l͑*&̂KPjm Q�2����gsyG�.(`�ʫ�����h�o��/*Di����խ��Ȭ�9���g<x4>�7�t�C��U3{T�T@�ho�>-;�Z.�~U��F| �߈����&�Q��l��ik����y�ь��f9�T����.2�:Iq,L�#���5g�\il��=�3��]?�z;�$F��|�m���2�]SL�/LZ���̦/���MFd0M�94[�˷+�����aa~��	���7�9�_�@z�v90ȃϋ�ˈ8c^s���	��큘'WS)@Adp&)M�/F$�=n�;��KY��?���&nj�a���[����C#{�d-�.�h���}����B���Wl�@�����|@>Q�8%�fp�QH��Io�A��N�V{b5���Y�&�񐰑,�We�եM8�JY�yd�1D�B|m����R9��ݯ;r�"��;�q�X��#.�6>����vLaץ��qS�����
�Ow-���uS	��$�u56�A��ӻň�kqU���6�kG���+�2�:J����C׭ ���j,��"�V�Y��1��f�>��@,�y������4S�t��G̣!i��W�t>�r�z�<i�E���� �����0/���	P�f�u���H:b���U���?���V�]�R���N��'O�m�.S��	[��t|�=~����ݻ}(�i"u�2�e
���)�w�o�d(�d`����lr�"��:��4m��<��f���25}�Ph#��=��pU- ��:��(
�d�=��'�cU��|̠�	��cY��z�ʔ=~�!��Y�����OO�M�-D����?��>Xs���=k�;���4l��I��-/�*���|RY�̤�V� �x���'�?N� W)��7쒰���Ǧ�(]JY@��%�Km�w���`2����q����%��}����?�H�}a���l~��ݾ�hv�7b�!�h7�.F����i��zCQT��&Ә@�nG�Ou��3�/�V�a�ȃzT�ֱ�%]C��{H'cE�
m	�r���u� #/�i�k#����J=s�+���[yԈ�l�#�<Է��}ė�4�Ӏ����%�T�r�^?HrRӃ�����q�+�8���sj����Y��SClTr軬�>��-;�k��r�{�m{�煐*w���O"�^�bp��'����7���Y=<��	6/˶x���#;����k\���7+������A}�A����gȐ��ӄ½ghN�ޓ�/�2��<@�+N�r��+�ߐ7E3%N��RP�4\-���c�.�=Cȉ�Qt�a�]o�q�M<���ﶵ���`j�5��7�d�F1���0�e�NX鬗��`��e����݃|����;�.�F,�.Fe	��zQ9�����E�sωp�I�rB����{�H�V�����p��l�^=i��^��ce�mV:�Z�~��^S����>*�`���M}CI=o[��ȟA=뗠����b߱����ыP�&Xb[��r�W��[5Y���X�`R�S��6�Sq慌?J�C�>�Z��������<���+Z\N'*�x��u�3Aײ<�8��g�l�6��/ɯ�E����)�}Yb vL��A:>��h���r��S�!�H�b�"�kp�6j�ﻇS��e�M��1#N�;QR�X(I�X6��WV��0�9|>陒����a8 +�jz����o�y0�n����!�V�R}�E��æ�.������ڴ�#y��zC3l2WY��Tu�ojL�cɡ�f5@ˇ�
���%*31�k~��r�xr{��9���0	��.s�Z+��Z����:�P�Cx�l��r��q�~�Mg]P��l�OSb���y�!�K��[�ц*%x27�'�=QҐ�l��k�cP�S.WC<���B�4jgs�.ґ]��j?lSt�'n�-aR���¸/*�.��81��t�\l_��ç���$<	t�3�%�E��:r���.�(ֱ��u�F�+���n�������:-�ein�6����5��Ya�j���M�1�v��=�ܼodr\b����i��ڏ����4��+�Ɉ�}D�_:.Ĭ��o�����)�ge ���5�Gq�ئ��������(j7��%I��?k��9�/㻉������Ӫ�"�K�I���_��$��(��Fl��Gg{� ��������叇�U0�����Ί*�B�Ć 	7`�w�p=�P�B�|c�MȒk݅��e	���Q��2f	Rܸ`��f\(y]T�읎�ZB�=�)R%��������h�vkqbm���Y��/�����\��߭W��(��j"������|Ԗxlb����o��f���~���T#�K�O�B�u��(����꒞�$�7V�Z..ʃ��6�� ɺ�#`�1�;
�O��}����;y��oi�.�-"�Tg��*j���u�͆t�%؂��7_�~>C���񲽫R`F�Hg:1�_����HO�����|<|�5������^ȟ�.��|'�����+:~bIg:����Q�G�z��O�q�_�+�ţ���LC&���/��s�.�b��fY.�k�����[h�8��-Uf�:b�sJ����^`�)�^��mPh�B���������Q8^M���=���������!��3Ŕ��H��2
z���Q�,W0������X &(������'C�����~�ң$��bB0��&��V*�w#Fo4gK��:Ï)��h��z�1�ظ����ѹ,V�YA{u�o+x�k�P���yB���w����@Oԉ��l'���D�iT�㙒O$��U!�]�B�eao��H%%����"�#v�j@�%�n����^�g�1i����Z_T%<�n���dΛ��%�Ϩ�����?����i=���̓SK�A;�;��l��֧��)�XV� �<4��cX��,VՆ6<�`~iz۵0x����2������%�����% ��H)����^.�D~H��E�H�+ B�����l��dg0��y�2����)!H/�tLz��v�|LE?vP�B�E�����{�Ғv��r5��a�L�,�k;��2��]�)҉�� v�Ay
&?�.�1Q*.ʝq���sp��ԍ�꩚j��P�=?^��Fet�iƈ���/.ʽ�	}{������R�Uw�������a,q���n��S�Ȱ���������O�����CQ��Ih�hs���$Ӧ]C���)y����5g#x�%'�+Y5�ؾ�o���G���Կ&5x����g��"� ��H�#�r�U�?�l�bv#7��o�NL��ɎJ�:��0����!�_�!�qI/��T�g�yYZ�y��?����!R��4�?x���X���6��ĸv"ٷhϸ��XU��P�t�!�0�&
.7����/*�t�{����}�N�� )_N(��9z�5ӛ�]7�2��on���3�״3�D�]��[�B�����U[2��V��1.v0h<����TsÄ!����Q�����7ۘ��9��
M�j�`�w?�l]�v�D�v��7$A�H�Ԩg�s�!w�I\��rI���n�nA<qG�إ�â�Z��_���ʫ�Y��Mv�,�{- �Ε.�d�4@�ʆ+B���2$
���XUR���A�k�bt|�Q]X��ߚ��^� ��,Q�)��?繆Oa�ɪV������Wo�L�Ѽ�=JN�����UTU%��T�i�Z�?P�+���F��Oc�%��<�Qa@�01
ȱ��eH��qo~�N��� ��h9'#�&$D�M��X�dru^>�ꉅݟ��<���v�gdd}��+�߂�`h���Ψ�\�I�^���A����1���cc<����`@Qv%�1�2GMeds�#o,���33������5ۡ�ׯd�J���R%�y|���֤�OQ��^T����'��k�)��>.:^�Stm ��G���Kш�+U���2��Znxj��(�����[ڒ����qq�4�]
����9�NZ�B�u���Wr���� �е蚾x��,k"��3�~
�y��:��Ҥ�$X3�H���Z^"á��`�T�<�P<-���& S�}ݤB��G��L�I� �)-�T�Ka��}�_$���B�Ƴ�u�	��A�^�ϤD;�Ղn%
���ʪ��+Cj����F���ʿ�C�3�HP�����qS Q.q�.z��u��Hs;��v��h�c�"�y�E�������0q�ȼ�1�q��F��}yp�5���f�<ܪ���"����:/��RV�HX�"9uFB��H�<�U�͛����]^i����YiV\L��>�v�C��}'�����~M:��ԥH�<�5��$���]8&�&�$�#H���NU�]�j���&n�n�<����(\���NYM���ppb-�8�.��u���<F�;��!w~��d;�l�X�젞� �,h�e\�x�v�+�!$m+�8H���8A;�0x���r��dْ���?����w�a�$�՟��J��E3M ��|����r���|��=��J�_G&Ǧ���!�r��yZ�c��r�"�ꆚ��Hr�_q�ʢ�NA��t'Q���j2�_!��09Eh�\�U�!z%M��z$��ՎoЙ}�l\R��N�/�נ�u�ݾ]V���+#���ϐ�/]���Y2c�b�<���N]`MI����*�P��գo���q�b���(v�����6�y�I�5%�!���l��͖z ;cr>�����]8������/����p�問ʼ�$�l� �V[�nFQXB��|d��?�({�VmŸ'67s�a��q��J��I��@�yu���<Sa��F�D��V�%p�3Ŋ�v���D��<d�˛2Y��7l��;Іp��ƒ��������V�EB\G�$½��U_f�a߰^��-mU��;nxw�pw��J��]�Ч�Z�h>�G�L�u��á��Qu;�%i�-�ӵ����I���`)Y}�bе����,���������'�[[�i��*�k:7w�\M�Q��>n���V�[tp�x�1��g�w�UĴ��M'L�$U���<I���p�)����~�
��d<�� ���b3������?|��r5Q;�=��B^&X������׮E@��6�GȄ�������P[+y�V�Z��/B����$S~w������G�����-HC�@v nl�B����Ou`0�9���Z�!��20h�����"4'VW�^��T���d��P���Dpw�yz)� ?ʬ0��d�lR��#��B�&�,Xo�����_��V�x��ˏrW�� Ce�?�L��`2kE�^���y(i~�!�|���W<�!� F���x�	g��8�j.�s5�5���e�������?�E{�~E��o�|������0�g�\5��̜7��b���RC����j�ٞ?�h2�[����[��fLT,�I�������N�$P�M~n6(�Wnc[k��Z)4p��)[g��Isc���\Bq�/�8RT,d�1�dD���MR���R�F�z�6��E�Ӎ�h��JAZ8� 'R��C5������3:��%:���2G��G�^��ۚ�a�ڻ�6�2�{��� �yw��iH�ص.ו q<� �p��8Y��\]�#���õ��F���#%k�^��$?0.ePM�e�_�(~��X���7Ly����%�m/TM�]�o#6�`����?D<�@�J�[���/���pL���hS��-�̸
���y$%0Y��>����v{�{PJڟb���;%g{Pr�v�.�gYֱ��E;v���Y��&�$:����iϾ�$�by&�eR�70�����X��I��흙��t2ʥoӔuk����:5���	���<��/le�C�)�SV˄'�P�.]p�(:NU�ьO���p��ͳ�2D��*��YS��"�&||wUB�Ig+ PZ���ҍyY��v�˖��Fõ
>7i��9��4�֋��j���V}�j�������?�z��B���#����-p�����dN-��M��Z��v!ޞ|����̲�����8|���]��:54�x#��5Z�A��qr3��{�ɓ ���@ێ�l
,�c�i]N`���N�QW�ˠ^�h=���x�q6�ϗ�'�zU�''*Ԑ�W�<��9P��($��6W(І�sc޵��?�İ�o8����t�m�m�ʤ��5��Ze+J<ڶ��>	�U��� 1}��LX��'���b��� �6n�0��bߛZg,��
]����Hv�=�9�WtX�j����d�U!?���%M)��v�mf3��4)b0��-Z���)�(6g��1%(d:=
[�v翱����TK^����Z����6	�0/%w@�g�_�/��˛��Y5�$��Dx��~�t\7��n���=�(z ��$	j4<�I������z!�����X��Q��O�/�թ �{/��Qu�?C_ dU���$�V7� I짽��j��7��(�)^j��L����M�үcmk��b�$�C9�a�P$��I=.��̦��n�++cFzՇ(!����Q�q�� ?rr_�S��S/��3TNj����Ft����o{ߚ��l2_k.}�qCI�~�^���d�'�v��}���_cn&�!��-|� X*c» w�F�b�����Nu�s}7*M�ɭ��_��sO�'|���0��j\��}��!>\�X�}�?�.5t�Qg���A�d��Q�e��p�x��]��j���z�]�\� !t޵���m͆q?r�0�c�)l�Z�*��e*]�L󮕣��ٓ��2��+k�&j��ʒٰ�<ڠ��5J�p���}�Y�%?IU���~Q���Gݸ�5��4ةgv�����pxь4�'����?�j7�aBT�-����g36��t�
�G��N��V�9W1�_���K+��B58)QW����z�ke����h{�H�J^/�
�Y!�"��L���b��iB��{�?�a^E�m3���\)7C�-1��/
��C�j���^���\�̿�%���>�P��j.�S�hK�a�
���c1ϋ�ǯY'6�����Z�R(:�l,���ye���ͥ���̕�.���9�.�qG�N��]��8�_�{��t
�pߙeq���*wEt�.t���!!�7
ZYV2�*��x��%�
�ȋk���O��c~(����h&I=���mU�w��mI�R��;f�����))�Cq+���-\��yK(� Ԅ=���!\���ͬ�E,0xS��Wnu"�O��|�oP�9��0HT>�b7��>Gj�A_|dJ�N�G�&�2�c��X���
�pև�HbdI��Ӷ.�E%��$��ӝ9	t���Z�꼊�n{?�᧗�^�ڕ�(��� L����W:5���r�:L�8�p���Ӎ�V��t�ŉE�9 �c�3"G��3ΐP�I�ѓ|*I�@Uv{��N���A>���2�B���#Ŭ�Yak+���sG�?�HD#��.���t���~�s{��bb�Z�?�B��r� �~�-(��|j�� ��	���9Bx秌&�׿}.<ԪJ�*�p9+6>�dGB�'����-���Y�δ�36_���_���?_Kߏw��<��EA Y��Icj?��� ��l�l��(����g�EAa�g��!� bx]\f����"?^�0)]E!�z,�����P�����yHǝ���J�e���>C�J,�2[J�gRm�*b�'��p�z��=�r�߃�	��� ��(���@�k'TS��iY�O=r��Y�a�T�V�޵q�Iz�+^����6��{Y]�ĉ�]�ĔZg�hu���y�f'ϱ�5A�/S�d �2��W�hQ⢸/�ÊL�Q~9:jM�֋��G��x6b�3
e���6�'Y�1�����}�	Rg3YG�&Q�ocD���z<�#N���V��e�� ���¤�V+!�jq���җ�$�Q�d�0�m�.��--4vpʍN���F�v��c�	�F�_5��~+����x��Դ���%�ƹ�낊��F�x����)1��Hr��l�����dd�i��'�����3 ��N6���@��Y�b��%�$�-�>l��Ц�x�����$Kd�\K�Ng"��C�J�u��$k�C$I�:S��S�$�й������6��"H�� #��q�=� ؽHI���K����~^�%����-�֕��M�q�0���v����T��"̒"������k�U	�pgX;���`���	z�P�?��K�a-K���z��Q,m�8*�25���.�(�Y!�����#*X:��+REh�	�:�2��&F:م��g�����pm��"�k���O�
�5��w���))7���WQ�����	� ��o\-�Vd�.]�o�ms�dH~�/\��/�M�c"A�|2П�m��!�m���ĸ�5����:��>����8hZ9�n���>j ��P' xL��C�= NN��'������	�,\jG�ğ�bK
-:����,�#��h����v������G1�Ή8*�R44��m�E�/�(��yx����C�o�i�,�[���LU��jQ�^����_y����?h��>��Zu���͞H��P ֔�i�2��Ξ�CL�t����U�ҙ	��*H�ɢ����9�J�� ���+2�L>�����PBD��tPs������MF�|�fo�h}�.O�3�Ǽ�.¸ �설:_�h%\�Bi��boQ�Mu�S�J���[��ӆ"&��PW]i�,)�Y��	-�4�M.}U �^�����;񁸭����s���>͕bq�x���芝�$	:��i+�C4l"�e�?���2}��@7	-j
w"Z�\X�/~wU[�aϢ�:v^�e�^���D�9��l�fd��g��0�.���E-\���ӑA*Q6���'�)@C��H�3������� ��#�u���?7���H�@FD[�?�϶T���k��ȳTU�����K�)��:k3g�»=����s9]6�N]�y�Kj�o�( N�8<Y ��?fT��1lSz��2��LF"`:����1���_��\8��[�u��IE(��P���E� �f�t�bU;;cU� `�mj\��X�3�栎JxC���	��+��z�n<S�N`UDk�� isY���%:u��AE���ɝ����Y�P��H�H���
�	܍~�4my�_�s�:����n��4�F�5��~���-B�"�'��b����1�?Ҳ'p����G�K�� .��B4��g�c$[iu����Of��?��]Qı�d��x���Ap�gy��V?Ն�馒M:MEq1ь}z�j���)��O�H*�3��4b��C�E22����X�J�E��L������ⳝi�4�-�c��3eT�_��G��sQr|�)��y��;�Ɉ�-\����,�u=�t#ۏ���ٓ�&��r�T{T�s�n�����9H�P���Ũ����!W�Pg.#�u�rP�Oݵ��#c�k¬�fR�OC��rGr^�ǟ۝���󔓵/V �:�d��G
}��~��c��O}�2U��Gkc϶�ͰVMT�9�	M�6�)<BS�Ύ�D�4�{�B��Jc���9�{��Җh$B�jSن�Q�2�S*7g�hw����ah|��f��kZ���6�4:�ʊ��z�<54j��\��6�7�ͷr�g�,ӱ���?)�yw+��pH}L&�AC�T��/�/D��"-:Qd�F~�@�V�?�a��Nɐq��N��2:���d���C�vf�����Xz����i��U�����wW1��P����Q})�l�	9Z�SF0�4x��W�(c��e ��F\�)�+��D�% ��e��U�%�	���L���g���2#���]�VC�h�~[	�T��y��,��Ŗ=B�|J}��6� �t�ӗ�O
�EǸK=eϮ�K��:8;zc�7�.��ry� �< W��0��psUq�@_R�%5��}\���*��{��o���������Ny����d�%j�U'	n�J��Vď��P ܹ ����W���6l���CY��;��f��c,���n�`�CKi�dQ���Av�K��(r9�������`<!�|b.�6�g�M`�ƥ���o�#�^C��DO�z��Ǘ�ۓY-!��M��.mX�հ�^���ݵ���#��N Γ
U+���ɹ�RlDCɨ�:m
�x�m�8�]L1���Ae�H��-A���!N���u���!���@&E�Y�)�)��I�|��|尹;�%}b���[C��됹���3��C�z@l�$����w��sRAC[����/F�L��Q?�s���)��R�0APb�۶L˙6򹓁�Sg�4��}�r�~AFNa�����r:��g����Ȩ��"+$c !�0P�^��8���"��k>�G����+~��u/��9����)�!�D��6�0:�%�0�߱%i�VVUI?��?�'�T���@#*�Rhh'�`0�:��+zb���ϣk��t�v�+`O��bg�����4�9��ۯ��U���#6"Gm�݃#ב��o)6�A�ל�xֺ �|Y0�2���$�sZ:����B͓`��n�s�5�;c+ᄍx�������K��+�ip���67�����$>�uU	����ԍ���Wu�ͺ��b����B�d��D�$�A�~M;��)�ǺR)7� &|������ϗ�ʆ���n��xz��]����2��#��)���`7�5`@����D�dXc� ��L��&�w�ZoΙ�9"8�N* �*X0���%ŉ8���3 �a$��o3�k�����I].��D9�u���%N �$�h�po�w��?h�)�K-Cq�_B~��
�|��X��)�c��e�����m���U��]CH�
��_�Pw��+�=-6e��=����o�@����a���B-�m���NU)����7b�<��=��܉ ��G�Yp�.F���8�"6b����۴2a]&�
��/o9�z���J�/J, 6,cX�#�5]~{	 q�i�/��T�ϗNz������0t��`�~������)��. r&�J��{�a��0n?�2,s ��\�&���W���yF�&7{� mn5��(�y=;�b���NA�ٷ�ƥ�{�6�Ԭ��])���()����
,��}9w"��6���AFIQOm}�-;�����RoT�l���"�
@;�D&-�m(谖 ��|4]�??㿁���J��8L)kɜ�S���V ]��h���*7��b�a���yZV�ˍ�ͫ�qg��"IC�a�b[ͭ�먪3��S�ȉ�!�"����\p�h��{ov�g��$�D����k��z����Ɇ�;Do3����
��o�7\(�&���Y��(�i��wt�\�"g�@�R�nx�
 �k������co�4�hꝧU�#nw�`�¢�A�C�.��H�>��P�{���� �R{a��4�В������Z���f�m�C�i��(�V��B�B�/�l�pk�Q��-kHO	i\��w�7Y�ʘrv�W���2��2�/V�i��� ���`�2��m�_C�����B���!����֐���!�����+s��sT'f�,8�z��O����2N�ҿE��}8�G8V��FA�&��a�!�=#�J�ѧXҔ`��%g�7�%r�<�n^�H�+�)'N6K����s�k�'ʰ�V5�O�n�Ή�h�;v�N�?��EH��i�;�_�e">у[Hc�|�R��oY�Bz���XV�0� od���b�x7͍7��jY��*o�`��=�n��E8�}��3��$�'(����sy���QJV� dȲ׿�}"�B�ɘ`\mիʲ���&�=
F�r5���.�`U�*���$ȉ�zeh��3��c (q"��8�oz�td�)E�*T�U/4�jo�U���@G�.6��[$�qc� �Z��]��d��G����A6R�K �$���G��8ؚ�fqق�n�S�ْw���%�Z�
n� R���+7�v�����}�G�
L�~�<e%�v*V�KR�*��Ͽ\�5�#z�q����3Q�.��I��)�U��wr^=P��+�ˌ��AHlc���<�L'���?��ط�@8��t��6��#��e��r��hh0)����O�^|M�Ț%l�6�}K ��6�'Zl��3JAv��熘W_ �M7`0��)��lc�دr�p�Td��$�k�,4f�|�cC��=��W=ZU�m.5�ϥ�6�PZ�
��$5���>o6��&�|�Uc �|3���<OC ��5���墱kQ��OΒۊvL6.�թ�x�:�ǧՋ�%	C
H���
n?+��3�n��
 �X����~=��Z��V�lK:��K��\7�fOf��/ŕ�6g*�<7����	�K�����%���o�%n���h_VV�����Y�y�$8�����:}�.�g�<b��[@��bZfC��w�d�U�!�B�� �,���g��B���Iշ�Mz�ĕ7��]��Z�2�&�?t�f-��z�􂐞�'�:������@K�;� ܘ��������]��|�-��xNy{4�v-�a��y�����ND�4�V۝�;ˡfh2eg{T�ING��IG���) ��zw"3������U<(cH����Q<v7��ܤ,˄c���3��F��;�o�O�\n�̀�jD�YamP�-��!��kg�b\�"$p_>��(T E�{�p��@�_Mh���0�����xg��c�:�s���ؾ��W�B��K2�A��َ�G{-�c�ք.#�P���+B�3���o�;��\��A��`��$W�q��a�ZO��?u���3�=���rRzo>�E��tf|��t	`4:�I>�$����Mk��a���w2�yd�#BR��,=@��<�U���x�v�h�y^1_��38n6��=�X����M��SPkJ�s�l ��l��k�WW��&U��ghi1��C��pm~	s�m�R���Y;�G�`�(��\ˀt�Z��!��Vy�m�+АpJ�m����=2oi@MZ�h7�=ѝ�!�)ƚI����)XT��
Y�<� ����$�5K9���ͭ5,r��6𝤧"���������㕹�!fE��"�Łr3�)h��/\�R����$�z|C��z������Q��DHYP\@B�֐�7���h�8v����M�Hb
0f�ӟ�qx���ϵq\�IO����j�ˁ-�XVq$"Ҍ!u��i�J�D�"�uИlp{�a�����gq�:�ZU\��.�#S!�/x��S��P�0υT3A��Ϭ�x��O:�X���jh� A/��mkOĄ��hh ҠpD%��I�V����o�u͝�{��u"�M��[��Wz����X_����0,kִ���S
eK;S�< |�:+Z���Zԧn���Y�΋�mIB,�?����+���Z7��ұ����W�F��2�n���#[��x��B	 �9J.�N�V D=�7A94Nb�;��a$�0��lL���WHi�Dd��	�7����J�@��Q�W��/$<r3�t}����,��ǲS�"���I�� ��J���)`f:�������\8��ac ���u�G�ni��/�M��f��-R�Q��,���$��uHW.o��?�k$;�1<�=�2���M4�X�C&z2C�v�JiZ���r�)�}#s/,D9�6��N���mZ�[df�V�>{eK������Ts}��S������ٕ�������������<��l�:f[��@����+��)*��b6�m��p��l�;y6~�l�B�*6��.����2��-LcU �y+�A o�v+���ݽ�]�.��X+%�g�ʨZ�ڞI��q���	6Ƭ��I���]��G G�k��!Tu�Ə�� ��υ穘Q1@� �-��mE~mXt�d���
���zdf�)U��V�Ic	w�x�%�C+W:V�
2�L���`��2�/m���\�2���R�Wby1�P�7�9ހ��if_��UB:(Aq����o��"d�.���&8�<�V~.'�å��LT,���� ���驣�Ӑeڱc�Do�Fa��|��u'��'	��
��W���m5��+|�Eg~��_�r�����7����m�3��C�E��ݩ���Dfy��Eԟc]k�Vt�B�Iy��Y��<�Vk�Dj/�"į�X	��l�.�&#F�>�eE�d�2�s�tr�p��v�8��	�,�T��@2 _y>
�D����"r*'w��6�Z��|]��v���f�h��s�b�����?x�hF(݉WeF�>�'p+ٷ_����*��u;<8᭶	I�V�-*#���Dn�A2Ӭ,��FN�.=���b"���SD�}4�1��
�����8gS���h�6�FB�>LڬW(:SG춽e{p>�j;�8���:�S��l�D�m��O4���^�6"i�,G�GԊS�F�* N��Ż�ƚ�۳�"O��y�יg�JU�'����S�{������
{8,����	�u>�蠄���4�i�!~��(#ZJ�8���#f����DQd��ԡl�����	c���M�R���1H��v���\T�%e���!�2w}+���)�	���6˘"/��neY)e	�d$Y�>��O�_I�'kx/֛��?���UN+�.b@�m$n�r;it����j�S�b��޷e���;��C�����!5D%u3�n �6&����Ip�ʄ��v���Z���,Ys�O������$�vHC��c_|�l5��қ��H�O�<� Vƫ���-��� [�`3d>� V,3��v}z'�^-jJ�f;����O�� �����fR;n�C�p�N��'T���J�Cʬe�l��w��߯�{_��x]F�)[8::nk�����Ky����0{��p�XM�:��n�c�ܫ�n������⠜�����#Ok'�lx�� ��MWr��B�����ǽ���}�Fۈ҆�W�sM҉��L�D2���K#<e.r����@��@Xl�����y��Dk�=��u8UxLn�	�է^���jU� �"��\yo]6�F�������K�Ց�+��E���4댟��� t�\����L�B�ϖ��S��~�=����$�
�D������	鱂�����xH���?V�o�v����h��iw��0�A�0�L��_��So��:�O y��h%��M~aɧ��D��ψr�Ϥ� ��㨊���60b��G���&�wj�&\��P�n�8�ν9(�Y���s|K��u����[!a\�D_��	k؝�6�
��x�W�baY8�t�����3��!�cc��M�[|��_���ү�L[�u���J���Dn�m)��L%�Y��K���[�^����2,:��;8Ӵ*�L���AvD���%\eq�7����$ZM�M��i2��{����mT�;Ը�lD��L��Բ*��;x���eD�+ŕ_q��n�m�K��U��$��^�ј~J(�g�����2�p#vV��'�ʡ�m!�K����\k�����T��.'�����.'���wz��륦.oI%��8��������|�υ���!�CV�M�C��6'a�P��Tk���={9�US�u]ZJ�ƷqsN�P�� B��7�#j�煿k����n��!�"'���*u|�!��v����}�p��"��ْϭ0��A�����0UE���Je�<5�֎����[�c��ܛ�o��C��S&���,ݗ:K`��Q�E^yS�~���zpԪ�\9���噝<Wf��TԄV��:)��6b��!N�X�L�Ae�J�#�z��&���I����ߐ�{�_e-M��q��.��V�U�o���>���f��Hl�����:���C�l��k�$�R��I��)5�X��TEY�`R��V�{�
�j����ϳ?�� ��u����$���*�V���d��7W��'��h�=�؇	�7G$0˫݅�(M�J��k��Z�h=m��I�Y/E��.ۇ�L����b>_1U`c~S��N�;eEI8P����.��z���f3/���!���i	V3T�fN!��j���Wܥ¢)s&�oi�ɱ���]���H+��H���,	�,HB)Y����Ќ�S�U�\���	��t��5��Ź�2������j�����Kέ��1�cz���<Ӑ���A���-�(�ķ<�J?��/?^�|ōW�Tf蒕?qf5�ᥖ�i�%k���K͐�r�b�k���J�Z���Ҟ>���$��(O��	��B�6�{E�m����^���F���`d��W���/����{#�gO�kG�d�Z�ф��W�1�|�׼���:U�l��
N�>/�%mԽ��y� \��2�r�}'Ȕ��yܺ�n/T�ؚ��*ҥ&@��Cpj$8ķ����2�}���hP��zȜ�p�`(C�T��c턱�&��I��m2�������ǻH_�"P���E
�n����!��S�edӓ�o�X5�('�AV���X�r�gG"����҅�X$�9��q�nmO�(���Uˌ �zW��;�G,k���f��DN�y*�f_��3
(Fbgg��'*n�̴`C>2ٗ?���� ���h~��LB� 8�&���U�\�v�C�
\3>_�8��Ig�� ��.���q��t����������_Fr��dL���U^:�F\"��e�ʡUK�P��PA���A���ǔ��[P1j�����[��ML~xAMYP�����<[T<qjB��
.$+A������_6Kdn��*,�w&�O?@��_~g�߼��|IQz�;`����qZc�e�\,0���nZ:ME��PwC/X����T!�,��7���&L��A�
���Wt��vUG���!DP?	��g���V��q���Z��w
C�s���Χ]����7���>U�~�v79���IԲ�e�K�T��@�?Ǻ�o�SȊ=�,b?�.@\��f?RH�og%��;0o�P.:l�<_oE@e�S'ڎ��z*{x�\0��l�[�CP��9��nb�N��J�p��+բ��Jd-L��� .qU�i%���A/���1�41r�
�0����K!��A�6X�R9�߆��8�~�Q����{iD�{�=��6����3D�ِUg`0���pOi .���]��1���}�I$Q-�W���Զ�w�$3�R�	hx�ԥ�'�kF���"���j$��Q��N�(�J3��o�7y����C��1�*,}0�7f ���S_S�Xd�v ��Y��	�����ĄeM+M��c��r�C�d����*�� �V�Rm1ؔl��=�
��(8�]�����fz����F�+�R�ݣ�;Q������u��c4�3YN��F�Ax�	�L�ә��0Mz�h�7�+>�h��H����L���W�&�e�7�W��a"�<��[^�q��thbCV^J�+Z���	��G����u�Zږ@�ض��}��#�	���a�w���ݬf��ֺ�V����s��#�u��v�����E��2#�n��Y3E��X�<'X��}W�rP&k� Q_󱶬ugcbğV��/ζ6˲
����m�l_8���{���m"�1�����k@qwѲ�BOx��~Ռ��Ĩ�-���vT�4�X<L�,�l>�3"_��s��O]*��e��?a�-?�0��&Z��oLR'�õfǃ�"��v�˵�
zt��(�eS���pI-x�9F�[�<"���%��ڃ��GYL�®0��ދ�?2y4�j��m2l��V�ǲ�WelبL�w����:c��.�Y�b�i�-U�N�0uU+���ZZ�,Bm?�-�G��T�P���� �Ǟ�Ӓ:�o�d.'�~�_[^<�LBz^��c� 2I��Ф6�>|������8v:�Wk��ߏ9�V%���Qҭ�N���Q�l3�jJj��Jz
�j7*;��lL��.��4�I�)>-V��RE�1U_�=��އ 
OB���D�6.Ɩ�],�Lg��R����-�i��i�<���)���HU�R�-e��o�8�z��46ǭo�)ias�x��يr&ªo-�R<��O�%��_焩X�G	U$��ï�16#����'�<�
M�l��b�8��(a��7�Z�!�h����L8ê�H��$-�:�^���r�k�Ԡ�?�]�5P�9k��������y���D��sߘ����3<�_�_Wce��0X��!�O+W���G�Q�9�ZS�ֿ/uE��-���P�)�s\�K�Yŀ��Y��1N��122�{��$��G!4��Y��Rl~�*w���Y�~�O��ǳ$jG��E9�~���/�W�T�Oxc�5�#�s1T����5�}��%�u*����~����EH{�9�=��f�?�,��HdHF���ߠ�hl��̓|�hּZ�qe	h�ھT7��L�6��[��\}���-�BO��l��Ҧ�{��w�_;6���(z�@�Ѩ�;<�F��QD��	e~N���JX)Hf��f�(�˾��~���@ZCW�2�d�}3i�N����5X{d���*F�0ڲCp%����-�P譓.g�����t���:73�)�R����2�o�5��U+V ��Lv�\�gl�r5X��|�N�,��؎Va������'r��7����z���lo �q['A�K��������5U�¤ٲV�
����p��"(:���7���/e���Esl1��o�4�6hw/X��c�V/��4L��.	�K(�"����((�,���w@�H
M�
�%Z
(~�����x7��.9�����=h��R�¤������^��XL�V3*%d�S3�c���	'?b,�T���g�;�!OF�)ŃK�?VVc�6�
��gt���,w�����͕s��_�8�Ეc eC]GZ�a����.?8�Ǻ�(�NPzU�D�sY�E�Ħ�-o�H���C ��i�8ܬ�Hh����N�%�36̥�c2Vvg�"���x&��E��a�7�i��2���'��GC�b��f*\��4k1��
�,�2�R=s��ѵ�?�*��mQ�������i�.u`<]O����T�s��y���mL�T�I�K+У,wUʧ.I�-l���Ӧ�ܝW89d=�x9Φ���q�6�p�;>7�!�~�r���赚�o��~7��.��iE�_�*ۓA��2xz��cwM�SI3P���XNm��0���dlG�z�1�ܥV�ʝ=3��y<K �Mk������ �r7�\��|�Ȩ4Ku_1n���O:�{�m�S�ہ�{�#��?���{,��!�N�8�!����J'�ܟ��?	�[W��b\a;���0����m���:V�m{T��U�FE���UJ�H��ڐ��n���������V��,����n��^�A<NJ|L��s�CT谭��8�݂�X�K��VkU�*뢠e6�\�gJ���:P���K�2H�`���X7R4]�i��� ��$^��v�����[ko_NiD�먏d�Cd�=��l�[w`��I���/�D�b80-��S��5�R;^��Zn�:����˨(=�K�8�Ƃ���,��͔�f3�#a-� o��y��� ��g�HN�_bNy��8�1��'g��2&gH�ߛ�U!��o�����UN�:�p�U�:��p�=�N�q�%"�����ۏ9W(�H��`��d0��T��Ѹ�!�����H}�aK#�FQ��E���݌`c�xƪ�γ����֐��$v��-��٤F�����4�.��H�P���&~���j�R7������Cky+I+��m�.p��{��@Z=k�0΃�	�-w��5̼&-7�BS�u�����uM��R���y_�|� !]��'��2��O����TՔδ��� �v�w_�5�����/���H.��\����4ֹ��KQ�������V0.y�gn���
*�H���rXc!�pތS8�K��U~Gw��i�)C�Kjš̺(�w+�u#7�ۼL݊7���v���� �mSc"��ې]=pp��B�y�ȝ/פ��C���S�1�DjU`71����[��yS��	N��㟝�����P�oz7�
׬�A�.��5���w�Pؘ����o�W]E����+���VREZ�%���A���D���`�۲e�8�)s�+Ў๝^����Y.�ls$/kC��tN�R��x��tY̌2N�(%\�B��}gǐ�F"<��pC�pkMoݲ�c��f2�8�������t>�
	�:84���è䳹]f&��M��,o@���� $�7����h�3�hYr��>�_2k5z_a�Qׯ*�c�ΤT�ES��y	1S`&�%<�U}Da8���}n����[���Œ�/�Sf���a��`#͑r.Zz�h��2�Ӫ��7��օy�	��6�1j��ء�7�yo`��i��%��� ��
Xˌ��7�3��s�]�/�'yB�X����Kl~l��#T�<�2������X��������Ñ(Ju�����%����s(�&>X U���R�]8"�l!�"���ň���Y_&�Ao<�<Ș/9�^G�3JQ��r��]�;�q��v����~&ۜ�,n`����B5C�Mh�&��t�gd�Xڀ
R\s)�a�V*	AY0ZR:W�%y�3�v���d�nvu��Q��6^�)S���	���'��B��k���c�t��6�!�!��WK&�/2�'��o=�>�,vHYਅ-[���R[���C1  gx���ރ�6$��C(p�5�7�g� ����0�m��l��v��-	Vx���V��8<���wK�^A@�6t���p��/7�ۧʞ��)je��������+_�v�'�+�w�,Z�N���n_����s�y����L�5� s��PP���:�MΠX��s�X|��⻮i9�]r�f-όbA탿��:D+U��Cq�
��Ƣ�(�K��pUJ�*�%���g�4�S�3����>�%Y�h�0.3_��|-��)G��%T�c{�	F.X%>iG��t!�V�|�[6�{�|5_*��a�Z�S"��x6UB6��˺��e��,�f�g�� W�K;�c��1+N��9t(��uo�D[�����ͦ�%Ily�i#�s��H�21���-��6�I�:��2w�qS�v�P��3t�`+�T[@����Y���Z3.T��7���.e[��-���l������c�K����!����P5
��JQ쟃�bDB7�e��sbN�X�#O�U��j5}��-c���}���OG����f��F������6��d+�j�Xق�`��D�Zq�0=��/=Ś-%}F�,�d%>�p�X7�P|B�Z�:�)��Z�����+���X_Gm�w� �4;5 �J��z���is �r���얖�Ur�k�=���?,���M�i�:˱�5�ix��gs�߶��"(�#��C!<�P3Ds+�GZ�o0e~�^5W ���>�$SBw�МU����eq��1K%����z5�ŚB�7r���m��D���yEE��p���0�� �*��sٻb����0�ɀEb�-�/ףޝ�X q��wܩ�_}�{�z��\3�"$'�}ƲɗV$G�4��$=׼=>wh��Z�2ߦ��^�N7�(���%]�<�ڴl]ܾK��G�_[��Z�瑫<���GS!�V!�m��q�ؓ�ss���`Xu4��u��з��>^ľ�r���+آp6�	�`<��n�C"Đ�_�����y'��7�P^@�9>m�d��KPGLvK��LG?ݷZ�\_[/�ZA|�ѣ�����9#n7X�Cl+Θ�� ��4{�j�O~��L ��*�ev����QP�P�� c*�F�7�{!�=���� +Oɮ�Fb��7/L���] �"8�`�AKS���=9��}����k���57���"�]�#En>@���%�O~|��g�1��������LC��h����`Y�=�f�l�� A�)��զ�v;�@{�X0��NZQ$�d5�ݮ4~e�U����BIw�C�;��~�z7�:�%h��Ll9�����T,U΄�U{�nb���v"���2-E�g����b~�o��P��#b�XԽW�J��v?��7y%׸�e��ʃn�����Â&$�! �Olb� y�7GYg��ܝ�*!��q�R�?H�Dz �K�|��"b�pL� ł��!:��Z/�\���5�L�H`��ZS���b��]	8�]��brQZ'��'oGBڦ��;�$�Ҷ�[u���x�:��-�δ0�"O�	G�;��A7T������*5xP�= ��1�_����e>;L���U�+���׃d��d���	����c��5g�xʛh��1�1~KoraGA�р���l�'���'J�6^C��a=ɞ��{���R�*v��E`Js��,J/�b|�v|����7h>� ͆��4�&�6��=�}�z<�1 'n��7�Ǐ�w�l����sY�1]bIa�s7a.��~e��}ŢΚ�
�gc2����s�gg����p��A|ufI�iLs����ߨ��RM�*��,'���y�Q�)5E��DD��T�c�R�e��S�';J�7�Ϝ��V��2�㙗�3�#�Ʊ�yJ"�����=���Y����Ds6[k*����Y��>���i��,F�հ*�&I�Ъ}��\�'@ZO'}���s�ƫ:	�%L������vTK�������t�a|*2Z]���k��:���߂��i�_���If#�ޤM���`΢���Gc1�ͤa{�!;�k3bΫl���=(x[z4�QF.�t�2�*��|�øy4[��6k���غ�kM_
6T�G4������jX��2�ˈ���k\�iܮ�Q� ��d�b�ה/䤒Y$
����������P�R'~Wk���X�����%w2=ӄ�{%*�������C1�-��L3�Hh�l�.8%o+��?s.�'b��ӊIP=�^/V�c.�+�&��ɭ�2w�oH�X�u>�N���y����\��;pF�����C�&+էIk��H�Ϝ֞�"%�"���7;x*���k��/�m�Hl����2��q�0� �p2�Į���S�V"�",�1ɜ�6�=�8ϧ):5~D��B)H�п|¶����y#y�X��BZ�JOC��ʵ��$�bI?��?�Ӆ�*y޿x�O���s�z�֘4�9s�/�X�3��"h�R�)�qo��n��l7�y|�zH\�UHyq���ݗ���D�`�k���j�$/�ߙg�q}1��l+.�8�۽�*�������n��4��?�A��OR�̧�Ҟo ��߲�A6�6��˵�>����_ �R���5�֜�&��t�,W|Y�r�u����2��*|�T�����.�^oX�9�M�������-ND���/N-72��D���񱚿�b:��(�G'`#3#7}ل���x/�
,C-��'�!t
(��ʽ'@?����A79�,��n�|Ť�
�;Bn���Ŷ��9�}7��}�bW=_^5M��R��۲�-��K��l�P��+�x̵��� )
�QE�D>E�,)6���>�&J�j�dGء3;����c�&p��õ�H�:h�zb�.� ��ʺ=)o_�)�=>�ߴ�;03���+��`p��](���L�d�O�
'��H�&s��P��k�����Z�D3����6�Ga� ���y��M�v���*�N��)��q�x0�@�`���N�J�)�D*��jA@�fU�=��h��E�����0��H=�7$?ː�juo�Q$���y�R�����̘�d� �2$e�R�i(�ڽΡ��ļ�8y^JJz��싪�a�mT1�%�!�	W~�\L��2/fK�* <��W��!j �qB����)z"H�j��{�i-L�z�5t�\P)�t>nŀO�7�w���+֔H�D��6���а4(�Rg�P� �4�M&�@:I��"�Zh�@
�=yW_"�	������#����AiR�1}fk�� MUN��*��dx��� 7��Y.�����.��Q~u��ar��f0 �����3=��q��`��*w�
��'�1��8��fݷ� �p���uRG	�����a�C��摾�T�O�*ݮ%�KQ�G�n��̟��y�C+� �:�4����X�Dˈ�[1�J?����e�����*TRp�!��`����:�P4WgmX�K�����AHd�i6�o���":?�Ou��
�-�}�j�
Gqvt�sa����h<k'j#R��)���׍�p� ֎�(����4�N~
U��K��Rq�`H����+����x�w���v����rm�F(�u��!票��.fd�h[�&���O��6�L�&?�ޮa���x�n;��E����%І�m�4xs��n�EY������8<F�	�3�wT���<U{�%r3����'��fQs�I;Ϣ�Cq��~ H������)�os/N��pV���MT#�;ʻ>ni��.���v�T��e,nô���r�����V�o{�qٶ5���U �$�쪀�kv���|��VNO�S:�B���)u��On0���b���6۶�u������Wn�cö�`�N���eP�3ؙu��|�3u��G���4|m�Ǫ�#�e�?G%����TL�C�r��nA��ׅ�KP�jcE�n�	w2S:Q�N����>�?w!IW",�H��o�)[�xwS(�qv�z���:;��p�NYX�T��JD?!���� }�=��iL����`���Zl=|1�,R�<ʝe�	�~�\e*O�n�D7]�/($�ˡ���e�O䊫���3��J�e�:y9;k��Kt�L��Qe&�x�gq��}KG	��VR��83rw��s�����o�����Ds�����W��I�s����,�h`�v�@3�er����X��@9��,�q)��������7 ��X�
d�
���Wi闭�����i��d�}��4��C:l���U��.�$�w���cU-�w
ߊ"BO%}��'�W~��֨�%1Ԕ |�9���l΄�?2Mm0$��Ki q�<�o�&�?I��\&^��Q����i�.,�J
������}}�ͧ��&4ّ��ӫ�xl�ٍb^������,c?.���'?3��_F�-Y+M�%��!f�8�T�\(;5��&c����N>�����{7}/�bŜƶ��Zb���i�3`RE�]iUu֦-��<]4�������M3�o�꼤��	��S�C�lS�T�zf���iH5�`h��؍M�i�@O���.^J�׷0`?@7��M�����-�b�hK���cNx�!������&f���4���� ��sn4�R<�������z3sœ(���~P����ԧ��#�Η�4H�f�a���� s%4n�H)0_T�o�q�����F��j9��s�7��5� p�`x�9�p��`������_�� ���]"7��\A:p�C���ީ���p�o
���*�����z<����[BF"�le�0\Ǹ�շ�@�>)��*�⳧J�ظ��m�Z�/�oD�Ɲ��zm�(ݴ�h��0< %eg��_N���ݚ�b��.���0=r*��`�>�F�7�����r�"�{�lͲlN</8'�������e>#�dX*�*Hp.�RrOr3&���J���\�x�}_T�ѷ�~t�M��l��Dնc>��gAm�K������:?����-�4�����[��'����`ꏖ�d�Ŝ��ӯ��f���5���zr���Xw�x/�3p�W��ݺt���Ep����������VdBhǳ��ު_��8U�WS����� j�`�JV^����#1J�Ѽ��u[���+I(���b�F�)b�v�II��P�߶��pb�q��D� �:��U�v�z3-��,oj�����+��^�	�_Ixj���7֧���j4�KY��N��Ǻ���W?9�3&#��hΞ�\�(�~�<�fR�{ƭ�j��2b�����~��'8`���'OQ^d�`q~��˦wL���!)I^СE7��v��j믘1q�i�3��!]��ެ�}�>�o�o�����	D����Z�*a�� �"�\Y���T0�l�	�h'�8�L���SUzRL�fY��I�,*ۑP�^@������zF�u�L {��W�m����`A93���*�9t`����C^���m�� v3��Pq	�1��£��`&�V}E�_/Ф��"fne5�o�@\ne�����d)"h��M��AŖ�����W��z;�{�=C��F<h*����-�!���bl�gy��IhӅ���|U+r��Ψ;���:!��mz�u�ġ:�W�����*"��pw"�������&t�qZ'u��V4x|O�� RǗ�*B
��L�Z�i(rݿr����`��T	Bty3��Z�8���Ԃ�ڙ��j�
�$ZF��S��~f���$J��*hD�:�7E�ǯw�b�(1H�m������y��]�p���������u�1����V�{H=���*�������/n���Дbn{����2K$��YP�-Ґ{�-?��L��<v�|,��r���ћV'�*��/a��7���4#�N�胣9t�A��#�_�ݢ�����şS�P�eI�����D�	x��~ϧW���{Iܹ��S���)�����p�j�7ԥ��î�_�G�K�'�B��6 ��6|i��C��؟���b{���tEq�����"��9��R3�B
BҬ����BJ�ĵ���zC['��L��Lt7L-�F���N�5����i�$�|���r⏄`�.L����_2k��o�;�>��1zA5�m�Ǻ�YI�+H��3���7��J;���&��F(Gw�� ��tr�?��� ��Ev��Cv������:�#�S�N�1�o��,����WGe�ԉv��O<����zK�b�w=�D�C'��װ~i��_f�&��<��X� �w�]��u!�b�}C�G�͂-�?��\�P��1Gn@jڿ�=�[`y�XU}��=�X�>q#~�g@TL꠺Аq�z�/���������[�[�aO�G��V�˿�/�q��%�ث��
.�cP�����eU�+%�/��̡s`�p����G�'��y����uF51:ă�3��mWײ��8G;�@M>��R3� ��N
�0˓�2�x�I�����=�.߲~0\��Y��s�J&������P�C��d�f�u��0�>K-�f�VFji�1 ��t+�������+?�~�{5�֛�9�w�W^�!ӛ%�:�У���}�ٯf�_'�U�s���_=ѯ@u��:�a��ɱ�5�:h�a�Kd����$q�ql>������]XN�<�o����0�I	�sp<iy�Ҁ�g����������!N�V%VOjʭ>G�F����(�֍VY�MB��[��l�%p%5`��$����Qӑ�LSʆn[�8|j��c#u�.r��@C�m�g���jY0��k�M�{��f�rtw�:�g���⶚��P�TNޜr8-d�oĔ����J��؉R!�t�֒�Sz1�3֮�ڼ-BI��\޳�*�L�eN�$�R���$h�& ��7@�K8�Mg_-��q\�r�`��M�O.D �X1�˴�1���ZP�~�u�̀�anU/d<�zV���QxҖ���͇
����U��s�{,�:�fy�ږ����z6
:�̈́���o�[����b�1ق]�鬁�6��7����A�y�Cd�-W��9����Qun�]C� �\��Ĕd���X�rp�=ï ͔壅¡ ώ�+uC�]0��zl�`�`��O"m�a�� �J:`�xi��=F��+^!t��]�)��	��i�l�a��^�y�j�Gj���E�)����0g��0M���ۃGT����:`�b��gQ��_��K̺^�MQ��X�YS:����=99"��c3�
�iE��4�U_$�i�e�p[�p&Y/S��"v%���*���<��.���f����9�ښ�@��#¡�������vR����G۟�0�h}�839�[Q��&4�S��>�ٛ�S���`>χ<��n4�vq��s��>�&�I��͢�q��f��a囎Kw���QW�+�DX*qL�/D�;(ǧ���7�7�T���� ~A�Eq�+n)�����|/�c��;}
����=�r �Xi�-�����.7�ZZ��VZ������*v�ޤ�Ms��9%��9���n�^-<�K�����UsOrM��Ŋ5��P�o�a�U5z-�Y+A������EJ8m�2�d�����q��*��i*)��a��I�GK���6����P��Y���m<��u^��,��3>&�2<�ײ�I�s��_AB��Mf)	�X���i������ � @������gv� �:]�Q�󡑑�ʀ;>�;��b,p�B��A,�lۑ��^g�C��v�70��K]�2r z�
���6��oÓ/�Y�"�ƇG�3�0��Y\�3��s�9�>�C k�����X4�H�'�v�v�� �0>B
g�GY��;۱
�,$ۉ<٥������6����� ?�6�E���%�ͮ��9=�*�w�<���.���,Ԁ���ۍ�j��,���Ϟ�p���P�oy5[r�n��z�'�I��b=&Rd��K�1On���B�Tjڛ^(-�ӫ8����yJ�鴩����e���f}*q}t_�,M׍t��z�S�M�hA�h�7WԊ��ۓ�LP-��!H%5�A?�rM� ^
>�� �����o	_���	煮�_u��(f*,���4,��kw(�U�|�#]�j,e�������ga��&֬ʊ�x�t�4\D٬K6"�Sz��.FjS���RH�>_8�=]*ꌥ��]�M���G����Lq��XI�wbq�������=1W+��ӎ�-�S�Z3*����G�.�s�����h��K�����ًL��FL��G����E��mc5��!VFq82�uj�䎇���=�!��Mi���F���ؒ^8���]�;������t��@�o<B$��`��<�]�<*&�#�Y5qVXz�l�*�	��>��|&H	�i�,nl����.�x����;;�1��g,ؖD�/�ٲV
��u<�A9�c�g_�~�@�u�2����U�4��:�;��gEǂ�������6��O�`u��z�q�0����C2�]X���W��ȹ�$u#fUE��̇<�Vi8z�I�XS؀����`���&�����W�eO��8�a������ދ��dR3�JB�tE��~��}�UϼP!I6���5���)�PթM�I}~k�\��w,��hC������V��p#[��hR���s+e|U��@��'J�A�8Y�߷1����g�vt3cOf���_���=H�L��ʄ���&����@�]0�^�>��#w#��V�f'��l�f�_�������7��'�
F|���b<�wD�/�AV������%֖#�!���Z<��9wM�������:���>���X����-߱��L
l��6����F��,=V��k= پw\&*�8GТ�zr<K�d���xp��B��V><���˵}r�)�X���)�6�Lo�:2y��a���֧��v,�� ���,�	�]1�o�J�$��>���|��	k��zN<�	����] k�c*	.�x��U
r����I�sa	Z?4��/e�1�s����kh`#d�sV/`��l��+o�(k�9#�k��[F�(�OM��|..%y>��gP,q�n���="�������ե0�#6:T�{��C(c���%���͐����>ݤ@��BT�"���#]{�����2��%��$���{;	�\��e�B�6��U�z��G��3�0��:x�U����[��W�dۢT`�#�<M��Ƶ/d�$�������%Q��? $BヘQ��W.G�[f$c�{J�*A�����!P���ɻ/}L5:�b�q�`p�ʘ���"j���_W� K�I5S��D����&^Ɲ�у�2�n�R�/�o�j����s��n��؊%����C̱�̄�����SqY]|.�����r����eK���z�z�f�ա��LZ�E]NdY�mQ��|��3q��܍W$�c���X��-?��9�[1��s�����r�I���_.SѬ7yܙY�z�1��E���9��FW<��m�,n)�u��s+�֢�LơI����%Q�t�l���������D����5/�?�Z�(VW���RE�/�t.&�+���dȢ~,'��{E�@�MʬG� )���!�j����O�=�
)1I�>/�vvLC���ku;�����#z���V5� ̵��Sis�7T�&�_W��Y�鑮���+LCX @�x���4�Q���h9�ӡ4�h������M��#�����f�����`T�����0k�3"����VJ��,�)�\�lg�����P3��~\���'f�Ѱ�K� �������t�<B����?Mv3��M�Y�%+h{��@؉��i�tNV�'�i�a��)Zq��z���ș1�8hA{�k�d,����V��MP�)gHJ���"��B�lx[�%_@��[��>)V@��[`�!�%6����0����vV�A��3��,�C�3��[r�p��S��x2x��z�:�2�L��%�.e��J)0�j2�I^��,�=2Nu:,��h����`8����>Ls�.��o�8�X�t��W��wPdg�f0�<�v ^�a�׽�L�;���Y�j��b���PI�(���I��YиEe蓒Ⱦz2����#�?"}:c
;k]�F�P{y�+�G?�DpKS�Ӑ���穡�/;�	]�a�z�@�狿X���֣�VSPE�$���HQ`�GWH�Q�T�s��e q��e���s�uKq�zd'4��֣�ôm���NE�lf#�t~����'��F�7z�`��%/x%����#�7���X}�A+����B>�BL�w�a��4�� /�;�|��AX��@�T��N�|����ə���tv_g~���T�yz��
�z��M��G�����k��%���·G:���]v� _�$|Y�����Y�OF��D�ʃ����w��D7�Cy<C���i:[���^;���$���LD��a�ٸi햞F�)�TJ��O-;�ޫS��!��yJ0t=2�Gdv �\#�OwY��gD�5J^_��o {r��I��b�8�4�j��$�h)�]�8�ǘ��&�V�%?|1�lOE`~2q�[�[b���~��}"9��[�m:�S3�р�t�Z�x�� �`���j���[o2�j���B����
ҁEw�����by{id�7G�]�녈?�b*'� ��v�t^��\WyǓ�#�b~�kE2?�����������Z�q��O�@�<���
(��	V��픟P�a�K�_ݶ�,���=��(Xb�=���h�r�A�)�v�⩪|�o��N��뢖F�^����Z�Q5����i���U�h��5-����5𽎣�F05��G���g��}Ar1�|��C�)�x�Ǩ�>Z�b�-Y��J%�^Ll�����[�m~vIAd9��tF;K[ qP��C� �;-��q�I�s+��Qd�>@H7�μ��cJ]����'� c���5��iQ�q|�l[�!뉣uY$x�u�?x	���F�6�ܺQ�>.4C�XC-��� [Rm�;�F)�v�&xZ�*|Q�[��sZ*$/��ԭR��1�N�W�i�����V؜�#�5�ÛO�8���t]A0֛熝����֕
jp�4f�u� qӋ�/�>'{�}��`Xj�G�_°�!S�Q�.��KY[��L1�����v��W^�^�dAM+��pE��I�!ڌ	}S��]nyG������M��M4;H�(} i i3���'BM�4UhOXߞ���e L��1�$�.-觃�(w�>d
����(�W���`T�,���!��s\b^��j��
���W{E�?�M)8�D�9�bH)�VX
�� �C�z>���m����bӭ�б  ��F[�#lѻ���b�sĭ��6	�u�d�
9�i�v��Ͽ�^���*=k�e#��������Z��T�{ P�.���|���0tT~�p���8��*��F�Ssc��y�o�O>k�<�"���Y�\=�@�Xw�U�@��#g��%�r�?����G}
�f�đN��I��tb�M��3�ƅ��"$)��U�K'��ph}��1i�G���)�����D`�&�?/N����i� �dgJ�.-����5�}��4�ex	��7\�b�oҗA8=��&,L^�������D{d�Od��c�?n�H3CF�b����2X#]
�/6��O���K˄��A�:~E����c ����ɘ�������9�k�?�|����VH�)s'���,{�|��GZ	]i�.�S�s�'f^*�����䪭��vJ�',����~�:�=�X�gV��+	)��֜�>#H墒��m̽����Ԥ�u�:L�_C �q�1��!͊�@��`_�'!�����v�t�s�Blw�Oِ�e�Z͑��Ӕ��$!�*��:m�h�o��^8+�D��3��&�_#ad8�z5Nd���T��v�����E�����x0m�2	*����Ho=mr�C,����^s������8r�hɝ^��ek�����h~��f�%��կ��d�Z
e�i�%%�}|��6q]\J%�	d+Yx3���|E��Pݴjc��u�9B�_7���:��
eZ�E�l���B����e�Q*�q8ʫ����WΛ{���O�w'O@�T�+��CH�f2ޡ�����w概	f�?7-VԔU�d]C�14��t0 K�-��f��u��0
�y��,��֜*�ϓ�pQʸD(-��v��H�(m��Tgcgi�+j�_��G��gxP��p"�DS
��>�x�"���m��S]�YF���(�Z$ iOE3����O�V꙱�w�vC�3"�Z\�)5�E3~�E��dM���I���p���|̌��E����#e�
��V�b�����9�b��5�T��82eLaIg�a[=ߐ��ߝ,7|��)6C@��z��~�'���H�VUK�ޖ�o�S���er�imޞ�u���}���0q��xL��L�N�_�` 2:�JPc!@=n��5x�y�����*�.%-�?I �2z��ǐ�۸y�.�H�w��Zp��';gC�Cu� ��N�/��je����"})n�j{���tǔx	Q�pp�����p��q\Ƣ�*��!'A��s�>-�H���d��U�N�&���fa�	E�!�F�F���X=�4�29�狰�b�31�E�.�U���pB$��1e��#��NIo}���x:c��z���[twqkN8�P���K���0J@�?��3-{~�,�p3�n|t�b�a�T���g�(���ƍ|@KQ��������M��y���.$�ރ|2�m����ܕl��0���=��� :��KtdrI������~?�dVW��o���r'��X#�/~������>/�f�RJ������?��v*��#�!�� ��Ҳ�7=����6p��m���n�N����Aخ�vƣt�(��Cr���7�)r��qES+���W��%@KP��@*�����eIG�y�R�n��=�q�B_4(�}O닮�u.���EDfN\�f<�nw;>���&?�L?:�۞�����b��R�A&({>̣ȍä��"wM߃�0���� ��E��B`���.��ў��p����,2��7��4Γ>��+������k7(�!z>�c�/��"�&o���켥V��f��Z��U��k�0�
��R?nmQ���&��k�����_��4�xr�:�����]zq�\P�q�**�E�DmZ7�7%���e�z� ��Lɨ�.Dc���7x�v�"���~u+Ȋb��B���?��9`V�.��u0��DV�^_�T!oMX� ���L�5�u���+:�R�#��ڿ檡b�ZV���\�2����9�
��#F�_&jG�H��5��5���*�*H����=M���\�6gڂ�\��)f]�qU�Lʅ�#<��*��C�2y���A�n1�&��j{A��W��j�d�f��#�q>;՝'���b����I�zI%p�J�
/�VZ��f@���A�<��مCFU����
���	
jaT�-3=���������������u׉��H�?��y�8vi�Q�TN��t��µ\NtB����Tϑ���P"N�w��魱o�⎪\�䜬�4吳a��L�	\�b&�{�d�~�����Y��:Y���!��{F����˕ۘ��L�O<���\I��h��m�86V�Eڥ?���Y���2)=�wFJ9���K�"�L?u��,��q��h=�C�)�iձ�A�Sa}�_h�o�!���qb]z�uꊂ�3�ulT���S���Q����+�<��6X���+:�C��m_m�I.�wO�l�$����!��Өu*?�A9K��Ƣ����mb=�����D���3x�	��1�ֻa��L6o޶��"�`h+���Z�<k�yt�S����zn����`8ů��@��e�6Է6���$k��.�},�M��ԅ;-�L&l/��]�?����gd��rm�Ľ����,�9�n<���>:TΟ-J�o�}#�F�F��z���%l�w�dP�0I�T^��t�:�0mr����.M��ֿsK����u�8e�?��'�I:�@�H֎��n�oGV�k2�^�9YP�G�Th��.�q�W\������@5��EåF$���1x�l�텶WQ��$�w�FjZ����,	�A?���WO O�L�D��:�m��mr&��u���Y�(��y�R{�xnrH�^v�C�U��!!��cwP��b;
3��{�F��b����m�P�߄�S@H��(t|����\kT����'��B%(��z�*!LC���%��$��bIeH�$��%c���)�]]�Ljɑ��L0�����7ק[;.x�<��@��Q��G�}Dz b]�iη1R
8��*@`F�8A��D��;��(�K��wx:�s��R��Ro���|�2�y���O�؞lʛO�c�u��(]���>�瑡����d��W���C��8eX�?���>Q�]m��lb����<��)0D�eͬ��w�a*��@N�ԏsn�B��C�b3V��/ ���Jð�hPMhpWa��s��÷I}���E��\Q��H��ї�	�M���OY�ᐎD��
�;�覘B)��Ce������SӅ|+�t���2}>���2d"��2���%���4�6�z�w�3Hϋ	�U�:�8��2!D%��TP��=2#s�^���^��~C�(��S�e51	c.�D��.�+$�� #��>��?�/`�|�^�"l�I��xK�G���гV9��c+���6p���p��<��E�(�Y�ʯ�c�xzF�]����#-J��c:��VM���<r�V���<��G� ����FUZ����~�,
�A�,���H�U�,N^�l�"�_��n��P:x��M�ڻ����}"�+��_�K��G���S�����A���������^ ��e��D�O�лm�M}�<.�]�4l�z�0��޾�9�dyLR'��wW�H���Ą�Ut�ew�Z�G:K%�Le�$^��E�X��gz�d����Νk�h&V+�a�����@�F�my�ĺ�/��r꽫�����n�{�x
Nq˰�.ӷ�����̝^��7�]L�X<����5A"��@ւ! 2�+a����8�������TGk.�i�S	K��l���A��)��z��z?�"���1:3�o����8y`i���IfD�2g�qK�d��i=����
��_H�С��26-�j�PM�2���������|7=�7�==I&��!y�%�3�Y5-B}��;��%��c��R�á�' �ٲ[��t�wƚ�%�UA��������k��'M?�06�.Y�GI<}��_e�C6��;�\l�5�K/%{K�ٟ"��q��]����Ψ�dF�)��%`*�`?��|��ꢠU���?�X$$q� �[
<��;?LRW��/�����h��Ĵ,P?%�)��ޏG-�[��8K4 ��i�ӵh��J�v<��&Z�����j̭^W�3�`Y�)�)7����`v�1�g`g � �s�dz���U�{���57@���lx3�p�)�Yʕy��_(����BԪ'?��,���vZGQ)�)&T�~������a�~,�?�/�?t�.���~���˩�٫��k@�N���P(Y�!��u@2Eҿ�])��(M��Hs��v~^p�y��ڂG���3_��{~�M��[h =��|�ŋ�� ���A��2v_�7�E�bb����#W�^���0⡞b��q#n(6�b2?;˒��ҭ�ѓ��u�Y��g	/9R�G�F	�ɸ���Q�s�Z�G��=�'�!Q���hc�<o�z�R�=NxS��
���@F�}��B&�L��P����6B����ym����+Vj{��K/���Z�W#��\6���^�c�1O�����l�y��I�~�G䚵�P'l�hQ<%�*їK�c�RA����\�7W2��h�j��g!���y�U.��	0RO?��d��v:K�k��u��(/9�|��A���VF��H`$\]�$��*�*x-)B�|a��,#��1�Y�Gxn�5��+/��\Qu_t� n6�-�4�M�'%擞�kS؝��](4�|�p`y�ɚ�t)	3#/�{h�:ŋ���9��r%Xg�����#h;�H����i���<�o�3�vXQ����@��z���`pm˵�'��;�G��-	�Э�bM���Q��� i߂;��0G�
 a�^�ˈ���)����G�qLEJ�q��C�ϓG����tkP�l�ma+zz}}63��L  �_p�4�ʦ
0Ρ��Q(�G,��F����}y�\h�3�O�,�Fb	��H��	4b3ۘ�L��܊;k�]���l���'�p�XWX.�8�7zܶy^c.�xN���yGm���&�ٽF�nq�E�q`��}ǭ��߰/�ä�1�:?'������4��|���A\i�I���abv\�W� �iM|�H��\�Gg��Qt������m�|;Rio��$�E�hM`�8����[��%Fd0����)�5�� � �4J��Ɍ��<G��T)\[�A��6X���[�Ow��墐7�G��8fˎFF�z���y6ڨ�^v�*ͩ�� �Z*^,�8��ry@���T��=�)yl@��G�0���`H,_���&�R�)�A��bVԌ)�m�WDk&&QE���A���R���OF\�FMm�V�Nް� ���L��э�|<����T	ڲ���:�@x��0���9`�g�Ѓ�f�}�/�xW��u_�mT3Q��]�T��e������d�vB�!j(�,�_}�&�N�Ц~�p�����_Ƥ��=럺�i��ky448��?W�>��F��:tE}�n�o�]I���DD'�$i!6B�ۦ�&q�V̐�79���t\�"�������X�wk[�(�rD�]�iV�D���'�|m@�Ya����ՙ�}ix [�C衭�N�0���]$g��X�[}�~��=��(3� k�}��:.�����4J�=�Έ�FF(����U

���f��6�>JjцԱ��5����lL���!ϕ����Cїu���A����s�sc�x��|��*^[��6d�);�8vdf?H)�~�ir�h�x�8����'WgP��*�A S`�yIU�zwD@�<G�U��]��o�o���$K�*Y�i	��l�X[�{������M�0��?Ѽ	q{�����]��\�7۹.�l˥�ϑ��Q0�pb�
C���P�<kv�:��M�V�<��ɫH�߬�ѕ�ʔu��-w��g���Uros&A�G�A���4�D�7z�e��]�qY��D�ܦ`f�Ո��O�Ϙ5�24�٧�6O�ca�-+�[T���>�;�	�Mʋ5~��}.w�R�1�S^E_Fw~�5��g��X�c�H��Y���+�Q_>󪪛���qa���R�W	�rc;���ȍ@&X���e��t+�wM7I�~	ả��*���-�V� �FJ�[�{�ܪ���H��f��ܖl�k����\�(P���U2`_C�pVn9���6����=?��ԻV�����̈́x�>��wJߩ��W��vپ�eOٵ�u1
^�uZ����g� I
E���רw��rcH<0ԓ�p��7���Sv���ed}�2����cI �2#�4�y�I)�Ķ�J�1�#L|ךt�I�V3��>�X.s�&����L�A6yG������]����'�F !��cTy,��<y�6}4��P��frɧby�^&Q3�|`_��Sņ[�aW�~��8����q�i$����6�@����	"\�3TH�cN4.L����r��CP�Z�b�y�)i$��:�<�ݴiZ�8pE�hv��7J��uZK�^/��0�>V���=4��TH"��<�c"�1�B���o����dFe�b.M�9�����=��	�[?�]4;04.�n�%�S��;�K����W<C�����5���<)�'�B^D�����qE�Q��[5���z��>pr�R� .���j�k����<X���Sh��ڷ^#����^W�f�Zo���uF�GKe�r���ӟ�o�	HZ>�4�5�>�n�p�#��R������ytH"� N+K��'vȾ\�ɠ-&��q�z�M<�F�8��ê���XIc�G�]�^���چ�$��&�Ǒo��mUN�,s�#4��|R�]�%��� ���a �/IK��	�0F�_�a䱦Iu���9��<�#]�O�Lf�����E�7b׏�%G.i�ę_���	곜���
�-t1#{:h��L��lm��K3���3�jf"��cW����i���DQ^v��sE3���X0d@/��yyӣ��w�"��l����@�h�f	�E�n&�4d�s��0� J�(���=�s�H�?R홼.�����u6������J�S"����h����zi)�ڸǭ�{����gp�%�J>�����L����R��-#meS\U���s�؊�QIb��"0dcr�;Af1�ŏK����ݢP���?Vl���n��B�wH2h�7���d��	�s�"NIA�ס�scͿ��&��V���*��o�X��$z�z[���9��8��u��f��%��y���<f�@�^8[��tŏ���3Ve��sյ*��0����Y^�o,�=�����N�W�)q\[��H�8�i�vؒC��� �Q���754�g�!�7�Ƽ�`e�5L#8���H�E�D��lt�Ū��H�H����E2���i�]�H0�ʓ?�\�'��k���ީ���g:΄rpї����T��V�
���[��߳|��I㢭�U;fL���1��)�#Z��w�)�o����DV!�x�>��(c�jn8�\�3o�I�D]�U9%���X�8$��躐}�x��Ow<���\'�rH��\�/���+zgƖX�;αA]f�?oDS0�n�?V��h�.:�Y�G��r����DH3�+�"|~���D��*!D�`'R@Z����t�!o^�n4&?���	���,Oᣬt��X�G���m���+46#�W	1�����
c^.�N��&b��Bo垲{(��%jHL59���[S'�d��jv�x~f��n�i�������U�m"�A��M���(���@�����ν&^�~]���L�E4'��J܊�y�FhH�G	�l�\:W2o�e��G<�E��oy�m�+��@��R<O�!Y+�q�<?�jf�
��AƩY6��w���2��ה��ʍM� Rll>�A�e��>��M*�|�-T�5j��v�.�N�0�k�L+!�Բ���I� �GP=���MRU<��>{u���a�f'ҕz�<?�L�h����&��� $L��
��_�ؔ�M��ŤS�ؚq	T�/
�!���}�A�� �`K�sk$3ق�.	��i�sU��J���9����~3G��ns�3+�,0��9-����g��a-��м�^��Ԛ���R���;�t�����խ�ݻ8�Lگ�jЃ�z��Nil�w'�g�J�"��E�+�_��B��Q7*I!44�0����R��GT�!��_">��~3�ة���E���{�pAZ ��s�h�*J�<�3<����W�*����tUi~ !/�l�`�wp����`�m��l����n_��Q���mh����F!�r;'B�7��\D�Ð)B��O5�T_�{ό����$�c�����AN<��j$ܡ ������]�Il0��/��Y�I^�2+rؽ`�	Wr���#�����@(�pK9��ь�h{�J��ޠm�u7���9T�})��U�d �؁��zg�u��v��~�}����K?F�ZI1�������UFko��ud�%7�w��9f���Q^�k����L(d!�jѶg&k���J=A�~���J�0�i�`v��Ġ!����9��p%w�P�֨^T�%���ɤ�*�hg5�	
��?cqG�� ��?�G���=֐	I�S��!ھe_#���q�z��	��E!��hV�g�!�P.k���r�����pA3��S��<a��b\�a�*��ɘ�-#d�ns*�Eʭ+u�s\70�o�6�cYx�7+`�F՝����&�d.>X����@���:ڒ��L��Nw�0u��h�h�{$6މ�t���y"��3���E�Knl3V-Nq�^�LgZ��N=[jTL<>`k\���_��~�����D�'��*�T��k�#gge�@����#���!�B5	q�ŕ������q|RǠ�}��s�(>�Xu��:k"q�m�f��]�/�6����M�FT���B֊��:�9�T''��,�u�j{�h��o�b$�=z�ա-�n��R�b����"�L�H��I�h�u!�q0�㹍%�F�#H����/�T��1|�/�����lV�G��-��&�>E�ﰘn�҇���b���Va��M��.�v`&�[T�$g�������E�.�C9j�\����"�S-�6�~��[j-�x!�T)&��+�LE�{�]癵�E�-����w�u^�|�C☼:��$음�C�/'q�,&�XX��Q��C.E$
��Eb��~d�_I��./���3��v���Kۚ�y���.I)��GV���3XVr�~��'݁UK�ƃ�]������^M�������k�8��r;�̃�e�%�K�B�̑yu�8��{��J�Yͯ6���������t�M�Or��wV�����m�iwvqA�A�[�?hǻ�y�B5տK;J�Ӫ'M±$���/�H��k��B�ĵA���W�xU!fwO��!ؔ��yћ���/_���d�8�E��l�0����Y�Pe� ���V>ICr���	Q��HGw���X!=O��dM�\_[\�hҴc�O8��#�f�pM~t�i1K>�B��e�
ޡ0`��;y�s��-<7��7֗\��R9�K��PT�Dؘ�P��U���,M�~SnTvӒT�k��z/$ޟ��G�+�$��$����^Ҏh��$�/[7�m��ɦ@R��+��LK)d-�I5{����H`W����*s:r���#�D�\4�R�_*!�Q��x��
A!չ�U��e����{ώ]&��;2��n�b�c@,�aJ�ۢ}�%�I8L��9&�h5�Urٽqh��s/kZ�L�H8�ț�D��B1�DZɬ.4_¾��2��N�h+� �4��p������U쒵cU��U��]H&.��{iAy���9���A6�LhK*Ǜ�ֳ��\���i�\̥����bWQ�*���X�����M�y�T˶`�n�j8�Z}�B5F6M�DZ5:h���6�n҄��|B~x�5WJZB��X�����Ԓ�F7SY}��%mlEF���������#��?�gx�����=h�HM�Qt�d�.l�;�u���g�Nn��'�ѯ�@�A�<J��ؼ�Vh%���[�V���n���W�B#}鋢���I.�P��k@ƞir������L�z"qRLB��e��A�&v�j�{.G`�{ˮ��RX�4ug��Ϧ�`:8���C����[�º�.k��뫜#:2�����槉�>�Wf��!h������{ꀮ���:�!�E��6�e�ô .]}�G�ò��O�Ys")���I!�7a�������3��c����Z\}��;[�Iݲ���Q%P�٢Z9:���@��,�k�CQ��/m�l��Լ.�������<��<��{3�2XvN�lg���ȱ��4(PH8F$y̝�K��ݚ F��g��E����}�֝��D��7B��Ne	�����9/���`,�h���-	k���N��7K��)xf�9&U�5n!�����#�Iv� 3m��&�(=�O��qQb�$K���

Q�mlYX&��0%�t_��|�4�)
 ��д�(!n3 �ZI��� X��%�������7a��6e3#�7w��</B����$����r��}-��I�(c�N��$!)aI�D�rWf X1ȆE2)Z���H�?��s5�6 �f�s����1�w���a~�st*�u;q�Q��CX]��~m%��h����)+���}x�'�͸��\5�B���
��B���+	�3�����A��.ځ�N�&m)�_�w�;� �Y��Oz*�9����|aMLR7�zm<��Xq�?f�1*_4��6������ޡ���Ѻ�uw�nJ}S\ýbZ�:j�Nc��K�J1�[Ui�wJ=���	�
d��w$��g�]F.6c��ǡG���	���x֒��Me�g����P]���<�g�ֲ��U3�\9��K�ǿ�X��4Cub#�������ؒ��<���Ԩ�"A+=:��=�M-c\:�7�K�����b@�Uk�;fI����){{�.�Tr�O�À�	��4w�b�B���'�lF[�<���Ne,p���36^c�}.���\ n������@�* [*�[��me�XT���G%m|Y�Ï�n���_�q.-�o�+Z�úC���D=$qG�ы�@�k�;�U��56<�:�z�$�%j~t䶛։lp�~�/�y"�V0�oȏ%ٸX&˽���pU���V
��!��a?@�b��/N1��o,$i�ۥY�;}]�����U#���j����#MB���E,#�%d|�4G�b�����`?j]ʍ0��⿄Ib��������'X�hՔl�i��e��?&p����Ά�[�8��O�����Ϸ����iqL��U�[+��vh�	���Fb�Ĳ����[]{n@b�p]x���jpJքH���6pF@3;�՚d|�y��~����V�lċ��2��Y����^+̥�4�$R�1�V����H��E�
og&$+�
S��ʌ���X?4��J�e���"����p�4�h~��X����ĭF�tSpm0�!�U�%+�j݈g���uGgw�Y��BF��䑧Q0�񇣋5Τ����S���ШԚ�脬�p��Ou�������K@8Q�p0�ŏS3�V��+������Z_tD�ҹ}��:f�6@��Wz媅�c�V��UU׆�[pi��|����/�ܚт�`ہw����K�+�����gd�YIޓYg�h�	6�`&�&�D��޻�s��@��|���qZ��ku�d���MQ�s��4�"�I��.���	m���	��N�n��E`�rm�������
#߀���c�*��<����=zj�<��J�v0bo(�����ڏ6�4���R��]Jf�u5�r�1��V~���zjJK�����&{8�jኸ�0�;eet����7>�8�2X�/z�1fP-$�\7vw�NM�w f��X�G��s��ts������s!�O����NA�:L�M�>D���a���\j^�Ґl4��+�=!�K`��fk{\�ƭc��Z������ޔ�A-�����#�6[�q�M+����*�C9���W��Es�� G�u:,m����m�'�Us��8��;N�s;0�;��}P�[����*��&O�0�[c���\�,��c��j�g`���cϪ�𢶓� ̊�](�ɫi7�85�5�o�����/��#{_���vP�������G��@m�! ������Me��x4�k+����q�1��3Y̙C��.��BM�6?� d��
j��A��>���b#�%��֒���q�c|�u��~AQL�S�º����ʐ��
[���R����t�n�R�5�{x|d��e���醀BN@�̺1�85o2gx`����`k�WO��{ǅȋC+�` 8����9�9eJ^��Ø������W���Nܰ�;��.�ᨉ�:�z3M���H�ْ�M5�v<���~�
K�}=c����C��U����M���2il�VS	��x#��a���R3�3�+�L�30��Ru��P�n�9�X�P��-���o0�q��D�9�<e����Ыg��IGQ���l�W=7��������;pu0m��ov��-
�.(�&�ܔO�1�c�QE�2jp4�6ET+����ż�I�Zy�)������#Վ��@w�y�;$��GEJ"*s�ŰB}�����P�c�>�Rg~��N��c�b-�j��@JB�Ό�
l�!�5��;9���TtH��lS%���{��_������8��t5b��61뀬N�sJV���o�\?�['q��[�j�ζY�����ɳi!�`U�Υ�J���Ty�6����,;��s�kn�4���oK�3�ar������=����:+�s�	YW_i]�hS�uXJ�@�vub*.���O)=�Cz��+��j7�]��@}C8)VF����y�C��k0QU�kѮ�Ȥ&s�}���u��_�-l���w�P^%y��1���B��L�j��������j7w��C�w���p5$Q��i�x�0lh!5iw���iʹVJ����������UT�1����)�:�Qq����`Hk)ɧ�3� ^Z��&5qE0dzx��璵F�Tުr�B�}���3��l�t���IliMJ��!�w�c5WO�p���FI��PI��������R����B��@C���v<�6�Ƈ���"��޸�$���Ԉ�=��L+EiG�@w���{�˹�7�;�K0�HUjk��a�l�n�d�.�3��x[�2�nPh2�Y��(�<�d��E9[7�[��D��hLq�*$�(]�,�!`��&�B�U�<������(?R"�Wi���b���6�2��l�h�&�Q ��-b�������=k�쿢�$"}���9�x#��U���*_�nﶘ�*y�	f2�J��c��6�,ȏ0�n�yx��.�K�2W�(z�̦�ف���w'"I��ڸ��4R���x��rU㴹,�]ۥi*�2Dr�	.�LR\4���J�4ºؘ�\S�a~��9`��Y��jY�D0�,� 1�\��rw/\c�� �E��b?�ҳ��p�f�E?��c������>��#'_g1�D�J�;����CWⴝ9�{s`�)����c��?��xf]z4�Q��ˉi�O��ǩ[�9:����7�aѻ獬�:��F����rO�pr �HN�����6v6&@����p/��.e�Y�&޺�{�EG�F��3���"�u@TD����",C'���l�~U"#�YQ������W��.�8EYM�#�����S��*QH��"�戙�=��X�S_�&��s�e���I	11�j���l�8J&��KI%� �e	^U��;����(;��W��/��#���!��!Yַ5�_�e��"��q�Z� ���bҴ��B̎	̿��g�Ob��dM>��ҒŊ'/�?�l�'��lM�w��}6���I��]����P1���>�m�>��|HӇA�:O[X�Pߠ�z��e�'э�	����xF��N�����������Ql캧y
�9:V�|����#�<J�R��M���d���T�bf��ʕR�Y)`� �����ZPu<oT�b�W);k�3{v�5�3�"�zlb�:s��W�Z�#� &��=l��<׼�}��nFrq�+c���VB�J#S�t��M�k�ސ���*�\Ŷ6[��m�,[��xZ�i�\���H:��|�ﯤU���[�rD�QQI�/Q��5K�3 �ъ]��KY�sc16x��@�\@�B�:�|�w�g6�E}`�_���+�.�}W^�ce��Y�ӽS�#	�L�G���;&�d�X���P)Ej���;�a̬�}�������J�t;���]��P+�VM}��@��J�bW[�K8�MD��Y�:6���w�^g��%)���J�	7촳�@���g	<��	+O6K�+�6�2_��*��:�|p���o-���V�:��5��2��@�Vm�6�|�f3J�t�;8b�>�Z�8ة"�/ha(.�Xf5����Oyw^p�)c�J����B<}�!s�r�7��@�=�I]7	���m� G!��mz0a=���Qaz�N�]z�+����8�"�&O(��S��)P��C0����<�(�ղhu^�8�*�6�|w�������HQ�_̥�~Ԉ���,1�-��߃m�;5�x���������<d��K=T�ϧ_	ǳD׾���;`�9��f����S��\��6S�Q*��3�M���`���#��-\zģ�#(��^��f��r<����Qr�w�M�{��ݾ쿘��!/�[c��\�Gɵ<����O���u��Ɓ"�_?`7`lZ�V�ђYhD����x"�;.>)8Y���*�X�}�|�~�i{�k;���s�F�٧�Gpn���Q?W��)Zi5נ��o�FT�Jڞ���v���IJ�s�S��O�zt��b%�8vfc�yCc�P��{�6�s\|�88�!)�#��v�%��i��F�"5�Ӛ@y��)�4!�͆"���V���.�#Yab��-Ł�@D�I�ν��r�jw4���sU��q��6P�?��E|����ƴ�����W�Զ}X�����i��׀:T�e�ՑI�l��B(| �.�^X�<_�J�(R���IJ>��rY��EL�<ڇ���b�ܺ+�w�/�Ŭd
���%A����ׄ����_tuu^(��&.�OHk!&��:��mG��5<�nd�:��f�s�F��Q��E�h�/�H���?�k@�����6o�b����V�r�Ab��\S�`
��A���7\��i�soK�s{���n�,�i=ߦ�ϰ��k��>��n��� �D��#��_#�м�Si���ȳ�W�-�b9i���3�o<D�~���ft�u\r��~�l�c��B�\�]��8�%%*�ISiN
]"^R�Ӵ��,�J@$�'�v���؃�����X�W[�S�0�p.�t�<AOQo�P�&i�`rkM���Nq���
��u��bkZ(_��Є�>��sM-��2@�q�es�ay������F&����)+�x��ZG�*.*3T�dlI�X��Ge7��Q�����\�Xi����`�T�ɔ��tkO���xo��	�_*C)�XG��`Z]��9fwEgK+<^�
ٙ���|�F}�+>���v�5;��E��5��2����95P��w�:U��2�Iu��3C�a���_�뿈Қ���
�ځ��k,:��jW���<;��aȌ|�v]y���`��=�H/�ܝ�7 @>�A �i��R�ȟ/������`>�C���U!CeL�<��1�M��	��8c�d(�%WD�(��}�F�8����+e�~���~'m}ݐ�^��Ƽ����������lYD��=h�l1L)4��}H0+6��nՅ����V���[�S�����·�dϧ .���u���Z �1C�3��P��`��a��s��B,������w�F�c�h�R��o�U�$��"�[�f����OQ�EMT%8��D�i�/R�!�4��c:�,���D�jd��]6���E��@~.4����ܥ3�Xv�dk�W�G��%<�[�-���m�-��R�a|���d�H�6e ����<�A��D�7�����8���P:E[�&�G%�\��8���^s���3�Q�z����蓫�&�kp�?�� b1�K�
�*	��������^��!I�0�-�I[��O��&�Ծ3�F�iNb�٠��W���Z�G��Ab���;�ΑB���\�tni��_������]�!�0�`<Y�F#p�!���(���48�`@�U��w
���k.�7yDd��K�钹���δ�|���.%���O�3�lD<�W̎��������M���0$�N�0X��Ȭ)�%C"�zJ���R(��9���Ӭ��Y۔r�C��2�W�H?3�X��>6�4X��ցss�l��d��^�d���w�a�t�g�A� 4����U	۞Vp^�!R�󱵝%�s�1i�CC]��.t�����>�f�s���P6���'S�,��?v�d�I�NAtI�N�������n�Ul
	���
IK?������&��}`�ج�%\�����m��t�,A~��[Ñ�ʩ�#���5J�;���zi�T��C-������³	��Mu��~C�4Ra���Tw.+��O(dm` �8?|Z?�>�⵻���B	�P�5��/Zƌ�X�-���B�!$#����(��n||Ơ]�J��l��FS�9C`
%�IU���2Tw�$���B�+%�8�cb�1Ψ�YF;�>�V�K�i̢���J_���cՠ�_�Hd��䙏�C���ب���E��a���fV��=��(����o��3��$+;�12�g����3p�
Q�Ck�8�]+����u=6ÕβT�)�8� 2\���f�"�0�-�eUpD�o�$�����E9T��$��OE��A�ԅ_���A"�+�l������<!X�+=9N>i�!�'�X y�2A*�6}}2����m7l�%C�(�ԖR�cv6~�i<
��ֲ�#&;��+��Ê�^y߰�>
O8���Q� �2x��k�l�nv�y�F	t�R^�X����� ���2.=�8���eB���`֣�� ���M��,ΐm�gn�[����v H�5'�� �B�G|�G��d��GI:E�����N�\Nz3�p0�&��*�~!az�j�ѧwX("L��0
���)�(k��P3���N��KX�4�=������̞=#o-}�3J�+U����#a������w��<�S�/�Ŏ ����O�]���/H������R�-�Gz��ء?jEs��� إt��CI�� V�t|��FT��.
�����}�u����unT�%otz#���T�+�'�8} x|vg�*(�e��h���|
Cs������bRw��u�\����Q���=��\ä�b���4��ʼ��d˯�\<�>�B*�l�����}�/�u!ilo'fӽ����E+�q"1��z^�� ��+��"��v5(	��S
H YW��Y�M��fs�q��@/�\j����$T2��o ��kl���(��=��}e�f� �&|Ŕ+�X�`"�]^��H}��0w>�'G������ab��Dk����2���A��W���S��`��
p��@i�~��'4���	$J0wD˶�Rx>��1�	�k5�YO����Ŧ�V�nIc[1lL���n�a[����}�w��S�G��m��!4#�o��y�P�)<oark�,l��T{:{:k�X<5p�"��n�a�6��}�VR����,.�T��H>�@�HB�.g�c�+�깓MpA��*CC�bUu?��`��a.�2�_^�/q�9?-�k��r`��� &K��)�:����S���%8q��x#|I8�a�D/{3L_�[�����-҉�+��pp��~Lne�3�[gkkY:����uر�e���g�a���M�N���r��K�D{9��i�����~�ak�u���}R���~o��jv�7>�j��K 4� <��jR�r��)���\�qg������5�����=�D9�k��va�e(���1�:'g/;��q!�y��іL@(t�w0���PR��jp�U��6N��"���@������m�r̮,���Ik�|�ٮ��9B\1������_S�mu�xH��_�I�UdP��/ * K_����S�)-����K�c&6�(��p�s�!�Z�l��h����>m�s�^��@���2��*8e�����N~�*	~�Ĳ ��i��<��b,�_\���gb?R[�U*���S_�擁`i|(��VΚ?)E�����=�|"J��ۋ�: W#��;<�2R��� C���������g��U��TU��pQ������]oĵ$:YϬ�r<�B���Q��]�RN��sO1�j ��_3`k���/�^Zj����ԭ+V�elHα�M�G�������Z�ҫ�	<��Az�����5�ܙ<|�<'d�"��S�ӟ	j�8�W֟nﾤ��.�p/Rb�C.�T�N��X��,�,�L�sT$_�~8�oE���b&Y��-�V�4�X�Y�yȿ�ߝ����=@|���cw
fLc�'uS��rAn�j��A�����r�ޣ��j
�$jE(�M���AHf�޶�h�����r�OmZ������T|Ÿ{�[����h8�{?O�yi׆��Z0�hn�	��Y����KK	}��k�&Ώ	c��vɯ9���.H�g�}Y�hq]���}ݥLn�g�͸$Nn*��I�"_Y�$���A�]���3_rj# {�R�0K��Z�_�i��Ҽ��C��.J2�;��M��na�%G.;׃R�o�7�b�q~�+;������zs�`��pP��Sn����@�I�S�MHB2�Rk���-�6��ts+k&��V� I��e!�2\Oc��}FJ6*��V��{�4���X�H�����ĝ�wu@�o�(9���1��!2��E�Y�)e�sW��YTM_����W��g�l�j��ӄ0Y������ll�4���c�R 3�b�W��E�iZP�J(ɿ�Lh*��/�� �̴Wf��'��ʱ�ї.8-��4XA?	�8�@<(�z3��Ii�9�� ��Ǝqh46�&�@�B�L�N]D��Z=���:�n�~%��{��|�r?�Մ��n��ٵ��ɰ6���uN�qD��:"kI ��l���E�$d���;�������R��{��h�a@Pe�"x�׺�Os�T�$��̷����D~���'�3�-(��Xs�[��m�X*q����=&�բ�O���K��^�j������[�=�Eu:�(/�sn��K�@�[�}���b�	������ʬ"+!�6q�S�5��A!��kM�\å��}H�K��u�K'�n_�Z�/��~�T�h˜x� !����,�a���%f(%z�B�>q� c;�1���|�������H�L�S�.#Cۺc��C|
a� mֽG�0��%-��򍧧��񆔦+�G�+(6����v�՜������Xa��,crv������M%�f.Q
e���J���O���2���%4|"�.`���x6�����������v�OG>OtJ���{,f=v��!�if��xʰ��!l3=1�r=��gUe �<T[�[i\@u�#c}Eϋ��J�..A�.e���!�c�N��^qT��^ɕ�����@jX�N�����)���8ے|�!G1� s��L�5n�l�?R���=Qct��~J��յ�+\�t���N�zs���b}�~v}A��px{�M3L�e��Nr��Ts:��D��Hj�Y�)������Q���n�}�� � ��)�U���@�� vȳ�2`��p&�,�~4ӧ���@�I_2��T�ѥ��q��8si)ߖ�k�@]px�����e-H�%-�(^4��ܻ7��;�M�OY���ND��K1H'	���[Z�����*���+D����Y�"��]�.��U�"	�f����T���E=��v�����=��]����<��
'7�ZR�$�Ew7���g��������D��L�u�!�����o\9��X]A
>�+P4�I�6[��:�]��R��e	fr��+�J-����ę����} ��P�6F���ix�O��X����D1�C\f�5��h Y10�9��3�ƣ�}y:7�$g���>pCwѐyK�Iн����]3��t�x�.(�нv��]��d�^y�%���}���J�"�O�S^U\���*p$��P���WWP�v�(䌌^�3k�5_J�ޓ�8@0���!I�/��*������z�.~嫆bN�)�Ȳ9s����k������P���̀��}��]�t����*�Q{�5�>�ҟ�g��&u�X�k�omLza滳(G��h�,|�tt�(�!}!8U1��~�d����xz#)�l������w��ԝ16���<,�wL����!P��g%��(<�n���ʒ{��z����-�&���/�Y�DW��10�]�c�h<mZǖ!:I0��fm7)��yn���Ih�D]���01��f��]���bR��?É�7�؋$�R�H��ŭ���&�#��ar#���c�'a=�NI�Vv�dQ�=�����)�6���8������g܇P؆�}s�'˫+��C�+B@�6;d�~���eY�$+7����ݬ�2���)~'p� T�����v ����Y�ΎGX`"T<jtzN����%ҵ�0�y䲾�O�ܚ���|�L�E�v`���E1�3�u5��$U����Y���{�qU%ۘ7��B�q&��f���زi�8$��u��mh%<�Γ�����y<�x�qpv��6�W�,��t��յY5
��$#��+�RC�3�t�[�����e��: ���!W�Cu��`Jc]��uhK_��aL�L'�����@�i�͌#�K��� �)��@R$^d����<��+Ő�	��fO3��-n��-�Z���{	���#��S���X?)^.�.�+s�?2#�ܤ�f�~U�G5����d/~���;�$����5���A�]�£���D�N��o���pP��W(m����J6�@�P��(Q��t���G!��y��B� �� "3��.=��by���!ݣ��k{(�f8=O���m`�nUɍ�Z�t'z]�6��oc�6B�v�����M�ɝr���vM�;MM���-]�>N�P�3�;R�q�D�$I-�&SEe��R�̞��S �wثߏ���߹��RY���n���K��ih��I=75��bN"Y=�k�@l�7U����y�T�I-����P~��Q���m���S���	ٚ��T�=���Oݽ��	�f�rV-��4���{���a#.ۼ�(�MX�rm��r&�_�LЮ_P�.��Xu1?�b,�/,�y�ISd獝Y��@�%�X����x?�g����#�k�(c���`^��9��yL�4�r����e����������k�x�d���h{<EtU�rfs��rw�r%� ك��1L��Ѿ��������LjH
j��<�"2���Q���I٭�^����e�h+_�k��3ؖi� �}�,�ї���b�FPD��=�s���+Vw<5�~�h+��f�N�[Q�G�Cvk��T����K��J8��Um�7ZSB�͑bځq��ۯU�S�_��ɈfR0�E�`h�ބZ,�MS���Νa���b`�B�)�m� �ʑ����:m:�{����:+���u\��}Kat�
]�����L��c���S���O����.zg}�9��ܩ�0^���4�m��_�1�-�W��9~���C�<��8(F�a��J{:�#�4��il����g����+,�[*�h�}���Ú�ٵ�K������*E������"#pP��_�~/�����_Lj_[}e�)�P�=\�q���:�� �:�9���� 9�I�dd��(]�*�~�b�C��� �	�Ţ���=�A����h~D7�]�?�����*��ͼb�:�ˡ�����}��Љ���#�EQj���G�����G� <սܴ�N]� �H��d9=�j�'�es����K���%�de1ǟ=����ڛΎr��[�ލ��ǆ��x����R�*>`���;���y�5 ��42��s�R�,��6�	�л�k2Π�Uq�H�<o�g����yt<�1�52���h���G�E2[,hZĎ�]�۲�2<����b2�J; ҃��c_�Ss�Ι�a�p����!:��,�+�n:f\�G8'�A�h�9�ʃl�컞�2�>g|�K�&���`C��d�^x���{�G��4b�Ա0��׌�T*m(1�m��u����B�ȇo�.��l6�8�MF՜� �<�.�?%U��BE�K���*� du���� aE� E��O�i)�����?Kp����c���Z��v���Yr(3�b�gO�GU����f��܆�#�'X��QM;l?��������3H�T��ؠ�B��#�Y;Q�M2bc��*{}&�M���Xݤ�u8SAE�L�p,�,H�x�G�/`|W��l����*�����.����/y���+_�_� ރ���]F�NAC<�#䯼R��V}���F��a�̚��k,��\U�m�#���i�2(/J4�!{����S�:���QU��5 >拧�ϥ��4ںހG��#�3���S��^BF��t�@�ZZ�	���F���n>��3
�ުw0�?�G�Y�S`�9����FN�|�flm�[����R���C��-�e���?9�ؘ��
L~;�#�g���c����g~}Hߴ���a矀�� oA��JA(�_�×A6�|�`o��'�7�u���Z���*?|�K ԫ�/�~]��d������kD�Ԝ��r��/:֘�%���b���L��X(
_��	�P<�:�����c` ��WX����K�t`RWNddjn-�c�B�6�\D�J�CZG�ݎ! �d[˭�x��6I��B��l`���(����d����[_FEM��p0�* �Z���60im_��Œx��~�q%�;�P�RAE�{��ƾ{�?m���,6�u��&���d����H�>����ce�zcV��7��QF�^��i^�Pwr���5I��R��9I�& �'7�1+���-ʢd4��^m&�yL��aȼ�	��x>�U�=��N`9��;���ʕv���v�b�kN\0�\ [=0f>�~$�U�%�6��*�K����4�����:-`��J4V�	J��uz�u�L}˜ҥ���K� ��4P�L9�%�Y��Ϊj�K�<���k�svtjʚ�_)8�/oB֊���u.�ĥםM3��H���}�+�];LY��7�r����.[*�`#��YR �^����F ���}�B��̶BH��OF��'�-����~�X%UZ�F�an7��9I,���jkĲy�Y���$���<8���ޢ�����(e�D�ٝ7o��'O�ފ܏�C����+��ο��o� ��W�q>erQ��q{�T�W0�zV�n)A��aj_���9VW������P���{�n����,���B�&roR�8���G\?Vy�պ�+��'�Z^���].���f1^A�Ü{6X$V[4k����Gb��fD�����$d!@w*�z��ˋ�IÅ�h�-r)�~[�_i��b��ەlG�7�u�G�i����ȥE���qS�ЮП~#:��亮$:�Q����zF�&������!B�s��:�Һf�1d
&��2>��pn��i0��W�b�i�E19^�g���l.��u�@��"�J�/ϋ6i���r@\A���R�W�����NI��8����JP��	�
��y)E��ɐ%��o�y�����}��\����x�h2��1,�e�4_[�=��}C!�to� ���7�'�y(�(�.�ݞ�3(�V�L�l��ݩ-MT|���-#���s�A��D�j6�n#E�� ]8���A	><�����c�ԁ̦sd�p I�� Xm�4��l�-���źe\/)������Y�G �!�fQ��[�_oS��`����_���Q�,�!TU��P�q��~K��[
���&�ޗt��T�n�y
������#��\I(�G{[��^[Vt�L�|�	S�x�X`�F��X#�f���KvŎ�$!E��p@m�Ֆj#G�Ҵ2�|Հ����&��m}km>t��l@���(��F3��CʴC���sr/�R�o�G��b����P����6�6�V�a��V���ӷl��}�&��"+��H6�������55��v	HX�L�6��� }|�'HW��t!���=�2��U�8�H6-.^��v3(�[qy	��R�~-j���jM��^I��q�kl��:?�&d��o�u�̣����q@���o�r=�%����ļ"��#Sr�l5��Y��N8���]Q=��D��GX�Aв�)�����Vy0��3J��H�Í�5���.�1�ȩ!@*�ꔜ�c��������*l��
=��Bb�uv��� (?��o�UP�ߊ��F:+va��S�� ᓅ��7^˪I��g�Y�t����B}1~ti�ڞi�?1��'��PBS[H�/Z��N������_�v�=��H�吙 GAy�%��m�����n��|_ Y�!S����ԉ*ۘu�'R�,�"͜�:b�M��b�^g�(���J��+�G��.֩C��g����:N�»2D��7��{�u��v��L$�A	2��d��XҲä�g�,�7�V����: }�am�
[�>|��W���M�B(����TM��}mr���uFt]Vy��>!���:�6����*ěؖQȘ�3�V�.mܪ@����%A�����p�'�p�C,8(#EG�]�h�����`�
���[��Iϗ[�AA���_j����(���;�n�B��f��[$a��{��)=�ģ�]���<@Tӈ����΀&��)�q�i{�p>�:`9�Sk?'48Y �I^�A3$�qA��L	V���q�ɕG�u1��dM{#:.�> ����ǅx�SW5a�6�
��%��5�s��4�J�OwJ.�{�����u�HU.�b��G]QFC�j\���i%d���\� o����4����
��[�[I/ge���,Q[���ER���A��~�ng�0D����Z���X`3� �yeژ�'Zٍv;ꞇHo��p���8�u�J*�f�Re�@�}���-b����é�U)l�����N��:�]��rE�����B`��.��a:Q�v��6�5c2�V�$�5~���>hqG�V����m�sٜ'<���}���@�@ӥI�RZ^t\5՚
���PN��������R��l)��[���>N�v1���:y�h+�K�Z"7�r����B%/S���ՃЂ���cz�{; 6769=��"ɰz�8���v�wL���W!�������,��O)_�B�P9���L%�:$+��)���R�\ %�S��Z�(P�����,�Ry:?0lꭒ�@#qq�H�̱��千��ܮ��'[]��t*%�A�\/�"D�E%֨�iaŷ0�4��Mtz6���Jޮv���{��!9������C��>���[��P�_( �q �^B�^������D���Գ5�0��dV�X[�kV�db��<�I}/��[�j�J�'�.%�~��O
H�ػ�D8��E��)��ߣ��ś�0 ���C*�w(��h�PIq]c���V�1y�n\{��L5��痂�H�^U�Ώyٶ����o�|i={�9t���,$O�����-�?��&Me�r�|��I�� �D��8�>tG��V�t�$��#�`��c\�݊���	N	3�[�S�7-�.�^u|w�4Iv`d�ŝy�E�P�Z���	�m�_�^D*_vsC�u/?@�7�r�|��~�v�
~g~^a�����{�5�iK��lI!GE�jb�Z�q�(pf�.���%�S\P)�E�?�p�oz	�d�?3kFץ,&d�F+4�_���]�;�6��z6�\�g���԰ ��^�7W��t&��1��J�%��]qk%�Ե�˛_&0��+�;�'�0y7g?(qz}����O�c�*�w?2ۮ��x�K�_�.J���s��O�A+gW�w���Ix�X����%r�c@�����$��~��k�>�n��=�F�j��s��ȟdqhlaMQl��,g���Xsk�̼$wd���24��=6��^����_�i�zT�{�?�%�^��Y��1�Y�J:��LA���Hup9��_����F��y�{�L����%�0��Q&��Gm�V.�:#�����>�oQ���]خMa� f�t����R Wj/CJ>y��b-��v��rP��)�2��%Њ�%ͦ�F%�Vn-j�\yΖv��nl���j	j��6�a�3nٖ���p޺Z����Wȳ�Vˣ*�5�\4d�6�.�Ђ$~��Չ��|�kc
�*��j���:ã�╣w����f���XR�"���%��L�Aa(�&nF��i�:'u ����ϧv+cKܗ�7����5�4�;#`w��euo����-�t���O8�*�n��jT��hZK"��I���<J[@��rEj��$mN���\�r�Gd�^	����{�M�����ӈ#3d5"����Cb���(|�0�$_2 ��S����8����Ѝ<�ӥ%-w��,5��kzoc\��/�[d��s��$'��R�%���J��p�7���1���!�I��rv�E�����f ����Ŭȷо�=='��&d�"j�	� #-��gNˣ=},J��Q��������4)�|�(7^s���뜜3�n
JS�w��a?>R�;���6�K���
��c}ƛ(��QB��O?MqV�2]f�q�N���A2� ��ED�7m��!�m#@���n)I�6�!����w��u�q����R���e�?�v�>o����+E�-����>�(|�ziu8�Ũ��d<�\�.i�1~Ƌ�j���8V��lk?Vh����G�W��)�ߖ�8����a�	�լ��jfE�Ul�	��w_�?`ݨC1����H�W
�M��M�����ӽU&���� ��jͮx@��漯�>�'X���0���dT����`��f42R���lo�s������Y��T�'�-�k�<H������qD��	���/�&�Kn�0a*�������k�t����J����-�A�w;d�����WRf��kL���	�l������#�˵FV*���m��B��)I��cÙT�"Q�1ޜ�R8����B�|��Ief��-���ܺ��z�e��h�;�-�8
��U/�AFm�ޟ�Ȗ�J��L��$�¹�n��e 3����5y�'S;cxHt��r=��~���8�BqC���HqA��(��u�l&��C�-
��ҹ�>iSHډEͼ�iZ�)��i�Vz�]u��A�%�8~�],�ms����T�[?f��0���\���{HQ����vL�ت����$рA��6�U�t���2�P$���7��61u������3v���y˄�co�
<k_��83��|�~�d*��1���='��](��
�Y��<����mr�!����������|]T,����&o����J�����3¨��PsȲJ?����Wg��r>��^M�Py�Qm�)��B���H*�_G�"�RQ'��Mp�
؏&��S<g�CDFkX�X�I���0V�-DS�8�k�@[|�z�|�sc��<ҷ�ޖ=�0�s��@�X�ܕ���JQ�RC�����z!��#>�fo��]��LFަ�SsHP3�[$K�0��H?��Z`�n�u�r�)�Xl��Xm�+�Y�u�C݈l��~!��n�:[���&�����4xz6�>>�^�L���.��D�`�U�,��7v�	1����?B�����Ma�W�ޜ��0|��7���ck����ƒdOr�뫄�41�^^Z!'sCL�7��� S��p���#-��+j\"�E�]obY>Ѽ.��
��}�����]�-��#6�����������kj��G�A\�����@����~�%7R�}���+�i�y"�zcz֠�	���݋k���W3������ٛ55�)��\�u�){e#y���F7ݏ:�q��y�I�nY�y4��p��� �5-�ڜ]�c��z4��u���LD4�J#��.N��]�����?�8h\�F��b��CO,o����ET���K��l2���J��c7
�\թfŰ�)X�r�=Y��n�Gfh�9	�\z�](�E���	(|6w�X"�<�ی~.���SmZ�:"I�g>��hƎ��w����(�e�|J���/��v�i�����U�x�\��#� �]�'a�ۮ�\��z��q=|���3�I޹5-��u�82Q"�������J�ĭo�q�.qrɤ[5.p>4����"g� ���#ר�rx���nC�
p"�����UHo{Um{�Sbk��:ײ��@%O]� T�	�w�.`�tg���t�BЄ35	�s�~������>.g������q�Ш+�3ю����uG$�y+� yn0G� �#�̈��|&=���2D�+��W��1��m��h��.�k���F�{�&�L}��G_9-���j^�?(�խd����+t?aQ��D��2?|��6BH����l��Q�fU��Ƿ)o�\��*���VHz��S9���Z��h����R4Վ�K�Ha�\h�8�3���$��P�U�t�q[CL�'�5s��~[��fOLP��V(ˎJ��-�9ksVڡ��Y)�@�('�i��f�/g�T�Ar��\�VU���4^fmn]����u��f�򧠁�Q�^Zu�a0��=�����C�c�/����z`7f�`uTr����.cK��'�J�G��,Ȇ3j{@ܾOB��ս�6����0�e.����+�O4��g��S�aڐ-���L>��1�~.Pa֑�ך��z��tl�1�r
��9	�5�^";����`��L��S��o��,榹 ]}�HV�C��&My�J�e��=<��kv
O.I�=?L_țپ���L����[y�3��d?��q������I(
U}���y�"�
A�oҞG���H���#}�r���:M�R%�j97�'T���;�h�w��M5;}��Q1��"R��.�'�Ȣ�ˀ�6@O}:�U؉�m�d��Tȃ������ǌ��[�b���{4�=���W�ɇ�B�n�ptx�y��u-�Y��wʲ�Nd��!0���W�z� ���gޗ���"j���C��"�x֓�XE�m���p!�N�~~:�����A�� ~��%'!�2NE+ᐸǪ�K7;��~c��e���\�a��]=iF�3�R��������ߜ��llm�T�����:�}�L:pC���;o9�>hIE:����+x�E��Y��S/���g}����$%��J_U��:2���}����o�2)����z��nv��h򊯍����m�ox���޼V�>�o�R�=�����P�x��P�#�Ԑk+�X�jqB��Yͤ��q���e�a�
]WD����1"^d�>��']٥��&Y���]��ɚ_��=׏�X#M�?xb���^������ȇ���zVޑw��m	
"��g#̗	܁r�L�޸�W7�����=2�� g������I����:�u��,"��V|���yo� kb�J`�XB^
�/��ɋJ��u@��ɢPF:���s�w�f��Yhv����	=!����90v��{Y̊�۱��uX>h���y<�g��R��tia$r��T�������Q�8-�(M�,��_�L
��M���ōTr'H �������b������lj��l��� 68V�%uW)��t�����P�C烄���qw�B��*t�mؑ����Od R	�Ɣ*��U���QN�H�-RΩ+	4;d�<���c#���v.V
2������p𦓨q]c�����y���~N6��6�|��Ӂ�5���E��񹮋6�c (�%}��o[P;4\�2����R�����#|e�>"�d�OU(-8�I����7�iG�=�OS��	�&h�o���%yi��F�VPSw&S�뱩d����;��j��� n��@�rw��Cs���qE��O�o�0B�w�7��XQ 9�
���8���@��|xS��SC�~(ͪ餍�Y&N+t���	����1^�1η专���"� ��_F��	G�{���B���m%�X���@CU���T���'E?�ޥ�v�C�)c�3oCxD�F�-P���5/_:,�.�� �¹]O�t
݆���᳧<U�.�K����|���54�����^������k�� o�\?T�ld���<�cqQ$<(TLJvx�x���� r�� ���RJG0�<WY�c���`6-�Ȃ�ن���g�2>b��|��,]��z͟DI�SZ�����\�DD�t��j��5jHsp�Qj�q�����p��5�/}_����T_�*�c>��9�ª؀��j�r���b�i��5�gtcW���0�N�.f�|�	��_Á�3���tl�˪5��il�Z����$� �b��~��F�h�z]��d��?���K>�����y)�^�HtDzL�}�V̧��=(/�%󸳰'���겎�K�3_
�o%�]R��Ó�(_
6Pt�����i����h�s�?i�����&D@>�ސl�E�� �w:�':�<m9Sc������^�������e}v�W���ll9��qh���"d<D�$��:0�o����� I��o�>�����m���D��P��Z&Jp]
6�PRJ����d�I��%R[�7���!�*@��5S��VUҕ�V�?=�Foo���tu�cߞ�B���+��8� `�Er��5��)���_��P4���=(���"� �q}�SYBH�ja�f�.g�Vzs��b� [�+�I�{�V������[�mI����~�f�O�c�1�Z�eP��sI�t8���/!?�)�/��ap�u�=axY��Ί��n��Z�K�.ai�xpv�e#�;��R=s���I��:io�0b�������}�w�O�(�{r�1�Bk�Ίw�`7U=���	,rq:�e�W0����MP(��T�m�jN�A��%��{���~CC���_�'��W��A��.��j	{Q��=��C;_��>?�A�IXӐ��k�Ϳ�E�?;�u�}b��?� ��٩����u|��m��Q���j��*��y����V�73��;�>�E���!����E���f�O�[�vf;�ΥS͙����Q�|Bb��9=+.1F�9�{���x̸!�����ށܦ����k��P�2k����̫ ))�,U�� `�6=/��~Ω�#�sU4F��'�>�� ��)��3|���u��MX-������G���q�nЮX��WY?Y���V�JϷ��U�D���!_}1��}�zDЁOt� �ܔ���gŉ��o��C�?>c��������i?)<�LNP�񰲭<C�Um1G�'���Ȑ��T�?$���5��O֒����\���Ć�]語���w4��[��>
9& ��yC[�]��^[4����q�~�ow�b��̀�iDW2z\z��'���$��팏��-�K_��ltӦm��X�W���pG�� k$O���[k��\��h��J�_����A	�����\o��Ywř��JF�ķxĴ�J ���`9���5���3��{�~q� [�E��}U�wTW%�x����`�S��x���~�ikr�������5��^z��!�3;o��@�sV����J\M��U��\vq.̮�]?�Af�n�&�|�}�}�|�գ�����鿂�g)v��\|t�.��⭍0b�s��B.T�7b{a���ԥUB`��*D��������8�F��!9z�bވ�{*��s�+����\�eL���J��qIb�H)=��GѨ��R<�kj0��������$�:'Z\a���f�ݔhyB��c1|ǅ˓��$
���'��Ѡv�{x-XͽmJ��:5�+������� H�y$��]ج�aG�5hÓ��B����E�:YA�N�G�6�Xf)��Awp����y��]��I��th�ָ;
4FfLi=��_���3'؅�@�'!��e�-��"!��)uv�0o�S�F��:�H���3���/���I����Zf�/	�"�\������Z���[�U�w�_BD_D�Q?3c�z�Q���n��T(�T)6"�H�<�pfN�AK�X́ڰ�^�$O�R��r{��׈�UQ����e3K�f�&��i��G��0S�=�b�ֽ�kg�+	~����5��E��ơl����Rj#�%~p�	N�f������N:g�����ú۟�:�3��Ί�Ϲ�PmY���H�@���~���{Z��t��� z�̸����,�"�!��a��-��V�d����)�6W���2b�ˊ�H&�jYs�"�}9^�g�3��U'	^�EM��c��D�V��'m��r1��g�����^o��3g��b���v���zW�s����8ki�����h�	��m�-B&�(Cx�)#0�]���?��;�o{�bm{u'�H�Ʌ&��8�g�v쁊����v�Ya/�\��!�ʫ�C��!��y�"��G7�@�1����������1!�}���y����z�R����"�-ګt8��/rU���,ȝ*MM������?��? �v[�p�8�ON�>�����5�m;�C��Y�pw�i�Cb���C���
�R��!)E9���a���ç�H8���x<�i�`�����k�<C.����E�ϣ��!B���r�;�]E�Z:#􆨽E��xQ��Id�&�*!u6�Y�ad\��XV� �Ԇ��_�{($��1�ߗ_�`�+e௫�����9?:�	��d���ųս-<��ڲe�GI�H���Y���zW�x"�A���g�K��_G/�sZ,j�h<��yZ��m�2i�<��^�d��'we0���g
�r�sw��{�xiQ���u�3u�ѾCVt�&��&n����"�ǋ=�/D*Tz��T�s׽%P]��.��޵�=�C4r���2�eH���$C�\}|��]��S�툘0m/2��j{�#�����p�З��ztEq��8�D$[���� 1<-`�RMe��!ѓ�y�/�i�6�  �"Cx�Q�������oxe�����? Ľ���xYM1����� ]��y�b�ޑ��%n��P�ڐt�L^���_��tȰҧĺ_���П�����v�G;3w��㖻�]2 ̅��C�s�ƱR�2vE�y�ݴY99��U�RvG�UJ�x��N끉���>V�W���O���t*���y&���i�2gh��a��B�y[��
�&�A��ɮ*���wR�F��E��N;@��'��������T����+�XrR�{	����#�as;����4'���P�2 +L��;Ԥ�L3�0�iN@�N
�FR
d'~�\�1�n�V�剕��ъ?>]�4�6�f��6� �NXf�=��)��=��kƔL�L��g���m>��Vߦ ��zb'i��41�9���C����b��<JUVgO4�8��1˘882��Ay.�}�)Tĵe{�C��E�t�@����[��'������<���;v�r;�T<�`&�ۥ	@��,'!��	����S�eȺ�~��H��p���?����s��w8�`�����lz���T}���L2��a$�������WDŏ(�^:����Pa3߿Q?�,/o�&�]=)�Ӫ*�����>ͨ�K�@��C]I���VH�Ar7���К��ޟu����6 ���w��B���jаB�!Q�C'筿��&�ȡ��m!���v�X����舫�4����mk�c���
��l�c����A��$ ��m�/O�󣎈W��2���q����8 ,�`tW�nEy�=es��I��fP��{_� (ܯ�*�D�+�X�fDj'*�*��)26J��Ԓ�pH�0pD�{�3��m`���f�l�?8Z�oT�c|� �t����Q�p�;�c��������x�V�]:�'�Sߺ���0��D�R	�-�������-[��n+/���0�9�ʄ�Dݔ�"��FFͰ�F��:�֏x��R�4�rB
�(`��%�awJ�"0v��WxԞ�ru��c��J�����u�r���$��1=��W�Ҩ��Ϲ?"�Wݔ���D��������\c�6�p���*N���<xxq7hV�<f�fZ�_�j���A��I�o	��Zm�Yq�l�>-�󔾙���+�ނu�Bu<��j������L���-���{��b�i#o)������Ї�*qp�=�,-����N���Vt��w���K�y�fX�P-"�*8��{��zN�Ĳ�D>X�(�i��8+WxKN#�;_�y��|�w��/3Y����v�/��@y�N��n*q8���s�K����y�KE�IC5"�k2��k}���Au�v-���9_��mUU�	���#�V��Fw�J������+�p���,��E�c%�X�hLA;�������LS󼰣)]l娰�6x7�	�n:��gK_� W[i:V2����M�(v�Dp�*�Y����ET�x�J��aD!<�$�~8Cf^sK����"�=���il�\)��?��	=�O��G��CAf(�T
I�/���X�uk^�.�xCů������)MO��zb��^�M.������E�k"s�8z���n�p��tD���QDZ}�]���}�{�H8ĕ�d���J�4�5�a��'����R�)�� 5SǅI�SU�����/,��h�������1�;�'Dg3�A�OxB'�fy���0��;F?����/��Ǖ�����ϻB�~�@KF�O-�zV�fj��:M�,jxz�'�H�q�4r��1�b��.��b�!�M��O�}�e�l�`\
e�*���fa��z=9��AYy��ҕV5��cjD�w*��-���P)�\6����"YB�C��ꃍOh\s#�	h�IG�=���,���&��B�pS`���Jم�ƥ�pMR��HG}���2�c��#�Wh��X�w�~�\q
�����n�@j���N�L��&�lB�r����:
�oL�IMK�J���X1�3�)�C�uP��O����U�u/*���(��c�긇�~��cև�Z���F��J뉾��'�+a�̺�cK
��(�U�7�1d9�lk#sRqG��sq-�Bvh��E������F��_��x�q!�n�{���_���U�j�������ʃ�/��sU	�}%tv9��N6�M,Y�����F����J9e}O�-�d�]���)�D���tbC�ۖ����b�#���/�E�����Ӻ��!��6���"X�e�
�ލ���yu4@��p�$D{N����Ê��P��<��#���a[�}t��_ܪ��w�1	yX�!Hb	L�D���__�]��#m�V<j�ퟴ���k�Ŝ|U��ܑ���z��g��#貂�.ϯ�Q�g��Pc�zk��iK���Du��3t`�t�`:Ĥ�~W[��A�˚��՚#���pL�F�x�5�v㯍|���?iՑ=��k���6�[)�ԭ��Lք�r	���ZF����G޳)G��G�*��#�L��]����%Ș`/ ��݀�O�z�F��V��;N�f{�ڱ�Ɏ�H`XWE#BH���s?�QҔ)H�7{��"7�����rb|V#f͞�S֠'0󀥜J�l�'��E�u��0��zG��[�v(����0�jQ�,�E����%/�}�+M�j�)$���Q��6����3��&���������<W�PB�jr@�ۭ�wTB���@� 9�����vfm�F��|�  ���8L�����JB��Wdi<�����	�4���z����H�p"�1�|\\p�f����ܔ�+� ��ɻ��W�fg��ܮռ��C�[�t����>@Z4�Zq�M���c������u:"�`?O��!5yK|���?l��@��K^��zcA�`�)�;���^��Վ`q�X�ь��bD�5���Я(�?t��Z{���S�bO1�Ɣ\�I�e5������ՠ�^$<R\XA@�X]�%��u������ś����:�����`��=���#�S�`��������>�0��dDz��Oֵ��NJ���t�N(�L��}7�a/!�л&l�*`�ȉ	 Z?���P^�l�lg�4�8 7
e+Ѱ��W�	��x��*�m�<u���1�+\Ai�Դ<��./_&��� z����ڜf�s�,�-�9)�a��aw�[y �~:8 o����Qԥ�����@���+�`�>�?F3���$�t�'�Q���Zqiс��c3�f�*�aE�N�D򯕷��^�b�7^�YϷ��2�y~;�R]��5����N������:{�y�y [�{�_\�$�N�c
6�\�`;�����KǴ ��Zy4&� ��&+c�rݲS �1�a�9�c�n�䱊�ejќ���4�X?�}B��U:�t��zo~�D:�Zu5��	C��%��,�0�b)�lg��j�q��Ʋ֚
.`S5*!��i�T���o�C@7c\�����1]�a�=׮�	ZĪ�r�C�_wڨ{�����r�ke��ɟK��?���˹Ϛ��E �D[a�Iޖ�8��\��,e��)����@�� [��j����6�>/p	�N��-S[V�
XY�M7����l���W#`$�g�CRQ�tW������cvUg���0���c�Je}PG-��<u'5wjl�=��o����>�/�O���*VG��R�<���HG������|Kyr��OV�&	hl����k�@XO�I���@�%bσ���6�ym��qb E���$��wNsS���T/<`�SZu�vԸX1u>����}��+�t��Dy�z������=�NdK�GƒC�!i�W*(��O�x�h�'Hb+b�j�;�<Ұ{��y�'|0o��F��ۉ�+�@m�~���ЯNF������Z��i���Ю7�!{��@gsǡy�n�b����Oܾ�>���4D"����(���>=�C^�|�t�s�<�+9�?�P���!@��FxFw�>r7>�����5�x:r`����u�[{-���sP�\������z��8`�,�[e�T���F (���%�-����Ed�tȰ���z��j��HC�Xv����T������:�B����vs��x��3� ф����X>^H0)��O(��/�|�E���$����2����$��#&��S٪�t���}����S5U-�)�N��cF�(I�Rh왛��O� �.f���`����k�3��<k_p�=9�D�[�C�nR���.�h��kѷ_���\��E�9�s�Oy���R�}��F��o�T�������\�Z������m�t�n+�[��bۜ�E6`��5��f��(�VR�Df���q�����7��.� �&�5_8(�	n�~�T��bV�)�W��˕*�H�
x7��9���d�-�t��1����Ě���	�T�)����ǱT�~��gHsD���=��'��W6� M෯Sw��͔M�� Ƴ{�xf���3�B�)5fo��i�}��D!|����������q�	f���I�-c�Z���R�n�6�#|Rt�)E9�$"��R�|��>N��jӹ�ov��hF��3V���p�{�_�S�|��,�>_��������1�@�k?(��&�G]�)�
N�kD�7��T�>�8(��YFE;=��jN�!���G�,�f��c� �H��睞b���I���;�����=P�����[O���v��^�s&��)U6��>e���P���`+���QY,R�ZE�`�8W\J�i�p�2E�ڊؾq9B|Hk�t��o��X�\!.B��[_�B������i^Z�"b�;��� =O-�`5s��T�Do���s�-.�C�4��{$��%�nȶ�%dXK�_�־���f��fu�N=+|��5�k�ߒ�����H��\$D�o>.+�G&�����^���Rh)\���/� e�%�򙸪�:'��������j���<��L�%�gP��C>E>�P�x���x'�-��&j�	۱e�;�{]ph��gf��������l�B=f�)^5\A�gt9��(�i&�����Q3�N����M4	f�{�V�K=�jU�����.�(WKU�V��8�;Z��^�4j	�'
��p>��U��\B�c�o(���ܱOu��:���ZL��s@�-X/�g��kL�+��Eq��h�}H�`��oY<r�O+�$1`��2�wC�����wG� -}&�ߣ���=nI���-�ԦZh�2#N�+|6�I]��=q�a�練�tVׯ~iϹǑ2��W�\���a��+����|��j"��q�ii���ɛy�G���zO��c�9��.����.e�E+䡓�H}n�����d�e,�u��V�C$Z�����5?�����gB�~Ҽ5�V��Qh���ŀMC��&S%�	ŲLc��8���}A�I���EPnP�Y�^� t%���pȜQF_1h������,Z��o�P�@-�F|���� ��L�O��%��H�u+e�۾��P]H�2�Hp �#�l+Kp�8<�4�Hȣ]3�R�/srMcq .:=͏W�-U�h������/�57ݴ)nD:̉n���k?e���&���o9�e)���2e��ܯ3g�,�r���D�z��:W�c)"z���r8O?�df��*��<zO�;)�E�h%]��F�V,{�p�4�EJ������r�Z�Dr��\3P���Z_x#S�v:��e9���S�D��6xAd�D����I��*���P��H�Zo�LUw^PU����N��|g�J����Ձ��gB�����S�ZB	?d(8__7�g�L� �}�l	��Iހ�tFc�{��F�:Q4+��r.�!�R�R���mF������0�#"n���ϙ�����U�Sm�t_u�ˁ/�X]�����.����o�P��������\�A�.�^'��Z�?-�^X�4;�g��a��Į(;��3��7D�Ƥ�b�y��=�w����8�u�'���y��Qb]�fD����8��v���-%�a�^����[��D�FU�K�^�J�I�d��L��EƋ�l��W���(��P��9A�8��[�I&]��}� ���8���XWD��e=��h`<����>�91����?ba ���)�;�*y^*�F���R�#�n�G �h����^¦���2��&�f��\_pµ��T�tf���	����4�6� 7�o��<@�׹�7a�f��[���w:��΀��kǮ��^y��[��Q�P��H�oK��ϭ)�P�r�̀��jdЫ3�Z����P������oC�4����5���g��䣰x��Q�t%?�xέwԼ.ne�eyזy��s��o�r�W(~�`�P�(�+h; �]\����a+��B�u:�Mh5��f*^M*���ݲ��7�X�^c�[Է��z���U�o�N�e��j9Cg�X��`�����癨i\��D|�����:�W��^�!���e^�����ļy����JÆ ��Π��d���{Ob	t|Az�01v���:�4�F����0#o��61�	k�79*���y�ך5Y�*9�Q3k�٠�h��;)�R�.9V�D�!}�7q6�ZO�N4_���,��x�UԺ���J)�%h@qt�!v�� J��T\��E6܃F`+ ��N�+DRa2�^�?�&�����ˉSr=�uN&K��U��TRd���Q� ��Ap�f���N��/N������X�����q��8��٤�=�/n>Q���j_'i1�c�4���WO�?J�M�[��^|5��G��6�ɩ�]�,ߨ��Y��g���P�w�ۚ������bs�b�h*�u�'��|A�2�Ci-!���qm�e�Gv�"T4��Z�yϐX�Ӵ:�2�D��+�}�b�b|nZ&���rGcό� GI�ضm'�Kq&a�
��2��9�$��B��U�a��R'�^�a;��:W�\�D����hO��xe�I&�j`��n��`��@
~�[��E�%����%���o+-y;V���?�ߋ誤ȋ�j�&E�@
I	�^�Ȣ0zW4Gԡ��/ӹԛs8|�C&�5���4�B8�T��7�q${��2��n��lH$	�.�D3��&���F��{��I]����f��\ԅ3q7%�Rd׵ғ�t&m2^��`$��.���,��9S�V��ZA8��ފ9M�tCT*;�'� ����~�;R̻��t$t�A�ys��!���Y0a���bښ���0���c�|�Q�L+�?�����I��H�������!S��kD�H=�i{r�1�i�K�����Y��Q �&�_ս}h�"��a%�֔�O=� CǕ$9\��M�-V�����i2*�}���hk��0Z�-��rYN���x� Asi�Ӊ���Fv ������o�=A�af�>����۹��.s��)�7��\�"��zǴU�n"3���n�\��t�N�O��%MWw"����X�[,,�I>��.���e�����
��>�%~���uJ�o�9� ��G�<sX�^��r�N^�سp<T�4O>F���WjS �/2��)?8��@�`��՞�~�Z���}�t�j5�ˎ	z
杰@Hl�;B��ʹ�sap�3R��S~;�I��9F����[}�?�؎Plՠ��N�SEٕ���&�1N���+�*z���ٔ[m�����7��;�F\u��0Zý�I`�BQ UK�%׿uU�&�0:i01(>y��qT$�pb�xw��Y�i=N���?4�A�h.�2�_��z��9_^"	f��l;=��-��x~�i&�3�b ����ڊH�A��z�d����g�w��-{#.g�f�V]�[~�2�����!�u��c[�;𘻚��W����J����q����A)�
(�)e#y�i�u�eM�-)r�1ž�;'K���d"�!��D��&}�P���(f��:c��{!_�# ����%)��q���JUѓ=������
���^i�m�U��ؗ�c}���"����)C�����۴]�$b�fMd)//�����lM,��E�Z!�ۄ_�\��/�YFÅ��ֻ}뫆u����{tm�Ʊ0ڬpo{ĺ�2�iȘ�
�o
��������VM�7I,�0��^�MGC�/�/&��|�}�@϶%g0��@O�P��/n˛z+M���6߬I���7F(�=!���
.�ՔFOS��e��d({�yPPZR� �G^Mz�	�����t�C��0�lĘU�JFq>4�T���{�Qk�-��M�[:D���.��w����ak�@�s��cX'�^S��5�%���:�l��f<��z��0+�=���S��\p��.�&�Y<�74�n�2P�+�2v�@�Oz�{�mYۆZ?�	�y������+I��E
C�:k��e�Hl�seUT�}:�l�LVg[?�P.��$G��)jt�0���EqtI�s�&?U7�; ���>��:�'�9�"/ü�m�V�n~B8+T���L�#v�0}�'��A�r��ǭԤ��b�?�X�8���M�X4�a��-)gx�W�*ɿ䏙�@̮��ݞ��Z��8aĤL�~�!�Jl��?�u�@y���06�۷P�����H�bO�_)d�E�c�^H�i<�%�:I6H�Bb�
�Zy+���i쁛�0@���#!J��Z� }#�\U
9<�2��B,������x�3��= ��x�rVV�	�7hM�ـ}=��^�C���)�lI�`:|�~��M
#(�2N@QKd�1��ڑu�;���z"qz���(�h�8�&�d�xm��:?��B1���P���٭S੫���\�P˨3-�A3���T$����������������]�X9<����Nl�!Mn��h*����꙼u��$�ya;O9ud���Jc�\��q]�H \/�֎�ۻvz��ʌ:|� �O%|�w#�{vwۂ?� ��vβ�=Ǳ��@����̭^NZ�k�/�=�w�L۽�4j~vB����nC�q�;��b�%V�����_��X�Z�B�~`ue�[���@�-� *�ަ^C�'?�Mwd<	��23D _Yd��J;�๣Cw}��Ve��,?��$~�^�����`~�ׇ�^�k�3�i=�Wؚl���Q���i�5t˝VpS��;1�PT��mc����|�B�V��z�����V=�8��� ;�X���$-�V�3jrpe�ۿ��GZ^�����1#�ts4{��#uO�|o��_���\'�.ы���� fhI�^]JNG;�'=�Dr\�T{�	����7�S/A���[S�^U����n���\SNX��&=�>�8�Y�+G�4��"�}RW�v�z�� �*�+2 ��2��h������E�8"�B�
��N\q:�xՕj&��b�2~J^ڷ�?>�"�mg~��k�rY���Y_��J0�����.����`7t��+n��ϑR�ެ�X��>m��5SV� 6�43�.��8v�r��U��^�o�Pߙ�M!�(�F�64�Ӫ����L�hl:g,����W�&q��݄�e���`�/�c��9b�g�����F�����#HK�ҹ�4��CT�N\��y�ϧ�s 媐+��_�"qڟ�m�s��7!g=
�xx��P�0�.�R/���.=�e��̽�a��*Gu  g�$��i-܃(B���Ȃ~;%���.W�W6!�i�V�٨������S#E� ���b<F���毯�IMkK����%dg#�%2�^����)��'��3y�}}��>�l���_*x<�O�$�~�s��8����e$Ql�>a��[ ����TS�1��&K�
̓hh��\	�+ �Z���-��%����%� ,}�yO�?x����M	+��ak*�Ϩf��
�0���>��I�B|����+������2L��]�a����q�9�b��B(SP�ׅf|��{�@_5�<s�^�|�I�+Jqv�%��:�Pd���,�?��#����bs�^Ir�,�\��qt2$%��1]#c������4��gNM�mxW)��?{6�i5H\>�ފ*�=�
����&��c�c��Cb'R�6)�b`9���ľ������L�;�JA 2>$�0/���ҧ���l7g1		���e���9���� ��v����~��ɟ͆�#G����$�>��F+����0}�r1&p3�"�;7C�h���-P���;�����U	;�ͫ굽�&��oE����� �>V���K}m0N!q�����-�t��aFDa�'M~^o��O��I��_>&���%���R{��mM�R��v���;��7�TtCq����ǌ�"��0V�ѿ�{�W��:P<���P:$,�?3��)\���R�U�^�nӇ�Â*�|r��r̈́�_�Q_�tJ���+��%j;�)+�.�CQ0� 9��)�^\�A������:}U�:�
���*��	Յ,�)����ʓ��� �S���g>�<����͘�H�LK�:T����n'V��Q�����X,�+ٌ	�tU�e�)�������~�w���>�Ȩ#���]g�g��@(��ȢFpU�ޗ�_���&�ex!H�Q���O��'S������@i�=W��+��G����cP�BQ�hQ��x6������+r�W7��h��(��,8�Nօ���e���(a׹�9+�y󩼟}�H���#5��&\{+�Q{���#�u�=���@���ƛ6�_K$Q\�VLa
�9�J�Wh�g$_��ǻ\PaD���)�^��헮��Z�8���&D�7����p�q%8���XV�r���$h�on0.��R\\IHxn`��"Y�����Ç���P6'�=V)%��J4x�?P^�?�gʌ����^rY^��;~DI&�oP�������~�wt�Pc�]y2�����b�.v�ȈQC+���o�X1E�+��BUQ��#�'W��r�ߋ�}����E�aW��Re8S'�4F�;��<�@z�tݥ#����@Z��l� >����Ox�f�ݿ���ƬN~������+��NrH4ƀ���fՆ�{�Z���/x�pvh�w��0)ui1���m�N�^��K��[3���[�����f�&������i��������X�ڱ�VO�K4
�R��Q�@O�=/�F���񚉮D���
���B9jm�R�����~"�6�1�&
��}��K�żbf��3�I�7I+Oaw�-=����p����>�n�Aq"��vE��h��KDַ �P^�%c���{�Mf,U�g�"�\�O�s�\#���&NîV�uz�L\J���ŌL\�IuG�= �*����[#��#2���DEAQ�S�e��щ/g=Ǣ����⊴3~AE��j��1� ���)2� p�v��Z�Gc�^��R�Db�p�q�Cy�����N;����	w;nu3��w�n�����L�"�>��N�ݒ����&�ų\�d68�5״1 4V���6&�I��ez�A1T�>َÖ}��ř/����[�ID�z�Ս�VZC��YPS"���wv'>��Cm��q��}?i7f��r���"y�_��%"�x��/��6�ɪ�P��>�ड़�����+��l+z�s2�DP��uȭ^/���OQx��p/��a��]}�%
!Rկ~���6zZHk�=iC[�yte%�J7�c������03 �[���v&�=��f\k��?8Jÿ�L^�$
�fr����_-�Q��J����lW�?7�}�ctPx�|�r���w����Vq�[R���/,�Ƹ�jս(�IU�3����t`@��>�hU�;�.�	�A���W�� ���1��%1��`���yv��5���}-���-�E�yiwe�g.'���˟�T��|a}yT"�/祍�<v���u��O��C�xwG� Ф�9���b�����3��{����srS�b�yfD�(�VS��{�����1H�����!#��Hɀ�)ףU,LM�z���ę 3���YR-�%W9z��1�\~'���� 	n�2S��,�W�O�yr.����+i�Č�r�P`KP5́1Oj�0�!"]h�*am���-����?�f��� �"������2	y-����S�Q'���
�y2�N�+w���YL�:��L6�e�7�U}�wV�?r;CG�E詬_)�Uݡ�� K~i����+|���u>|p��א����׳	��0ף/3�������t������_Ep]u!���qZ�2����T�2�`�?!�[��7?ܷ����&��^�g��]�u��b3_ۼ����/�:v�V�ɾq�m�/���Op�B�u "�m���̃�?�P�ֶ��9r��<�6T�c����K�@�J4jD�m䌆��SF}~Q9$���U�#AK6?��y�jl4��5vl���v�2��8S9%�}���f�����X�$�j�U����,��RU1���w�nϽ��|VoS�
�u'�_a7��n:�ɨ��QH���C�RR�6�����N>:�����_A�G�՞�,Ѵ�c��m#QEj.��/��1�Ӝ�@G����k�2��� XȾ�7�Ѩd���l�>Qj�)�����C.B�؍),�5��f#V�BQ����ɛ&y��jD*�I�~,|����P�ʳ���}X��$��nEOqq�o�8�1ɲSG�O ����Hܸ_@S_��P��]���\b��˳��)!���T� bB�zX?�b(��|&`H����T$�!u*!܈+`��R�!ة�It��u�)#h�R��G��v^=aw�1_��9UzW�HS�2���U�5��}��b�Ī8�
���Ib��A�o�/<�|�V�U1E�K�d)�u_�VH9���}��� 6��j߯2[~�s3�3���E)����`G��V����(��[�+,5�/gXg#6F�w<!����iC��H�#.�в��S�Oe<�)�SJ�[;� p��yK��!p$aޟ[^"x��!`�<�%�/��?��V����4
8u��A�Y���nT��E�j�L�OŭQd>\���c��?�~�TZ�ϓ�p~Ց2H��Fq�����;��gN�.��KP�*Cb�}���f���h���f0�O�XW���X"�$�=>>�F(�$�9�W���:~��|�_,�L"���13��5�V�%W:��V�z������;�[�Q�kt��~�)��b��ӆ�Vc��l=�x܁FR�Z����N+E�xo� ֲ��L�_���K��.�d�B�֊񧟼bH?x�>��<J��a�	�m�ߍ����s�E��Dv⠹���'�G�Җgx�ΦA5Ī��`[���q)%χ?%�-��vM�Q>p�	����#~�Qǫpg�|��V/����p�)xǻ�� f��G�%�t_3Zo�q.��~,�ɫ�,���s��ĔN(�rm&��#��e���T{6�ޟE��b�=2a3����Z���ǥ�V+�3M��=%��ΰS=;Z��4��\QG��h��q�����s!�����န��s{�y�Nn�ǀ������X��g�-t�%�(���!WU&ޞ���-�ljX� ^e�CO���I������K	�e()���W��8;f���>Dds2��	W]�v�ʔ.J�T$��e���vSr���$^	ཆ��.:�_���&�$$�;Dd.&1�q��P˗:~Ɲ����"�7�^L
�w�M�52�ٺ0o��YE"��iT(`�i6�X�`���h28�c�5���H��8>8��B����b�"	�c�����g��'�r��8��m��8��'��d@�%�V���8���3��H\P7OBS���r��d�j��ơvt�ϹJ��ҫd�dE��X0Տ���+�����F&�+��鯭�֔j(�a�+R���`m����5/�l���+��q��vЀYP�?�On�"=}����4}};��t�F�켠�Sئ�U�����=yכf'�:��P�����;���9�?a��E������^r����n��}R�1����_����Դ�7��� ���,���f��'����ߑ`�H0�1�]<n��^���MRa8�T�_�e1���NF��{��4;9l#�YDr��~C�Nf�_���sH�L��{�p(x����P=� �B�hh'#+G�|���rC�䎽ތ�i���J�vZX�H�������C4�Ɋ&��I��KK	�6��6&�%)�:38M�L#�N�� C��0�Q${FsW�� j:���
�D-Zi�g�c7^Z�j1s��)q#R��1B�S����4�Tx��Y2�b���G�
U-���Oo�y�;j]2X��Y4�;�o&�P��,%B�]��ɵ]1��gP �?�>���񨄎�&���M����u�o�.����f,���|��c1>י�E�\�K��cJY?�L�	:��a�Ta���9\�h��p�����
��*'�XR�Ԏl[�,=�Q'+��0�D���l�g�v?<@�Z��۹�cT�=�Y�]�	�Lr+Aq{��Ԅ�zY��q���h4�:o����t��
�j/S(X�\8f�dӠH;)86aL�yx3̕��Ǚ�jY�V&kk��:�>��k���XDjZ�M_�wc�;6��~NZ�A|��u��)+�	�N1و�Wn�c0%S��6w6����q�9`��Ԟ^X��\����i�h9��X%T�('��@�`��a�m������ ��!ި��6�G��O�A�d+�pL���paXV ˜�.�h���c���xMK��t"׬�giH9�`��٘��n��Hx��=�4:�g�ҥ��\ڃ���B��Z�^+e(ٲ���N@�D�Ȫ����/A�](��Xd�7(����a��mҫ��?2�H�}0��<{���*��n�!BDv�p.i�:���ڔ�������i�<��E�t�&�]9M�29�!gm��DoOd�lo��?���x���~�q�/c]���I���3�e5����Q��>M1!a�E	ܖB7ȟ*�m2��ֽ�sk����n���8�0�.pRl~�mK�O�P����tY|=!s����ٍ�����1D,��d�L������]xΞ�A���aR��S����z���XL��D 	'�gi�ث�� �}zv�I��KQ��6��tz��H�ݲ{���e>�,��o=$�9�*ՌE��[D��e�<�oU�(K��x�p�w�T�3�ym'�b��m&��PP:��O\`<�8�:,��6��� ��k��[޾�z��_�T�i�n�l���iֽ֡��U���M����$��Z�MH�b2]��'����e�"��u.)�є"�1�a�d��[���Dp �(وD?>�B?����%qdE�l]��r�K �CT
i@i�9��7;{.pI������Xn�3r�4_	��ҡ���Pg�ˡ�@T�K)Ј�eϗ��f�T��b��
�}��#֞#��l9���!u�S*/�<��q��ڳ��16jڄ�)��`=�.TKT_�+K�$Bʧ�H`ޖ�U�͸;�i�Iϣ�Q\'TK���IR�U��]�0�W��[%`	mE ���٢�]�]�h��6嫖k'9����Z�L
w[�c���`1�cRT{�lkH�6� p���I*QB�c�����
��@�����R��Z#�Z�Z/���w�Z�D���I�(��"�-ʋwZ�9g���e[��:�o�1�A�s��U2�n�W�;N�a���M^����F�)5��z���H�� =��wY���'�'� v�>�@�W���1�U�8�Iצ׭����ε�3��}��S
Ko�׌'_[s��O���;
���TЂ�����[��E�ݒ����4G�ag����1%mB�=��ԣTxv�CN��C��r��4�e����Ir��
�����4�9���z����#\�������D�/���W�^֦�=�|!��e�	V��=�dSJ߱GӖ�ĳ<뽰��E�͐c;A6ġ�����s��3pta>����魝j���dWF�k�l�B�*�2�表,��Q����r�HbV�:d��
�$�2d�����s���r�> 7�`F��yF�ٻ>/����[Tg���)��G��� ı �g��cb��P@���@��:��8F��j���d��p��!�H'Qx�����v�YT���ߗ�o8��*d!�f��b�!6bB������z�/�b�r$��K�,^���^o��^����E�ڣD.&��<	��fvӢ�a�|s,b��%gL�#)�8�ڴ�"���F�s��P[MTmPj�s�_�t�)�u��������7�χ��m9�!�}��1�r^awm�<-��!�
v����O���*�O�K&�`�0�H��K�̸�����
C�p��4*�Q)���H;�l��];۞�������H��p6=���?��������������c3&D"�Bo��#����k�	=��-^G��o}���¾���ڞ���-5��<�(�i��.�ϥ�߈���I ��lZ��F���b?~�j�1%<�J9R��q�J5�E�ޢ� �'���Glo7�~��X�2zCݸR»\c&ȣQA�a���D��^�f���*�O8�O~T��N�rH��ن٢oV�k��zz[S?U���N�����o���Q�_a�U �����{��!��F�m%��o�U�YM;#KE�E����!�������== ��1���J�{�G[��l��U��M��h�A�=r5t��I`ޖ����	���GUO؟��|�ɀo:�I�QG��f�{	m0pO�{q@�o��T��mbRW��8�ӑ�&�ѯ۪�g��m�	���3���J���(�D�����%E�Q�'3'?������m3�s.@��R���ȄK�A�%�bx�Z�-����(9�����t��!�����7��c�]5PP�Nc�Y#<)ǔ���N��ct��}\Vc��p���up��G�>�֝��L8�}���m�pJ��p���fr��m)
o��+u�5k�5|�>p"Qb�ږ}�a<�V��د�'��ΐ���{�iI��؆�{���?�3p#T�^�!U��@Z�>�}�K! ��rS�T˙�8�9�j:C������Ӕ�V�haV1fhXq�Vǝ���j��%)p`��^��-�������RX����21�`^�����S���9�ՖW�S����;�\��:)�B(_�Ğ�ڎ�e�~��}R���a�"�����	�[qi���7p��l3�+�6��(�m��5�X�)o�&����)�\��L�-e	lW]t�~kzOI��s[��Rt/�ml9ޡ	օ�x�Q3�9j�)���'n�!$�k��p������vu��(���¢��d��v�!��>�l�1�JP��2�ѢhI���λ�^f��ƕv�R��E��x&ЂàҊ{~�U��]#5e�>�w�鍁9�aM}�@Mb�z�b���9�"3byCS@ds&���K�)��e[�ƙqf��}���}z+�v�[�;��#%�uC��4L��e[/�8�K3Z0���R��[�t�j��\�w��v+?��|�{�d�a�w�ڢ)�n��-T����T�u��ҹ���1�_���Hm�⊸R�'S����� �(QM8�l̖��a�l��6S��ϟu���-���N�,@פ��k�p�g���-�X�Y�7h=��rcWXiY����)�����C�IB6b?A���o[�~�;��o>E�Aj�P�kh$��b9�s��F��b{���p����.9i��<q�nV���N����ԙN�ѩD��@�Pǆ'=q��N�ωmF>�`���N�6�
��oB-=��V�U�H��t�_Џ0*��	�<��'��~��?Uk*��v6>�J�w*��e	/[�� �������6���떵�K�\��VY��HH�cƩ:��U�+�ur7(��}{�a�h�J\�^:����X1$��^p��憮n��-���a�Ý��8JH��kP֮>X�HV&��kL�"D�1��id����i�ؑ�T{�w��K�:I�)=Z	}���K/H��kڶ��t�A7���X:���5��ɻA;<�C����	%�������%ﵧ<L�D��y'q�X�����7#����1�(���{|�gy\�E��\P�����؞HH|�����{}/���y�T�)]�=�3�-���B_�fBd'p��u�	��T�oqW�'�&6�L��b��Gj�|7���h-�Lg�Le���Ns��֚�I95
Q�~~[�c�2Uy�M�a�m�P�������k~'��ͤR|�h|���v0�(\FwO �CD@a7O<3U�f��g͗�M	�Q�;'������5_��J�7��{�7V�{iդ��)�J�Dw�]�1���vj�:��!ERmt����������&����T�鉧�#���M]pЦ0�)]�h~�h|-2�ހ�f���x������F����(VK�J��Ȼ�@-�j73��%"�e٩7���
�v��텠O���CT��ƙ��E�² ��6���%Փ?�)B��>|��|��:�)I�\Ҽ1N(8���7�R�=��P�Դ3��,H �����p溕�|,�5�"(c�_�>��cuō��m(g>C�*�F!z�bd��7�4��#���-����@��4n���b:uA�T�?\/�Dge0/lt��`���vK�������HI�BYȧmw@w�q���t5�9U?~A�9���*��4����������(�,� |
�?3j&��_J'u���P�����3��~�+k9:�Q<+ϼB��#g��[������$�����ʲ���O�>�����d�v����PWn�3a!�$�Z��J��+#T7�fFvt~c�ɀ%�+��#�C&�ͪ'�(��qn1�@���Y�P���k��8f-�S7����I�PF�\��e���u߽q&��Wz���T}�t�?�������~�@�߹���ΰz>�$ˑVC�p���<�Y?��<���TCJ컟/��l?��ڤw[�IW<\}5s��k��
�|�|�[�s���}��z�	 [ܱ���Xl�E�~�z��9';`QD�O�8�p��?'t���g�_�	K�Qhx�۰׈rJ� 9�(�\{��C_�������n'�,k����\��A�.�	�9W�'��מqb>�{�u�[������)��_0	rF�`���e�yM��E�9����2�/���5K@��ʇ�N�5�'�5e�r�l+P^��W˿�v�"21~SC�e��ut2���nZµ�:4��0��`����������"��g�{�y��@k������
8�t�|��T%m�I�p3v��qT�A%���^+�3O
K,enϝ�8�����c���ϴ�t��/JC��$j���Mbd�ٚ����@��
ym� ��tt��U�ђw�>6��G���(���x�� �uFd�t�G)�uX��o$�"�aR�#F�p���_�۠-j��Z�������?�x�3�����{L/��Xjq\���F���=�/Ӓ��B�櫂��_B���xF�n����^�4Wz�����������-�:)}Ӑ��nPSL7[��������2��bc���b��5��54�T/���y2�p�3��myK�f��8n�`WSN+�֞����?�����A�J��aj��Z��<j�����'�]ʸ���&��S�y0Oo?x� >2g��Yz�D,� �It#t>UؠL-���_�xQ�����T��w�	���nhh+�)�	�e��Z�2TuH]=�0kFּ9�-��o+}����EC�Raא����Bl�M������
>Z=�ĸ��2�1��<a��|��` ���K����+L#�)<x5m���O���4�y�wai�k�.�d�/54#G3?�-�2��!o>��϶�}��;R�� _e��&���C���$�FC���� ������i���l7n���g�)��f�1�J��J$�c�m���@���9���6yX�V���'�#��5E}�ذX���(�,�P�Zm���Z�T"�Mg��G��)�x� 3n^�V�ǎ�2�8���n]�0��]=��Ks�=#>_;Q�Q5Wx�dnc��S#þ�k�B.UN=�&e�οl��p��cj��V/*���8Ca�P$#q���;T�#��2�]�6WE�蛑�-��M�|l���VF��m��O�u� �QMC��l�T�pr&v��=�h���ܠE%�DrM�VOm<���U������!��XU��%M���c�+����k'ġ��i�
��GU��F��T������B[M5�RWp꬘%Ъ�j�eC|vFT���^#����a�Y�M;Y�	R d��W��q+��إl���21e5��/k#[8�0I���!�N��}�A��A�^����0�w��z����E5�4������2���$S�^X�����OMG��wҵ<�.�;*���ǆ^i��L��5/��*ϱ�	Ч�.�Ͳ��	姠l�JJO�;ߔ����mW�������s�����<�RP	ҧ|�C�����'{�����&F���1�p�Ӛ���3��9h�〾q������ҽ߿����`M&�y<jX�ʜ�)"��b7�94��ɳL���㈩���q�ʺ	� ��dR�N�g�ˍ�9Uo#�O5a͂�j�J&U�K-=�/:Ѭt�=�:V	fr�>��5m�#oV���~�F�p62�g-�n�$����-��FSE��',���^��g�K/7�F�6j�3�� �(m&j�f�^m�jҷ��f�˛M�G���r! 	]&EC���'Um�O�qK�vҞ/�o Аsϊj��)�J�'��}�'�d���^�>�qM���Q�?=����w�_�G���p�^�Oo�4^������Q��4`�Z��k��T�w�A�R�Es�*4	ѓ�.�ZYlu�����]��BrW�Ϳ����2vԖ�é��"�����M6*�������8-
-ey�bi%�*n��~9�7_
P� 2��ؽ���%�"�u������/�g	
�TG,��	2%ە������_5��ж��������zc4?+�i�xl<���VR�[2�xy�|{v>��1+�y���̰����"5�?|b-T�U�'b&SKq�O×�H��R	-��Y�r:4����u��]́1Gϗo[,g[jo�&�+~�ˤWP� u�b	d��j4�t�Zu�n�GQ��!y�h��O%�)UB�7�3#CG�V��dv����\�+զ%d1p4�>r|:��?w�՗&����4D֑�Wd���C#%w/eA���ց;[��(��؇6���.����u<���i�+j#���fذu�R�v��}���^�9�RZm��k��WN�m{�n�0�e�T��J���~Б�_�^k(2
�:t3<P>����+�Rs�̴F*�#��*x��0�ꡘ���>��'K���L�����������_>��j��	/�Y�T���n�X��]��XmJ�����T�B`�{�O#0����d���#� ��{mg�ݪݸC:�hf�r��Ү�uv1�2���&�O-F�3)��"c�@^��kI�s�B�a�?z8�_��"d�0���͖{^N��ޠ��g� �ߗ�ѣ���4oE`�����pЧE�y�2R6��`3���� ����@�w"�b-�&���#"wg��׶W"S��j�5;�R"d�}`XL	�P>��m^25�4&1�ʇ��+!�>d@�2���$Y�Zٸ0ЦQMvh���}�Q�R9m�G�6kr�M���fj	'z���eCu�_ �����z�p6#���#f�����q����h����a�t��Z_�D`�
��)�"e[`ȿGs`����5�4��G��u�;L�
�U�5*eN��k����D��ݛ��V��b���c;W�#��P$�~k�6&z�}eh�`aT�Y2�~"��3Cub�$��9�j�RM��ǌ���̀|GD��!C[��W�*�i!��9#.�N���c�������u�t>!��m(_ls'j�Cn�G�������^a�\�(q�I���kV�R��c�*fBǌ̨��`��R7�jQ[|�1;g$F�� ��<�x���Ν'!���f�hzn�
���q��J�S�'q�ć�o��mݔ�	�g����|n�z�hӦ��?���.�Cf�D�v���r�)gj���a��֦Z�G�m"���*�>37�̀��v�s�zZ�^��2�ϔ6z�Q������;wpr�j\�l�2 A��]��rV"hj,5q�RSdZK����<�ϖ�/�ͦF�y�g�����%A�',����p3S
070v\��ga���%�lҢ3>&�V�$�+��Jw,��������ձ~^dr�U�#�5�e6�|�����i/)�?M�'2I� �l��n���DB�񹴚�檒�M��N����o咢f�f�Bŏ�,!��p9=0�E1/_�}��1 ��k>gh*�eun���#H�\��ٿ����/���y��@G_o��y�M�$��T�}bq?�lBy���_X���C�C���K="�6�~�� گ����c���s�[�%� �+Pԡ#��YF۠�WB�������
��Dϧ3���By�+iԢ�r�_8�w��h��G� �Ⓛ�t`�,�&�}�N�c�J(��m�'��g�['�->P�{�S ���2���Rb���p�&6p��<�\�BR�8|㊀q��|�.�[��'��<��'0S��C2N> ���~�D/�Z<Z�NY��-��K2��ǂ��{�\�D�w�H=_�v߆a�RD'@3�^73XV��/|�K3�q��kY��{8��ܹ�[�K�~V�N���:���_!��`S$�n�\;,�F�����G��"$;|Wz�9����l���%�9�"�ٗź|G��(��qR�BPkH�e�h�(|��ә�$�7����
���~*U���{L�<+^��=H"�����=$�li��~����9��z�Nl��o�X� T���D[Rv�,u6�]��2�kC�(�]Q�,�"��	*S�H�%{��=����@�t�Rf<q:iE��z9�y��"Wc��U ��w�@�o���0�u(<�xL���1CkG�F^K��C���e>,BK{&��h@�!.CȺۯw\S��/�l|�-��_+T�����#��x�u ��K��ɓ�O��Ѐ���߄+3k�c)-0��v���T=�����j�T�[V@��y�0�����cw;hRDUT��wo`#��)��������/
�l2�Ϊz�e@e��0��x�H������Ef��O�	��;� �V�:�ޗ)�cH�<K|V�Z�X��(��T7F���@X���LQ�
�$�G�%��fUҌR�(�����E��r@]�p7��g��Oa�E�2�"��(��b��1��l:���< g���E�2�pmĺ�2�SɝW�R\�μ*�d*o���ˍ���
Gyل�(�YiM���_�W���8�A��J�i<��V����ᵄ"��79�uݔ�f��Ǘ�}�|Gwiu,��0{Z�a!��igR���36���,FU�,V��F7��
ZV.M��j��Y���)$���q�tu<͓�d��
y�4{�)�劝ӥ�� ��Ɋ0������E�׍� w�Da�
A���.5ɢ�.��h�����g�S4T�
��7�T��b��G#��
�E�I`2Q��L�م,lD(DE<��6K�uP-���k�h��~wr���H�Y����Ȗ͡c����My2�$	�P�Zc�<��pw�SgG}�>���MR4�6���l*�*�Q���T�%��|U��b@����̛_ BŽæ�6��i�<��|-bC��B�4�NXOgTp�9�d�'�!�����r����9�2���,y�,Iք��M���J�bb0O��5RyR���y2�@���❑�gQ1����N.|,Se�ȧ�S4�$�����گ&��\a�U4o
�#�~�Ɗ���x�=�Su���h�}̎%)���e��{�3��;�V���8��߃�8��n����ƂS��+>�}�iRbUH�9וtt$H��C�R��6�|S��J��9�hT�M��W��ޠG�v�����cr�/X袨]Ȯya'c���Љ�<t��^�
�����ӯ��5���K��e6�H�f�h&�pL[�`��׌�]xi���7D㩞��l�\��3���]�������b� 鋀��t�:��F#�XC���G{EUCfҩ��cD��e���%�Q�"����PUV�P�
�e��T�wd��04*��EU�Y])�t�=�bζ
���|�C��szZZ`jc#�yC�漰�`��M��Ť"����K<�Q��W�gb.E�����i]:EÛ�wbXs���B���v��Te��`�͝y���r_�w�KfO*,���� ��]M�G[Un����^����×�Y�`oH���nη-Ue6N�k��MX�Hy�%}9�~��M3�<ko$V�#):��$;��ɤ�>G�r2w��g���F����J�4%���s5N7���"��4d"�Ʈ~4F M�W|�ܳ����;&��D��}A"�J���.���,?�`� C��L/�#>$�=��,u��s�
��f晎�ܺ�ZZ;F�����@*��)�3=��Q������i�Ga��N��C��يu�<�Í^q�YD���5:؂�+[�u���/�֕5"��	�	8��2ir*Vc��>\��)�T��;�n�ki3��f�Q�GU'�%����V�J��0�(�6�"�=7����Z�R^�Y�%�Y�㖢��&�����t��Z'��ͭ:d��U9�;(�4:�W.����Ѵ�q�]o��`�Ѝ^	�@Goʲ 3�2�Qў�B�%u�2����TC��"�6�/���%ж������'햓"���;�femgj��$�C���]w�����'��E7Gҏ��=�a�Dhu������W����`���(�~���.f���ԓ;ҎŃ��,[/Ա��_� �j�A�9��ؼ��7O��\+)6
M_�
�p,�2k��	3ĥv����D��,<h�P��X+4���$_��`ӲI~�5������{�v:"�C��֛�o��j�Ϗ!���'��f�V�b߁�n@�Y��i�~�U}�ُ��v���\)�-s��9T�VTZ`	�xJ�0W[@E U�?jP[���gDI	O���o0���K�% F�Ժ�=�)TG�Gl>7����!���kk�����%���H=���|��;�����3���1����<o4\�H+�*�z4c��Ί�܉ j�E���RI�u`<�>r���gZ��Y�{�#��lV��_o�Z�B�O���F��6l�.5#BI��Y�?P��rr���*S�K�B+|{��c��豍������o3��6~z�u��?A�ܻ�떒����Ya��H���"�3NLh����'"�s&e�0'd§7D67��<��
&yJ��P��Bէ�\3]d&W�RČ`T{�=x^�ͣ�' �!f�/G�ڙ6h6<�� 64e$&y�K�Ed��c�L��.h2�fc#p?Y
?o`��0P�S�*�����m��Z ӡ6�*�zZ�?~�7U-��ߪ��,����V��ukyl�v�d����8�aQI(��4�K5'=�)+b�>#��q����T��w�i8�K;;�Ġ�W�4/>�8v���ԅ!x��~�d�u�/{��էa�m��m�X8�@u�����K���Z Go���x���Bٓ��S�HZk����:�e�R*�jǼ3$갊(M��?�[K긋�SѨ%�.��	���2���h.�˨o�+3h�X�OJ>�!c_�������4�|�:NL-M�P�Y�~xc��N�ˮ��}��O��rus%��ŦlIlLn���Pm0�+��"1��d�[:�j�Ұ@\ne��#d��(�����O,3?�.�X+]�a�E��<���D'Dþ�'�j)�^�,_��#�t(��2cY��B����;�'�>.�����2կsR�&{A��{;&�<(e���=�vZ���	>l��b_���'c̼����C��^� v���v�k�[��������6�hm�=d6¡��EF��2����՞�T	�X��ڙ%	5揲p��7�0���X�^$T��s����W��'�r�+�+�@�<o/_��dɬ{�.z�z���C��.���X�Ŕ�d�\�Ѥ���b�ӈ)��7�Q]n��S�}% ��7�.�z��ҹq1�Dr�����m8M��C~߾MX1�o��,Ub�)�Cpp�ti;,�YF� ����UL�$}�s�ìTz���^�B��Dl�Y<z ���u�V��3��1�O3�s��<�PWN�%9s{�ф�0M7Z gy��Qp/ `*��H)�_�e�k��Di�_H�9p��|�Cn�%�ڧ�p�D|H�$���2X�2<)��?�e������2��ՀG��ptxC=�m�EADU�R��)��+��?ie��Zƃ�&AA;T�p5*��g[1����$���p*^��-e��l-��U�+�n+􌗧�7�ٗ���]� M��TV��f�HFj�"�?/v��hMDPj�&�B.<����_��f�7c5 u'�{9K���� [%ox��fy�r/C���
��vK�{j��i�߸vdW49J��Fς���!(4��9���I�O�{�b�1.|���h<vՊW�A��
�S
�e+��(џu�� �����sǅR@~��ci.�Ꜯ��ۉt�q"���ºY?��[h"���@��	��b�8�<�܌��m�0��#�1��m��/b���ֈKI�C��τ�g�������!���ټXa��wg�����!s,�a�1����@��w0�D����o�s��v�rF,�I��qxYО٘etG��9'7�	����hq�8�(���8:����W��;���
�4��̛�D�K��Vr�#��n��:�=WA�e�K����Y�{E�Ƒ$���ĺF�p�l\�.�D�uq/r���qc�6���m��`2���<5W!�A�P�Sw�8�����wSt��L��	��*ە������m��6id��:�`���+��jݪ�nW��ga�	��h8`��k�_�0����
3B����k������5+tZ�G=�C�Bo�+k��:��%S�#��:^j\c�%���[�T�=��T	�6�o�j��	6:RFaU�M�ړ�N��A��SJ�٣�h幕[x��������mht�[1�T��@��2�_Q[1V=TTm�~�V�R��M�Ɓ��A�m��#��t��@��v�9�Q��<b%�%���@��>h.t���HZ�A��0��_�$�}�؎��|��G5�*���::�lokB�?Ì���C�A��MLs޸���;�Iml֠/�-��!�[O
��w1�{��Z����:��y1pwW7Xx4;����2��'!�Y���q��B�6���L��ez�:�E-��'�1�tT��y`��'��vo�,H������7����8D|wfc�mD0���'&������:��d82E�b'���R^�_z(�N�m&|`����{পy��L<p���g,;�Pz��jCL��2���H�`MOh��eyAb�=A	�β���RAG��C$o�K~b���%&g�:Ƽ�^��{�>��8�v���%���h)�;=E�%O���i�1�r���Iޔw��mt�'=��k(�����t��T
������e��ib�i�����9k��d��&�x�A�	���j?�0��}��������ʆ�|R�a�I��#)#�����A)k�v��@,��6�-\\d�T<��e?�����Wgf�jn�r;*
^�u+h��}��m
:�r���M�<�6A���sj_��L��p�X��i-8�G<-��!vx�[\f�ͬ$即�q���DȮ���<�m���#j��~I=W���F&Ó�u�8n�6�� I�s=".nu��a�~iʅ��c�m���;N�Wb6�HbT^*��	��n�f�l�R^%Xf� =(칿�Ę&6<&ƶVdq�:X|�L{��T��ܡ�u\,i���!s�x�>Z�u���nӤFo5oQ((�6��ǽӥn���X�]��~���1Oߖ�.A��UmG�P��Ҩs>dV]��,��v p��b�� Pm���4�٭3�:0}#=F��0JE�J
J���0?8{�h�o��1���*+rz��n�_Fz�#�R�
�J4��  -J0�@-]i�Z�ط�I���;�M�S��_M�*��g�����r���N���9�G�j�D����P#FN�N�>ҤTi�JO�a�I2u�O1��L쑌�P�c;�##����JjMث|(�BRK���	���
v#�'�73R�y�P��~�]A����hb��Ǖ�[�"p����>�ݕL�������mw2[��a;_�I��O�Ϫ� g2!oG?����INX�*]{ɋ�M4%���Ul�^��ۖ�TK�J��Q��-�"o�+ӫ�ap��6����Ӭ���1+��$��!��r�`��f�f�����+@�-��a��/���D�t6�U3K��0m��!(��	Nr�z��Jl��ݾvL �γ��}k� �|:Q�WT���u3��DMX_�`=q����.�!C�x�����ފ��	���T3��2_��-6)?���?����mX�[��?�;��U}���;����5'F�vV]&� &��Tψ��G������Z��
��
8D/�0��-�(1�8��8�Y������~��ۅ~��˵S�3O��[�hr�G����h>@ڇ,�2[�yP���L*XU��nFAiL�P\Ϧ�j�����H.�E�޹��@�n(�Q��kS�����fS0�$0�q����ʿ([�}�Lŋ� T�k2�c�d���i��+qx���i��	�q�*F����.����"0��xox(�;~#y�{F�mܺ����ǈo�C����H��*����/Qd9��w�="	�z��|���B���r3��_�	$nT�:D?I��4� n-E���c����t�1�����<E�~��%F�J�Vw�߼��~+�H�m��|ı'�a�X����M.̒�bbSk����?�Xڙ��lx�[@�԰�ãHNf,�������=~�����hoI%��7�� 4��c-�E�d+�*X�B�3��(��q�7���
ѯ>p�eW��	>�y;��A�Ğ�S���7�4*d`�ܵKu��39D�g/�ɰ�A�!}��z����K=DXP�_��	�- 
�3)7�rqg��O�3�G������bk�j�Y����J��%�D�-�'�43�jJ�����˥v87���)m����2g�c�ot��v�x��j L�'�ug���nX�AⲀ�j(󼆶݉��Cع޻�y�%����O����"Z9�Mµ�:��;�S�%#ܙc:��0rt�O�i|_��)�!z��.�RwT�$)"(� aա���*N���V��zL`���(��S7�Xf�n�v�b5��t%�M>X��g̖��-,��Z����..��E�����"A嘣MG�{`��YF1�RnK�W�P�C�ʟ���Al�k�}�xϷ^��ExF����G@DT�`;�����6W�S"�F5���~AP�?Z�=0��Q�U�~��z`I�M��a�a�&�@h�]Cݨ�8!R�1���\|�ۆ���*��_?OH������Ej�����U����t�&���\�8��@�Q[J�3f���'	7�7 xe�����eF���ݞ��!%QGR����8P���\��'�SR�o��F�eȓo�ُ1�a�B/�%�XA^2+TH��-NDɝ�<fD�(�@��L���Un�ʈ�|f���ʗ�e�,\6v|c"ceD�o��w�+h���W�+ɥpn���ƨ�6��P�/��m�U>���mn1��ݽg���A�<�S��l7X<�ћ5�Q2�AL0��ҩ�[y�?E?���T�C
˴_QL�v�\'����໐���Ni_�I�/�V60I���e�r�h�>o�g����#5qk���s�x�):�O��F�j���pӗ�9����N�ϑ���j�3�*Һڤ|�ݼimm�T�>Eم>����G�<��6`4x���i�:U}�g��D��ȃ�M�ň?�'���@�E��r�Z����f��]�k8֕�$��^�]�X n�޳��KL���+,�Zܫ��7���cGqu��0;���Hz<�B�&��Ǡ�g�������	�������h�9�fE�:�i)�µ�~�����i�U��;�NGp�p�H�m����3�|mD�F�ʘ��>�n��Ϻ�Qޙik���k�MfF��-��	�"Pe����gĠU����B� {'Vtb��>��u":�8�1k�����K�Tr��>���������d���?V�士�;�<͓z��U<��(��׊��wjA���_��%�1	^A�G�*�P	嚦����S�+��lP���G�i/�,��(�8������4H�Ə���,�Wu�l{��d���&�պ5#x���� ��=�̜iǍ[Q�j����b�z:D�F�k��<2�$te�i�F��_���rk�r�f0�697;�B�\R�^� �a�ߑ�/}�=O�,8[f��ȗ��D;B/a���x��sy����Z�aK`T�W��fŪCN!4|W��%;�kD0�����ۀ`P����Y&��a��Qopk4&�eJ�FwgA����� ge6���U�C�/��8�*��4}�n�ڝ/l7��R�V���x��|��r'���<��{iM��kM~:�Ƈ�������&��3��P{,?G�8K�R������! n7���kMU�
��j.�e*l".�0��T�~1��pk�W��Ȅ�u��~`��ƒ�%��E�#���L�@ȑrG	A�>]"[����V��2�(*~?=��@��XxqF����V��C2xAɝ� g:�s	6�g9��K
1K�P�+�mPU2��B��=�6��r��1�sO$�%i&W��8�R�cO�d%\�(��@ܦ��'�m����5p��i��%�לr�H��5���ѦluO�a��A@Q�C��1�k}��qCv�e��
��rW�r@$����{����yd�L d�q#�4mڳcm4Ahb�Ә�c�p���\RmT�8�+^�c@r��9�C��gĆ
�L��5�~��z�Lu��#<X�x|IT�����<��?�?B\��D@~ԯ6h��G2 Ky�mz�5&�+��>��F�v�a�Yc��/^��8)�b"С���RX��k����)4��ÓS/b���˕�g��{����P'�/v�=�h27W'�U�1������N����Uk����~��Ȍ��cY8�
��������S-��U��g�t�CO�z�r�7�p�#O]�2�m;%��Ҧ���E�%��ZC| �]�$t������
B�F���^� A�Ry�
x�1ɷ`\&�x��d2�� Q� ��H2έsy���E;�H,I"������|��l\��Tڦ XW£.t����f�TKF&u�K�TU��>{�����&-l��z����6�	�Ϭ[��ˍ���
�#y�-�83D���y�L�8�z׆�JlU��~������7�O�����E��(,"*���z�c
i��~B�ɳl��N�:\/*�!X  �t���I�[܉,;9aN��r%9��+\cS��R�˧��)�c�������5��Q�(�=i���ɌUa�x�߉V�2PN{����Av���O�Հ�pK�=�dpj�	��Ӿ���Z��a��ٽ�1r{�F�,�y'�jȆ0j�D��Ko_�mCs+�&�^p`'�y����V��$��z:2=���$���`��S]�K�<|T����T��ye|Z7�4�A�nW7��ݜ�8�\]�!Xz#�qI�tۍ����2u���?�@�]�Ƒ+.�<�\S�U���j���y-�x�o�(����j��([Q�GW��U%�0_��	K`���H�EW���y�XTG�4�_�,٨�4�<oTI����w�s���R ���K[X��A�,1���@:pa:�3�Y�OK���ԟ.�,��BfWP�*G�u��7�Z ^2I�,���}ƕ^��<���C$״N�G��y�Jn���D;
��(�NDLQ�ZC�j8���g<��e�<j֪hHpڅ-ׁ��jA�{\�=$7��s�jV�k_�?s%� �u����Z>�~�H�l��C�'�sڷ�M����&��=�|�Fx�u��w�,�Ӆ���=��E�i�u_,|�����W[����r}_�b�9}�l�p�2���fM�5u�)�tᨇ��$���&�f�8s�X���_ܛ�8�:�1�s �O��0<]}J|��{��9,��i�d�h����k���Q	��H������z@�T&!h����	ZWiH�wؐ�w` ��r�p�� :�/�hJr}�N���{������</��C՗��{�1R�����7�GﺪL�h^ Z@�Z����#�hh�K�Ȕ[��[v��q-,����~;K��ZR.�g����\l����ޑ݁ۘ*p��<��y���H"�}<��r0��C�)�]�/�_����6?4�h��G;��(��6t}\<�f�"3��]H���9�;#{&8%t�F�]/BZ�;���%�*B��a;sT�^,'>O���g	�n��}B��(��n��$�˾���8޷9�c�8�|HK���zuC�;zCsE���3��Cu5�!���I�����/���ΓWi���F임"�e��ت?�Z?#����$Y{��2n����]=['��AB�8v��q}�"l���lb���e��/���Gk+ʄT �8o캁��͍!� ]'����n�(����Q�* T���\р�/��p	��	r�˕�d\ @�_��JzX��hK'R��O�R�讧��d!V̞Yp������ѳ����oyj.Ӡ9���6�g�7�H5�pE��^!�xAf��lK��͔ꑱE� ���i]t't�/;3�㿷�Y�9"(�S�i׿$��s?t��n�~=	7�Z�O;՘]�����ڏV+=�B�~@�q�.�9 �y9�ԘkIw��ƌ�x����
ubm������$������}�#w$���� 	
2���\�b��'v��v6��S�	���c��V?T��Hx*���VB��e[�=j�hݛ�͕�%|�PX|�J���7	��׉?I�xbg��Ho�&��n��T\#7��AU@[��(ڃ_�ų�ڶ�7�	�������~B$U��Y̺�5�ͅ�&ޜ�&&�Cji>ֈ_�����{�6� '|��GQ,9'&��R&�C���zDJ$YBS��;wq`�j��]\�5�D�#yR�Mr���v��0(��f����U�,1L������������l��_�B_�?Z�c��T"S@�Q�e��X��@�_�����0�᪎kQ�ݸ‫�0A�z�n�����x2�IJ�b����`�����%�8�-�K�ߟ�	��7��(�D1��h���k�1�+R�3��h�C����J�s_eɣ���=��@���<�Su��[_l礌�s��I�J��y�W��0;�L20�R�2Vw��n��+�D�~ϡ��ץ��{O���e�]�F��n��+���!�]y�e�`"8>(�h��:���E��LT�mK�_`򰲦�|rP��������[�YJ���mP��ϓA�U�N�MG�-˫S��
pU��Q��U�$;2_��8�w�#Tk�Ѕ���s�k$� �-��8%���i_�C�A�-�F�BgF`�3�`p�@���*���'�^���X�,���א��sm�2q�+�D|�4=�*7�{��H�#���t��{�vE�I����)�%.��A��
*W���l�nS��k��4�%�]ƫ�\�0�����D!U9�R�2Ꝫ5�>����w��s��;�l���X�&Q{",8���/�``�L�� ���Ҝ�T�%���ۻ=x���A'9.֦ W�>�7�Yo�w�S�y�ܝA�̦���-Ly���4��&*����M�뜈���c==��	��9/A�6�չy���RR���������'�T�������@���I�B]v��"%�I�/�k��)q<jN*��n%.V|����q1*��m������b7�U�pC���X����)T`7 Lv._R<���r���<ٟ���h�.����g�x�Ӝ��%��V�ި\N.7��ivޕBB�ԉ�_&`�	Bu���9`����Ѓö �uiP�=uE��'�u ��XG=��V2$J��|���M�@ǂ�#���ތ5�V{b��h�Dp&��x{.��*�.(E�*^�匱�B�a�C�z;����5���$Y�fԡ��;��ag�>-6�mC�ڱD�*un��)/|+Rÿ�Y��h�Qg�t���+D���e�\�J\o��RS�WZ��E�4y��@��E+�M{�Meȯ��q�Q�P�h��Wfۿ+e�N
+T�'C7a�UÞ��p꿁j�+�.z\v��i3V��s�-�hE������|�x2��N����m��k�e��LU#Mq��hv��c�����$S�n8���>e�0�=���d$ �S|B�IMX� ���"�"�$b@I���4��U$�m�W{tXY/���MΈ~H��K�0zD ��ů0Jc�ؑЧ�$�%e��[^�j�hLY���#�� ���L:�uZR�e���	� wa����m�T��Zŷ&��rDF���=��r�Y��$��"��
��-s!u�R���z��(�@�������?�~0ME{���/���F��A恶����H����~�.yΗ�oJɰ���G6����@_�YH�o���*&U�V���\?e;��x��ia�eI��RnGX�wA�A<��ހ����(1�⸺Ԩh��>ڻ|'�����k�<,˙��# ���E����š��˩��y�1^�dh<O��s+{p��*��Lb��&��5�8h�\Xo�m,��n�
���Vv ޚ�T��פ��㰼������O�[�����t�D�Cvi�����
��:.�~S?TWc�<+�1}XV/�CB���n������(�^/	�FZ�3��l0��?�%Y+C�O�!`%��o<8iqdQ����Sk+@�"��x�  ��k�����`zE*� ��u{��,q��y{�	C������%�j��r>М�Ò"�������(����%��:@/�ҷ(�|dHu�f��e4��N�������|��b���풆4i�rg0���!�
A`)[���Kcܵ�@������Xx�T�_��]� )Z˼�L�+��R+u'ɒ�$��$���ä+R8�u]w��i�n�%�]9{P�����5�FN8I��e#��<�����Љ'F��\+J;�� �{9�ܺ��(+#���Br�k���9��r>��v�B�"�f� V�a�N�m��u%8(��w&7���T�o�7�$)�,��:"��b���B�'������k����M\b����y�(�O���bs�s7�9psH�Ȇ�����ì�4�	!���G���0��a�o��?�̂��X}:�VF�[�w����w��\3���K�'����K�>�8xlHN�&	\<WI~C:��hy�f�P=�tQ\���[R�4\����z{�\�[��5���)��>M��(5@�-�NRO�I6�˩:j��X~�T,�?��EQ��x	#���@vϢ����Ⲓ$|�(
��+��^�4ѥ�h��
���)����Fܝ�8
g�)��<D�ՙ�f��g�=~����^/T�C������|�:�2��.8܍�Q��01��_��W0�ط�	�$�Y��PR����AI0N\ר��} �<���G7�S�Y?Yy�B(��%��X�����K�"�>�|��w��	i�d�Z8k�l.T/�ײ2kX�<��Xy�����h��N�?22�sL,;jT;��X��dQǳ�~̺��=}����TS[t�P)�u��k�{�Q����͔��I��I)��8��E�v��� �8k��ކ��@z!q��N�З�PӐ�Y?������j(��`@Ytʉg!��Śq��*L�K����o(a�2�GH�W��D���>V�)#����~��10�8�V{�0���*�Y��c��4�K�g���V�e�{/;^�)h�������?'k��"�?�� �Cw�*�u	r��8_�����H���<Y���D'�N+5HJ���<�,E3���V��}D�[oܿ_���Rd>3����B ۙ��u��T��k;zWL�F��X�Oj����p������BZ�d�qK"A`��[fsV�1�P���VDl���vc}��3?���!p��>Wa{I΃.�PQ>�tT�R�؍`�ʅ>�t���ߚ.�1p�<�5�%�ܴ��_�F�E�b<�J�NH6/;��3��Uo��}��!� ��(����v7h���
�&��e{'��(L��
��l(�Њ�� P�m�İ�j-e�i D�r�ջ�jm�z��Ս#���=0T�ݧ�񑯃$M�ƕ����`G[�����F^�=���S�d�6��=��DG>���'���F�HXgwF�i�Kb�/Ob�zr����w7T�Ѹ>sk���N��U�8��a�v�l��Ƹ��烊��yC>4����u��²z̏K@�P{�_��Zv�A��] �`+R�b����=�%�N����!�<��1�7����R���Ù�?H��p�#���Է��]�n��;7q�[�􍦄A�l5����J<��0������c���!ϙh|����F�q�9H˲U�L7m�֡Y��R�a�~�qw�:�u��n\�Wb�S������'��y���v����$�	]%���2}?ܮ��W�J9z�.M��8=۷$�V��Y�����Wn�(�S��֏��̎�U ��4��?�>&6�Lα���a�Tu���42�rJKn{[?YJ��>~=��v�n��J�����i^�ș͘%m�Ȅ����Z�J� �bY�΋��-ʭ0ʧ:����r�h�9���9zp#�^�df>H����2�$��>� 6�,��2��A�p⼞_嫙�H��?8�/�n�ᆩ����oA.e#��Ű�l�;��2-��䚜]D�S�����#m�/�Pe)<�d��k9f���7��ު����}�i��v~-���%S�h��,a�8J��υm8Wc�n)���xh��\�O_���F3�,C������jO�c�]a��'=���H�Y�Q����#^��[�P[:��M_��hT�@ʋ,��K�<Dv���Ui�~�O'��W��6Z�'������������j��`��FȓVl���q �� '�Y�S�5�t����^�P<���Č��%)�	�+4.�+�k�[|��d��05h�~�a�r���pf7&g� s���[�;;���dΈY��yDR�+��t'�@�"�e+PWcC�/�S�ݕfo�G�-wC�M���v�,���g0��ᩑ\���Ñ���/��=�����'�F��V���#�\>����j�'�)�B;�M�k�ύ����i�o6�}I,f5t{�c+v������V�V|���A��$�P���1zg�s�'�#k�ׁ����~)$���T�$���󢲛^�:��v��1j��9�Vi,@s�OTR;�2�j�!m�c��\����g
S.��o�t~G��ߪc���ȋ�"�;��lN4�����?����SM+�~��c\k��cf ��ģ��bI7v^�T��C�'o8Dx��ǒ.��1�gqe9�%6	�(|�?���?�a���\��!�ٯ�N�.�	\�f�!�n��i�dӘz+�X���V��Xit�0�'�F2?�غ�b�WP+�o&�܊�����[K�z��F(Y�#��:T��<d�^-�:u��	��J��0� �� ��Z֙h�ָ�W�vIgrm�*m=�1���q6��R�:���J�Bz�oτ���q��5�3�g�(����׸�.+�?Z_��X8 %_�G�Y��kXz.H�q�3�3�����K�����'/�^R�`�8��x�s�ALh�i��/u���	I��~�j�۫J6jN���_��H��H�5k3�d�q����`�d�/[����(��8�jc+4�ж�H�w��,$"*���� �h��;ܾ��l�Ws�G9Ѵw�0�^f���noMu|D���p�n4��bh�&���՝*4";fE��lkl�o�8�
���,i����W�D�ȋbm?��	D1�/�W�u��C��n9~�_vi������/!��O�?$��Ձ{������u�|�Y�
�?�R��n�vǉɒ,�E��
7#{/E��W8���Hw)� �+8�Ro}$`)�O���bz���� A@Q	�O�(ZH���0��ܐ��-0\>�W��?E�{��pe�t�4'%$i�^��j�B�-��oQOS�o*��$کKZ��y};���>Nz����w��ΒG�m����Τ� ~��[,gEth�A�d=I�Ι �,���_�A��0��_C���xéޫi��SH��\Nʴ�`��������f:�c������2��˞	9J0���N�::ZH��X�I��Lߵ~��[���Bk�r�9)y3#��*�x��YײC I�-��N���mg�kM��Vq!hL �v��LA�B�lTn�
˭	�~��y�]�4�E[�:d`��y��7m��i�*���{q%�aA��&tM������2��zJ����0O�!`���a����D�4l�Kݟ��NxD�����G ���+�[�����^��O��w��og����z G/$G��ra_I��j
��I���&#��*�e2{��p��M��}=���y�ܗ�k�QvO�kZ���d�!�� �>����#�R7�5�]��z٠¤�����޺����HB��:����V�L=������鵆6D�pR�SS�UV�f�Ģ	N��C�B�/�O�N�pRFZ�/�r�owU��${STz�"@ ������X��6���P{��kuF�J[�������
�N}b0;Ӝ4M�#`�V�}�ڣ�&�Ϙ
�j3�*&�"@���4�.L���;qq��i��e�R��N�}}O������ �]�uUY[�I]��W>�3��V�h.!�ݧ�� �E�X�L�E`!m��.����bf�U�a`R���C̳!�Zb	s�PO7]�}��D�����'`�a��٪�l#ƈ  �AX�L����ܲ�u�)l��q�``;v�>{A���߸��Y�蘤��fEW�<|<4���z����X)��Z���W��:]KR�!�e7f��yc̺�g>,Di���<�0lc@�\�ɬ�+.�bu�����g�q6nHͨz�ڒ6j�c(3�c�$t�s��{��xH_�T�������B�_�&�u�ޗE���]51����Y�G���C��%��(ߴ�ѣf��Xԣ������,6����j�%�H�U#���?"e!d���=԰��"�?R���>���#�s���C��WM�P木]��:��*4�2�!;�p���S�p�p�U�p�z�=�� ?�s����6O�.|�c�Ń��]K"�>�Bz
��YT�פ��N�c���&*���V�T1���k�1FN�}
uzx1��cKք�΄�����33�/�8�E�\� ��ݢ�l/�s���\gj�ހZU��c�3A7�g�G�v��m9�oZW(�铼޷��/�{�'�����J���-��Rr#>Ba���s�?$COs��[����Q-�zBsS7Mߜ��I(�P딓H��;F��3@�Oq$$88���xᗌM{S��y�<�q��	�^��&=��g\�ﳽC����чh"����$����Y��@�)�>r]!��>�4�/;TM�hÛ2�oS��UA��g��	�����8�N��L;�j{�&j��s�Lp�,���#7z�j�QC�|�ޱ3!�c�X5������(m�^�m\�UcB:X��5���<�5�8���q5���mx'�-,�h��s�庴
^o��z
�|���)���F��^9zi��Lb�?|�x"�����b�o�ȸ|�$��=9���F`��%�MU*m�wF�~VA�uꡕ���1Bn��hcy�m�8ܝނ��u!�5-�2���4(xrM8�h��� ���H�5��Wl�h~zLK�R����O\����Ca���S�	ǝ\,Ba�
�b���� ڤ�7Кe¹'@?e��p�'%������x�ܛ�*j�P�A�����ÿ�����eq��0�)ɆgO�\��N����>�S��Jn�l��N�~	�������OT�
>*Pr���k�?�<C��o1=�I-���ߔ��'vֿ)�R�n.�̕��3|"�k�M����+?֑�`���d�A��$>g��/�������HH�9�哬�3
����=��EC_���,D�'�*�xm.!i���$.q��:���9�o�˷&�-.�8d�K�n/� �����3��V��.2���v�i������l�#˙����Q@_����!����2�DS(�G(3�h��p8Z�)SbK�X�Ě�<׀e_�'q��A�ݹ��%m��sF�
k��亭Ze��_Q3J�����l��ְ�X~��^��.���ês1�qx&b8* ����g�AR�T��*����^�|�HF���8���*�����+���G?	0�{�(�w&�/��w�� px�b�ґ��t�_tR���5�Sy*�q��7�Ń�{`�(�j��KV]�sp���4��K��6�B`���j���{ɀD��}�[�<q���$����y�����GVg�6��z2��C�ҥ�T�8�!��������P��΄�m/Q�j�a�Y�,66���6rgW]�m���j`��.��锢��~/�{Hlv�X� I�I�S�@G� ��%L������ �,���c"7ږ�^+��\���WL�����u��>|���P���?���<��U�/Z�M�:Hx�^��W:�w��8�+Xo�E�H �:��|��ʈ6w��|�)���zv��!�n�@�CS�|-�D�R�>��٬潄�Q�g�r��o���9p�pp�P�v���u8z��Q�R�%�N��	�r�uQ���E���Ė!�h��C��	 �2_���#]���`�ܻe|k�ʼ�R��g�oN�Ce����A�e_la)��v������E���7E��Oz;�rA�,�~�4�/W��Ա�6,��Yh��ե
n�e���SѴn}���ҁFg=k�;o���5�+c��l	�tB�E�Ȋ�o�7e�l����FP^\Y4�f��_i����L��z�B�|��YL<��g�i�fwR�fW)*#�{�?�����������*@ݧI�(�����G��e�z�K�a�"���=���5`�
s����>�Q�]����?}0���6Xh5z�긷�bw��O��9������7{�<aq��>C�3mȽ�T�ݝRf������˩��&L��� ��lB�S��]�s����K�.BlLtF4��y�_)���^ �_d��n��~�4�O�ޅ�17UV�BGs�u�ȣ������O+a1z_m�|���uԠlj��^{�x���H׾U���������wF��x��2q!O�'�/�<�8tN:&ƅ��v���Y�%t��ߡbgy�:�W�"4�3Q��*�nۧI[漹����a�;5'?Pߗ��?���ㇵ�P̆�tҋɆ՞���E�`���hQd�^��i_=@w�5�Kz6e�w�7�α���h�� �_]�{R ݈�,j��(Q�E�>7��w��=.'�Ӭ�{=��.�BNxB@�tg���}�:^�f�	�f[1����U���psP��n�ն*m ;��C�r��I��� =��9Qn���ܰ��p �F��������=K._���r�,�8� �Қ`�iKJ�� �g�Nw:���n���e�m�¥��e�R��B��(��u(/�e��Nbp�ef��y�J�
#1$�A��H��� �U�w ��Q6lW�8f�Ч��{��3�-`[vGGN�-O'�*9����hG �L��Y�"&��_Jq�`��6� l�v����'����db	�6|�d�3�9ܷ2J���߷	 z��������C[�x���!�Vl�l$b�	�h���;��d$�䣡z���E��!��D�]Dv��Y�i-$ʐNj@�1��o��
"o��0H�!��/ѳ.,��	�o��.�y�fg�`^SȐ���b�n����j��EWY?6�8��h�+h�=�I��(@�聃S�ЍU��
}�C�EvšAt��g�w �uu�5Գ�n�����Ӧ�r&AX����A�쒓A6��{v�|������[��F��Յ��k�2�B�P �f&�ϯ;ω\}i���7ƥl/��R�$.1aJ��pI*c	ZVE����K9�u���������~Nk���s���
�~��8e�axzr[��E��Tޤ�8=�� ��}�1��I�4*�"-,nsk8qg9����!:G��d	�7���1@�;)�|�}N���Ԝ<TȪ���v����+kO������ �ҮY~5�f���QTdBH��pFN�r���NpڲT�ddm+�l%��颣O�Oe�p�o��߉��7t%����ǺG9[!!8�H(�^�ƪ*j�����[?ge� �`Ie�I~r��8���1e��	��鉕��.�p70{��+���(L�.�~+*p�C$0�r���\���ٳ��~�3�׫������P�}�x&a&�~Q:���N���SuǛ3��4��De8Z����y�:��Rq&�A�4v?�
�MK���_��+K� Y�nj�yޟ��6����D����~b��ŋ�%:"Gغ��;�=�R����������Q���E����s�"�a��V��B��j�XP59[sU%�~�g���=
ԥW�2Hf�'⅊M�W�$8��QC�xE�pM#N�)@��[Ea��"L��,N�4BP��u�I%�S�����cR�l�.h���Fn(4z�2#(����0Q%�:�a�@ׇo�F������g䒉�y�1'��nXWK��^G��2�bj��������rƤ$eg�+ɣ,ˈ!��T~�>�+o#��~�TKBV��ר]� E�&��4��O�$�xJ�6��B�:�8(�&]R��L맄��sj�rQ��/���D�����7��b��x�c���[�h��<MGh~�;f��?�{K_��aiPׂ� �m�_����VH@qyzv���ȜB~շ�v�}�>	�?X�͏�Y ���`����J�=�9%�5kdr�}x����)N'y�G�.����Kt�`��
����ݘ�s������/���\^J���5���gBj��M\��_Pꉾ�px��i�U9,Y��.��Q&n�iB��,���+ϵ�M�x��Bw�{��j�p�v�$�1��oH\�O��S���,p�Q��gp��^�,]I����i�����>�J?.�Ub��_��r�h9����iG��L�&���(�ތd�!��H�CfW%��L���->�O=L���k���RR%	�Hwi��2;����Ɩ�::ZZ������V�s������Ų��������rN� )w{��Y�u�~t1m�eO�+��K�͗�'����I<a�Ӄ�n�r]�����ŝ�"6/�&���N��9�໶�~���O^k�=����s6�K�l��E�z��r��q;���TxR1��Q�8�Dn�(�Tf�GFYT3�O\�KrT�ܩ���IڼrO��ֶ��H*3�\;��ɯq��v���[*a㬢����됗G��N���j�@���%]�`��\��O}�!œZb��c����xl�����&���∳���|�^u/�U1����u�;�*�m�
T�;���X3w�E�\,3G�'>C�a<�n�.�,�'�"�1�
�G0*�9d �zMi�6��R�/�G�}� uHe�P������ ᫨%й��]��@.�냧�m���=8��Fs�\f��+M�������:�c'(h�=����t9��ut���|U	 #�v�c��˨��v�qX����]/���p��yu����m��<.łZ_\�3Nv�ߑ�M�V���س��" v�4�
��ʹ��M�C��O����^	�gK��K�h�$xe*t���e�����مO���!��2����w�O~�X�> �PD�2�� �c&r7���5���+S��H�"�+~Ҥ�g�qw6(��_�=�G��]��>I����z�$����b4�����2�i��a��t,2���w�_�B+d0�8���7I�⌙ZR܎�����g����ܝtIѩ>�W�OY�|M�|h5�By��&$0;�G��L��[�`�L��\���b �t8���8��Am{��wf�?���L���%6�p��ڔ��Ժj���"�d�.���_R���機�؆4YW"�߻ш4�^q��ڰ[��X^��)9����:�|���@���fLL�(-���ȃ�J� ;k)���7u�}?�_h�2:ɘ��ԟ�W/���M�ö��A�t�jR��Nt���@r��]$�z�P�(�e��"����T���/"/S1t>�iu��$��up��W&s)CzS`��^8_ѐ�KQE������`��+���2aU���Qa���OR-v����|p�[W�̖!���aÜ`u�@�q���u���y��4�X������2;8�j����ȷx���z��C8=��B+��e8I��d|�u;���ބ��R�s��i�Z�|;����c($O0ʅ^>,E�r�i�{��ԭPp�:��;��[|�����k�8{L.pk��K���U�E*��q�����/�5?sui����um���e {!���ӾҰVV�ؾ���b1=.>w�W|��g!�����X'nT��S��#3w�%"bx����o²ojfȤ�f�O ��I�W����s*�ɞh���?�R�p�a����� �>jxҬD���~ {�x���y�����z)�o�
��|��^89�8�U�]_^��KF�'ÿ�t,��E��ZS�e$�Xȹ�&t�7��5���核e��J�[=z�w��9��Ͷ�K)=o�AnU��KpI�x� �ڗW�@h!����T��.��<y��xM�ҥRUg?�=��@cV�" fs�ωh�W�?���С d�7����H�\�����㙊�V=�#�6m�4��s+��l��Q�	�r2�2"�0��j $��mB`� �����z�	<|��p ��g����E���|z�c-�������-�E���y��_sD�H�|ߦ]=z��tֵ�<p��i�f{���?�[���@��)��(L̈́�U�,���8�6U�x�]��+U�8U'ߘ+箊%���K"W��{�2�<k�
_!)q���+ۛ=�ξ�jB�Y�`3J��Vz^�����\EZ'�/&�&C��.�oݨ�R���|�:�� x>!�7��K2R:�/Z+5 L���~��\�!�K���f��'֬�-�-�{�۩��� ��C��n�P�C��a�+&�ֈ2�`x1L�o��+8oP��|�ӿ���F�s�y4�z9����5���A�V+(j`UO��#��@� !+JP&��c�"U�>#�7FӒ#m��MK���|�k[P��^#��bV��.���!���^�
(��M�3Ol��,��ד�FM�)�N ���^�3��j�/U�>(�:ȕ��NqŲ��`�eS^����D�$4}�ɿ�[u�'"&�v�|��?s��@�uF���ʽ���0=��N1ym�zn���Ai�z���ȑe��OԴ4J���xa&�3	9��.��z4����z<���JJ tr�'6�Yd����B���Vk%�0�G�r�Ś�f�ovԐ{��k�#iMј��8l*�{�Cr����*)T�	�x��D�����5�e�_j���m�e�mW@=�����2�#�����mT[F�-c)c��13�%�O[��HEe��ۺw�nX0�;I)�b���B���j�>����BL���l�SX���k�����-���7��m�
1������F۸o�G�痀huS;c���@�����.��"<�Ƌ�vre/����6����-���L��� ;�4�L~賻�f�Mʭh��v���A;0�iÝ�ɑ��~����IW���;���gDhx��c�Q�����6��k·b<{�a<�zc�z�GM&*������j|ٙ`��12�1�-��$7}�	J"a��W�ͪ���O?X��}�%Z��������=�ͩd�~��\`Q޾{G��ㅬ1|a�(�Gj���!�Z 7f�P���VI�+���=���t����1�(�Xcyc�Fǝ#�ax�^W�z�����A���y���½�S�n�	!�&b�3����p��M�R<�S�����R�8mr�a�4zDol_�ͻ�HP�����j:�D���0�_~H4r���'��hn�*���"�0���M�
���(���f�-�_�m��غx�<�E���С�c�ߨ��[<9%qR�<�P^1�3ف�Z�oȸ!�V��шB$�"!�ǁi�������-O�4G����/
�����W���t�]�!�R@�"�Zy�̛tD�K�Ù�� +����,B>�����'��6n�IZ��ʚ����F�鮞��F,�iJ��{y� �a-L`�i=��ؘ���8�nߎ�O��R�Dr���.̶�;����G�4�_Q\�4��þ��`��_�qp�B�������$��f�1����1��K����=+'����3� �C5+��*�sf����Q��;(�(N�ޞ��i����@Fٴi�������<���˸o�����[н�pPUXҭ�� �fr�mFc"(������6k/��4���'���
����پ<v��6�n6�h��6�TT�J~��� �bzt�&������%�� `i�n0�/��;'����yS�ؿp�6�_�U�}^0+'D+�*�,�ro�~4����[��+�AN�Kn���Ү�f@�)�@�ojQl����B�F����uw��b'y9���ԟL+ys��\�h��m�hv^ޚ���]=�K�θe�ء��@�=����d���E>�s��CĆԿ�:ưm��Fn50�.�zV�p
놉.��
*dۖNh܇���l�K���(|���Q6�AWE,�`�U98Vȉ��b}���S祍�1�.=�B\5�& �44��Y�Ka4� �V龵B��v�U���]��(�� h016c�E��E�sPv�2U�[Z"Oȡx��:���p׼�ww�-���c�������,ܶ��ݛ�[,��%M���Fs�R��gv��MYyY�_�R���EL)! F~:�v��60��κQVE/Ⱥ�աcV��!����7���#`kFP�Huӿ��EZ���.Ћ��YB�DP%9��VA	+5��k��Z
5SE��Iߌk����
�3�hYZ+�LE辌U?�N?ݙ�:ֵ��E�ҳ�j�)��uXywU�n#�z�1+�(Rk���T�����Z�'�������0UP5�����H��a��0U���7���\�9ř�4l��k�����۴�,�	q�=�Wq׽��k�P_��M�ڝDWX
�G�I�ͣ=�9�p�8$����7�Ǆ�3�3�7d��;��3@rE�;��x�"dx��5w���ٸf&x͊���hũ�&����W��(�Z���;O �̖��׿)��;��-�b�
�a��Ӆh�F�AJ�����x������7Z���M���_�O�i�;1�CN�S;��E������:FZ����e��1z�M�*�j#�N�b��a�r�c4��eiV �������O�O��!V�����31��&6�Uo�'c�'���ܤ�4$�����7��$��5�x����KT�<_	d�,7��Q���$1ډ�p{p����̏(��*���i+?<��I.B��3B)=_�.c n�%���Oǅ:�j<�GG�Z�;v!��Ay�r�ğ=���\�ȧ n�	'��$���O�e��Zo��'=�n�ʬ�qҭ�r@��8�gP��:�[u���	�2w����D���U��x-e_x=�m͎���X��/�I�\yMѝ��<fe�r=�W=p�(���D���|�E�΄�wA����Y2/���/��ڙ���ل�];Gw7���zspD�2�%e�|�N����I����x��-V���F�L��qĮbs���t���f��B,>�s1*�e�F��iyՈ�s0_�l:����Vʧ��[҄?{���YNX��s|Y�$�L�ݥ*��놷` Yp�D��T��hȌ7/zkB�o�9�&�N�����*L	Z�>�^d����Ӊ����m���OAsTWv��ؙHPU4v�rq���W�1���N1��$C_��xD�u�1���#��|<�AN�8$gm�������gV�郍`2.h*�ql"0����%���M�[�n_�@�xD�a�:v0=%DI�)J �b�M���͊`����Sn�Z�008���h��m,UxԌG��k�-��vQdv�>���f�`�@��P<��c��8�h�NUo據���Ñ3(�'���ϗSe�v��C'n��آ�i�6���_��G :'�T_��{!I�*�oRM�hq�d�$jLn�I���Y�L��d�g>�$�����M8�V��x�9�Ѵ���4vuZ�.���DO������z�P�oW�.sWWP�d�U� >Hˉ9�˅9�i~�+�-�b�]S�@�@������}�O�-O�NV�~���pZO�>*8���j~(϶Ͳ~��ϵ�=�kAD�����ٹ*�K��"_��֧NZ1F��O�7� ��u�)������(�By�����T���F��hy�fm�KD|+�xd-!���i��u���EP��Hy�뭼���� z�7�0��C������R��"�W��^FyUlb��
EөXT�˟�`gҵP���CM�N)�L�v���{��~gL�گN~�lK�#O1B0�I��ɻ��	5����2�A�~p���u<Y��I23�q��P��DA��m�Y0�����xJZ���|�zgH0�_ �Sx��Aqe��i��%�?@e�8/j�]K�X�ް��V���:��PUE��ix��Ӊ����>���V�BΎo���pn-�˷�)�	tBM��:�$l��8W��祜4ʾ�UǰV�C�4Z���[-��!��'��ԃk�3S��(LpK�jC�oK~�!%����X����07LK�uN��!�t�\1U|O���ִ�/'���ՄL�vd��B���o�779���m����|䆕��>�������$R'Oԁ7D
*ALhA�-
�@b��&*x�����'���jEYj=l�&��� �*��F��W��.
]�G2L-lr��b��Łt��cB�mQ=I��D��.�03��F�B�����sYK�M���u��_nn}~)$\	o#�p�f��^����LWY���t��X���,R����0��]�Ƥ�Skw��b���=2i'��M��� ��PS��wX����$]�&#�d�n�5�t�l ���d��J��6F�rR����%7x����M��G�=~�4@���G��t�Fyd� O��u�O,��e[4G7�|�fR"T��i�bm���c����~�0��7�2��ov�>kRz��JvJ�܄�g��ck���.���f��L���A����/�^e��*� ����n*M�$qV<��i�zW��n��9�^*r9�%P����<�B�>+������;��E���옔��Oľ�}����-�˛��l��W*�5�J��vl@���_���3�]��S���n�z@R�4�:Mf��[���w>��+�����N��`_j�gk��Q��l
Ө��Z��V�;�<�2��jU�G�k4fC�k(�|����OĊjN�~z�E\�Z �	�D 39ǝsV������n��g�w�i��ۃ���w��
�$u㊀��cㄶ��zBK�c����os���Ͱ4e�=�K�"�=�R&M�U��ͥc�aۄ��'̑�$�=H1"�\�2���Ɔ�0mːUoю�����
|��r��6�z�$�8	��b��'��}�{כ����ܷ���C?�m��3r���'M�g���:D����ӢWu�s��ş˽ ����J���&X�Ls��e�6[VQ�@�P��A�I�)$�B�pMHdN]||9TX%,V�u�?qv��7q�1\p��X�|�z�d̢Xg���,[L�E�>z�)y%��LCs?�F��R�5��}�y�e�h5}ě���ԩ�_i����� 飰g�A�>udψ<�
n���c!�N�q����Ƕ�~S#��G���g���"�z���R�m�ɑ�sL�Tv^��K2�2�|lhx��U��6��Ո�O �M�V�s�-�Ŧ�' "�����^U�4��ʌ-��9>*	\�����a�!��`��W-���w�'K����1ڰg��
�����v^|�����L�,r���WdԸ�����z6��<F}��+��9��m��f���0�K�!�w�ڬv'��JX�P�dN~�&v�'o`�#����aΤ��G�9Ll���z���A�Qx?�/j�C�����A�͍%L�d�-0<�4����"�-Uޜ)��hИ���d�B�d�
����]����;qB,��Ǝ�&zb���,�1�\r��UJ]��s}p����l�_��4���r? �Ju ����?���ݮ1�ټ�B#��S��\}|-Dd�Jz����[0�F/v2�����/5li��r~utGw�Q\TA��6�"����Z-��r�`�62�a��_�ׄ�#��f�O�a.��H��4��5�4�O�C�X{������)��P&�����x�Q;�y�qZ���&i-=*`��t�t�)�9����'Rs���5:�yBPX�gیb�!N��5%=@r�8C��Nx��}�֍zB�U�~Dw�3�r��b��7Q��Z2�`���T�dN#~m[|P�W�c՜�h����\����8�����B=�A��x�4o}R�d`s�?䙑FA�^�v�@8�������nt7�[��e�����;�z������YF<���d�G��(K��:�Jqgj�]Lk�ct4^2���}�ѶVM!��6���!�}XH~�U{+*��!�^�� ��vkǂ�v�bK�2�0�����N^�"^'�u��!������C�͂UЦ#4�e5�3h<z{r%n�d����S���)��A �*#�0F[X?���yp��=9ޘ��u��BY���<!���</��&��7�wrG$���+�H�d�����zX�0beh/��C_�Hﷻ9=(>�z8�Y3�=d���K�'#/Bo�d��\�m B�܃���f�`e�g�1�u`E���0Y�z��FR�q��i܅В���� r7\B�2o*�^�īO�f�ćD�{�mh�?��̲wTD�9������s���CFo5�q*2�H{�yw�tQ�+��I�oaBrf{���Olo��=��(���A�_�r㰊�'��WS�ys���&5,��c��Ӟ.������� Ee�(��d���b�%M+:
MB��}��d�3Ⱓ=�<��a59�x�l.}���^)�+䋵��=�eY�1:�{���8Emu����&E�����SVn�k2��%
��!�� _�ѱO�j�Wo�J��_�F;ɭ��Y��4U�����Td�(>j[P2�+tb}�>��A`Mq��p�쉿��`?��
DXq)��|^����$�a*�V	T��8N��UP] y}��e�~��K�����eG���u��Qo��l]����]]9����q��d$(���Y�p���jb:�v���h��<���� �1��ƅ�j�픋yo�&������x6��EI�laSi��h~F��A\�����D����I�y�!��O��<(ǃ�Z�1EG�g`K(�R[����}�J��A�w9��c�^;��;���~�-�P{�$�(��������c�bEf\�2Sŗ��l؜襙Q���L�E�O�+#l�2�8m;�W�r�Ԓ;"������!#�;���&��솬m�H�R.ccz�٦2$\y�K(a�$�9^u�����B?�)h�o��G]L�@?��4e#�\�8����\�.m����G)pW;���8NF���W��A�i{՚��֕A]��p]*�'`���C�?��c�����!�r!0�8�r�]c=���$�<>v��4���C�@���k�m�D'�`Է�@eu��:����R]/?C���$a���n`ͯHm[�|{�Q�]tH?�)�����r��ڵ�$?z�@�Q& ,� �i�c���X�K���:NO	�+�i(��a����P ����B�g3Jܶe����u� ���)��C�o}#��?<V��}����{�Z7��S>⯮�+I������
�[���\ۋo.Od��,y�6�������?�V�\e\�r�*�g���G��	Y;�ӄJ�]U��{]�$|^�� �O]��?�0r���B�Q����/�	
�3�vq�@�'j����_JL��G�~��o�{��d��d��U���Ȩpl�p�\�`�g�C? ��6q*"�R׋/�	v8�sO���~����8)%�GE��b��ԓ�:������Lh?����f-Z�����%)��_bIJ.큔�Q�m��8��	�:�PE�c=t=F�И�hE���K���G��ƒY�Dg���;����{��c��ȴ:��5���UJCPɓh&��Y(�3���`jN'�
E�$�X��5���s�At�\�+�`��O�4��|� L��F�)Rj���g�<e�Ts]�3�.ZJͶ+��N�$<�"�'h�����5Co�X�MN}����{�w������|�a�\�so����Ǒ���x�( �튷!��A!����d�КB�%�|�]�~X�	K��,�Se�a����4ЏΓ�:d��g�v�)3)w�a���)ETZ=�5A�e��7����j��{�'�7�M�f�K�=�z?�%�/��&�V�j��VZ\V����)��#;��4ƽJY�r�t(Ǩ�n��A9
_���|�Jkh�ҽ�2N�sQ�D��-�+���d�G��e$��pt��~��`2��bB8�5�^ j�5X�p��g?�K������݉��Ӎ3֪P����VI�hrF7 �ٸ�-f���f�$�r0{n����I@���(������Mڎ��k6��@'ߪ�<CE��9f���zK���nŴ�zJ+>�N6ݺ����]��+8�-N���Ŧ�GU�f�4BC=m��-�=����H�$%��D�[���b����@�\�m�R�� j��fC����0����\�I�:n���Q�ρ僃��˕8��N�7��2G��>*�I+ʓ�[Rp�3Y�7�D���wr�(Pr�?�m�)�0�� w
a�W�1��K��tz�Je�Y;?�z�9���=$6��@O�?���*DU��̸x^,z����"�V>a_��1�TK���!:�_>&�j�.�
�9�6o�6�ڋ�0�̱j��l
ѵ�;� "C'����ɨ�(��2ce�'���¡��/������R5P0(�iU�������{[����i9�tI�����$�&,�
�3�u؂�3Iޢ݀�y�I����U��}O74��E[5� ��Y*��G0�_-�ɰ��!��C�y\��qA)�O
D�Vُ�-�B�鹙,�z ���HW�D�~"����zͬ:9Ԥ6G@�i?K�iۈ��bv�_�Y/�$X8��<pE��h����i����}�"�{�e�X�b�V�-g�+�D���ɦ�OkXS��іʔ2^l��<��M�:��ՍH�t`E�˥D�cU�>W�EW���dC9Ք��Y˥[P�M#�'����{�b5��C�dHK'd����}�(	�I��:����IӀ2վ��n���"$C�S?���Z�މy~�3�'7�RgV��fI��ۅ�E�L������-��b)G9�Ӹ�G������z��Hk��2*Da���^J5r�X�]َ����_���[hc����H"�n��7:bM^!�@�Cg倥d��Ďl�M��/��0M���U!_~
ʸ��#��U�r���0cu��>qä��ʱ�R���kN��I��Pa�x�W��烞-;���P���Q��ëJ�˳�������[��{�J�[>[�U���/%������s�QV�D({��m">��I�E��k�d�မ��Y��p/��ǿ�Pu*�Ї�%{3�.�cc^t�9(TQw����+�I�=Î�*{�Z����R~��X�=~AnŘ%$;���6�)�A�����[��Յ�� p2N�^x�N@���8�7���&6�����\h������HL����'��|�@�F^F���{9��A������𐯳(�8iu��-����� �-07�v�f5��n}?��z�����؂y��W�rUKBvW�x1zC��.Ty����&��*D�K
���#�!
+��U�
�
�8�m��B	�e�8��{�a�>�.�"�lV�����S�6D��� ��.D���v��h�3d�ȷ�AR8�y��ҙ�΁��0�1��]Rb�����"��RU��+V��؅��-}��Qe���|�Wh������N�P���¤��OH,,q{���7�ǀ����6��B�.0P�/tcg�D��_.�T6g9�d%/���!���ظ?�#Pf"A���(D?���6�6�>B��2�;��C��O3����Oc���og���4�$��L�[���[3�A{"x�-X�����u��Z\p�6�Qw�e�{|_ԺX1�8������l�%6g�����~�j�I����JO��Ӌ�Iw#(��ƨI^T�#/ք���C��3��e>\{�6�7_��2>k����-�`{]f֐���A�-2�:�9.�s&��@��-����f�f˱��ь�n����V�l��8k>n�CI������֨[J��X���ѻ�#�"o�V���4\N�T���k� ZVt��@�G͆y�Ko�^{���߈t;E���B�]g���MXܪaU��0k ���h�����x�5$Bʋ�=xW��jt�=k1?������-3�sRϛ��d�7���,�M�kE
�|*n\��Īrk'���Bo&��% �i@�L�uG�iL�~JqU��"( ��Po�,�T~\��\����4��BD��V�:(�~�zUO�͓oӚ�=��M=H�0�)����P�(�#-s8jΖ����LZ���Q!<�OH�����Xpۢ]�ݸ6N��������@���l�w���� -��[��{xa=��sN���.��m!ٍ�؈��L�y�-�y���d��8�\���=�W��&�S�IcU@1�Ɨ�:�Y��a�����@&��0MF�3{4������m[���`�@ԭ`���4.~6}���g����~*�"�c���*�ք2K4���C'~:�o �ڏ��sY@��c���zC�7 	),��L�jƻ�4�y_�>K��@P��Q��hװ�|7]�I�5;㰓��P%9����˦�q�Zr*����PV�W�axX��@�1� ��L����,�����p����]]m��w ����Ē�#��Z2V32զh���H�R�q)����F�ȏ�a���
���Kn���+O�y�L1��_{�0��Dj�t�"��;Z�E�'r⸵->0.9G����`,�S�B.,EE�M�~l��'�_m��i�v�Q2�BW�nI���J �N�� �-���NS�p��l�Pfa�W�g��_@h�����G���!��3���_#�m�h�f��$�M�V�jF����Ǩ�Ev�^��jT$2O�m�n}��Z.�"���h�>	Ng��r�@� Awf�S�|R��̈|z���w{R,po5>���|]iay.5�`ө���wk�z��U��=���b���|� ���vZEE�D�l�ǵl66��b�@�$FU��L�:�N�>A����L�r���ͩ�
@4���'�K� �YŌZ��\Ӹ������U�"T"&��3�6k#�F-q��u��"���/y���A�ؑ�y:�:�uƫ��OR'���Xm�hG�ziA��#�#����٥�,��׾�%RHZ�ci{2�R���� !Ad������l�����6�%Ǳ�<��n������{�l���+X0v���m0�\6~~�V�_�j7����wb$�r��@(G����l���wg^/>��t졽y�.��m%��~{��d;��_��.����z+Z\�p$�1Y��)�d�d82�fY��$�u臓�
XL����p%^���4#7GQ�����B�O�)Z�$������*$�P����8ϑr�u �"	phV�]�'T�M���&�CG/���Yˁ���� ��A����R�k����mYp�ަ��d��8�,W�y$~�������X�(�;@�������Z.�Ǎ��v<<�m�C�ǅ7gǗ,2Fz�r������ܤ�{0\7�7���T�L'x'Z�ׇ�i�b���	�m��D��%E�{���x'Y�e�_���G���v<י��r�T�?y��\ݢj�S�o�v�|Z/>M�B��sß�ُ�k�q��괞a��~�V�#a�o<8���W.�W��M"�@�aN W�
�.� l��&�6�W�n�F�vCצ��\�L�}���[J��G����QI���]B�n&@�UANv=BT�rHK=����,(�����N�l�h���3���9[d����h�f��lD��en�+�ۣK�wwaa���"�C��j�A!�fD\�8S�4a�O�%�n�jGF�G㉚���e܁@|�374��FD��1Jd�?�@����ـ�%�^£��ˌR�|��Ra��o����/n�8��۩�R%�4S���:�֔�I|X��tg��ߖ�N�dfH�8Z,ƺ�>tU�L+ =�B�ڢ��x�`��qM?�D{0*�A� E�к�8�a5%���Z���E��M+Y�_�^y�㒣�ǯ�'Z\5B�̛ w��5�+̎�2�:q�7���)�^Q��s�2c.���z����A��ݙ]��	d�i6����'Y�ڏ��3����a�&x�ux�ծj����4�/.�%��ڜ�"�p��z��)u��gb;�D(��U�-yG��m %s�g���U H����u�������T�.��@ydu��+�)0�q q�q�k�X�qw֬�Z����D|� �	�6\��كg��YbH]�E�w�����Sq3��m69�u��Y���p:\;U�i��d�r��{��:]���"��!O&�5-Tn�^�i��>�4�w�� q���E�Le�%���p�0�^�N��*s�Bv�o.,_�o@��B�G �" ihI+�"=0f���p���ϝa#��4)&��P�4�5q��( ��<�5~M���ᣑ�Z�U�h��FD,),���� ��(#x\u�����5� ���o��'f� n���&k0�pTJ팳/
]g֯s*lI�+x-B�)�"����N3vZ��W��h�2��p�S�2j��S���z�/94� u�,J��G\�^}f����5}���p_`<�A"�������Qw��J�2��Q&�������T��z�ǘk�v7��@ܚ�׈_"Q�1~ٻ���ǁxkӤi�S�X����+�����4*3I�L�����S��>)j� ���|�%CO9�qz�4�/�AꝨB6*�2ٞ���}�:V�N�1�Y^o.' �^�Sm���`MG�e~�n���w$�c�p�&R���?�)������P���������z��g�$�j���i�J�}m��D,��0Q�
S���1���9u,|?ԛ�Γo�e%{�:�H�ŀl�����B�|&�{�&������S��/$���\�yUI��~���1E>;�6�@I 8Tm�Ջ���?��:'������(���q�K5�%;_	y�:��ӯ��5��pY�A�4�ơ���J�K�QK���!7�Ǉ��wL㠛�l	�Ռ�e#Iӳd�P��oW;P��u�B�7C\�|�G�t�4B�G�m�qTݹ$������'�)]9u�!�*7�@��^3�S�>��@��1U�gj;�o��,5�r��ʞ$��>R��oӊ6d���n`�+���;���W��}U�#؝�!�o�Q��Yq��,�d�j\"��P��U.��-Lˊ���,XU'��^�}U�d�M��p�`��,P����7/��6��C�:�ۗ�l/r�TgyB����K��r�| 5=����RG,x��F�%�S��~�a���5��0�Y�ɥa����\3&C�ɚ_�n��byM�Gأ��3_��C���nӯ'�Z�X�6��پ,�J)0��Np���qKv�L[̒C��q��n��K�I]|�V������,m�N���M��������B�"_n���LV_1��0]�Kҝ�O%B9����hH�j�5�݈��Ŝ(�Is�{{�j;�j-!l��A�;y�b�s.��a�sRä��x���Ϡ�b'~ey��F�����Iϑ?�ҟ��H{��.��SQ<����{�
]>�L;M�L��P���t���Z�o {���)�Ț~�Yn1'�=`䂾%�qd(�������2��-]:O�L���gNK�������M��sd���������+V�v��
����WA�n�Co���A.�#O,�$�HU��?s^��@up�����Zf�G���`:W�(���� ���)��U:��"aA�k�%!%�e3�~�Րzm�j�����_���E� ���r]��̜�g�u�i�k�Iw��9��ه"�R u�����W�H�B����u��v48K�uu$2it�=�~)���\@rSU�� �J�/���-�+d��=��$JN�߿��N�4��@a&�c/j��ȯ��?���υ�,w-���F��A{�\Q��'P�]�PĶ���|��3���od��C< JA���ㅢw���S�Ƙ.��D�+k���_�D.�$�e�W!�g�8y��K���5_~�RHq0Bρ%���l�4�F�U�V�&�K��QWf���W�z��G��{��`>Z�q�ϸjY��dÁ<��)֍���� Q��Ǒ_�m+et�&�������b:�ȝpuy�V�g�h�&Ǧ�'��K�@,(xڍ]s��g�p;�S:����I�$������5#�&-"4�:;��e��6̆b����0�py<Ld����i�`���EF�ֻ$ű ��7���v�j$�?S��4�O� �笹N�.)x��{4:�����3}��� ��6���
��É�Nq�a�q .W-�Čct+i���Z�#���-��	��l�Q���3�����%�I+,5�,}��)��G�� O���L[�h0�+�EX{Hh�@�T�R��n:L�,7�,�Y�JP}���@�K���?g���j��%�F� 
�4B��+v�BF��0�%��)��`,���B��s�d�J,/O �cMb}!��_��(�4�<4BVb�ff��uYB�1I�8�ӥh�jw�Aӄ�m���迗Z \'���j;���:�W��3ϔ�$c�8i^[H~f����л{am��"4w�h�p�S�x}�~m��=M�(� �*L%�P���/���+E+��a�^�ڶ���������v&e7[o�����|C�J�
L���피%E8a3��0�%7?S�2�,�Z��B%��*�rm)=J���"s���U�y��^�H0��Ԃn��|�o"�� ��(�P?ؑ�h��Ah�t��aҕ4nA��ǧ��Ķ��9���6�t��:gu�vYub�u�`Z�;ЙF�����?�S��O{�-�!9ޛ��4)�UN~ B����9�k��Б�/~F�?��3DM�}F���En�km��/�&_{l"Wڽ dX��"?�`�9����*��Z��J`	�Ru�R���X���jTOg6(-��K�,���V+�Qn�텯X$O�4�p)=�2^�����t�-�a~d��!k��ペuGtc�3/H����	n�S��}a���Ae2�5��c�4��Y����T�L�d���@��#�$�//����`��W���r�V�~��FW6�W�o���!��OĊW;�3���?
v;hLM�t�swLLi����FE��l8�V��F,���G�4�:%d��(���ƴH�1�،���[�U����,��p�`��SC)�_�6����ѿ(�T/��1�@'*�p �uϗ�"
;���y���C��k#%k8��=X*�ЍH�(4jn��բh�:Q�V��Ϟ����'-�J�\gL�����:�$Ղ�S�$l>�6�tv� vk�C��U�@0�
%�#�=WQʔ�2��I��RR��ڳ�NXs�9�tZh����æ��٠׊�T��$;v\΁���d�:O;sQ��h�E-�B"4�C�Gd��S�!�Nhc��d�iƦ�V���+|�
�����Hβ�h�	U�c;크��Y�t+��g�1I﯍<��]�pL�g���pe2򗅖�_��!�"�SY�R���LWN��:�`MsT*�⟧٣�u��HX�f���CwL+�8i����#U����Tf߷ۅ�s3����h@ v���M�<��O�1ȸ;���*/��,y���a!�����C�h�ߤË���K%�)�Tź,/ac����'����̷yQ�Pb���F Z�-�1�a��X�e_#��fMx�0Q�d����M�� g���΋qG}�}p�O>��$���mR��D~D�+	��{��~8���8��s.o��;�J�]~����mX�������w��r���Q*O@�#�OjҎ�~��vA4�_o��f����Y$���sd��t�������V�շo�2��N�`5"�!:�uY�8�M(~��b�uRy��[2'f"zp�@�o��V	��T�դ�:�C�3�,����,ۢ��IQi�	�H��Z�*ĵ�-� x���H�9��+�8Z����j,c�d�]'�C ���h=ݽ��3��wGnú�`S�P����;'eM�I���� g(1����K1:��YP/~��8�OD��$���0������ ���M�ok��v�9j\����)��0M@�%��p��E{_���ӨF=(mv�*`��i��Q��u��.���y�6��a����U+Fb��9\�FW�ܬ�?���'>2x�f��e�M����R]��&��}k�]&��
[������v�c͆�*j��X����"��g{Eη?0�C��s�yy0*��(�Sܗ8�ͭ{��B�5�Z%�p�${ƀ4�㢎�DP�3?X�b����ʔ	&ۤ	�%�zя��!F�a[�]���T;s��i��P��&e��i*���/�<�=��nʀm�[	ۿ��)r��;3fQ��	�#�Y�a��6�)NR��)6x6?��
�!����E�a�3*Y!�o�
�����������ؖ{^����=>���!��l\�&ݭ��8dR�Lz}x�eR�������)颿�Of���J��y��1�`����kb�4�}P,:h��.̼�'�I��xT=+H�����ah�`���B�$Q�?�6wKAj͖�!|A�z��I�W|]�3g�L�[!A��3�jx�lfh��MJm-S��ǅ_xV�N��7��x�~��(��=5�k�Ӯ�A��i���qQ����h��o��+�)r����)�F"��KLLj����4'���4
���̶˓X�k���DA�?䭸�(MH�J���\�2p��;��b�DS��v�w*4��m���.C`�S�����j������cA����9Y����瀱��X�؆S�5�>���D��K���mIy|�Z�OJ�"=�YV���:l��_L-�Uj��m
pt"���֥QU_�˹u�n-�D0�!�P���8]��^�ߵ��
�o]�BE��Qh+w� z�N˓��R��8�GDG�:ˎ)�P�8����Ln��ow��\_�v)a��;E��#���]�"95��l��8P�� d(=��%k�(ߋ�?!��(벷0w��e�h�uJ\!�x�~2�3���}�OG2�xa�!u��L�nUX%s���U7z����?+�O8qb*N��_Х�@�l�$��Bҫr:�ߌ��q��av���$��z)�BO>E���g�sX��D����5�1n�x�r�m���]'|EV���E[�	�z7�l���&��S�F�A8���EG��?��{(�r���R���|�U��P`�V?�?[��ƻ�6C�ћզ=��eZv6'�+�R_X�"�L`EO-���=�`�%�=\�X�t�nU2�[{�jMl��a )º`.�/�����+��NZ3ִQ-gZ�*J�j Z���PZޓ�+�u�I[��:��1y�*D�D����'��E1�Ur�/�DQX�⪏��H5��(Z�?��V�0���c����5��oz���U6�:{���n�4~�	O�t��h�\�wn���G���2��K�����U9�����&�ySd�0c��j0��{��7�«Ї�a:��s J<���(��^�dN$�`"�t�DY'풟|��w�h�_yF�����pVx|��7�0�젙����1�B<,}�~U^;`� ruF��g����W۽B���;�Wf���tUd�`d-}�܁���ἳ�k�=�q�(4遪%
��a����4��Ѻ���;�c$���+�h]�ؾ��*�J�I��V&p��)IeUMb��2�\�4�:`[�)���`Q��l,��NHk��6Ϣ#�3��b���6j�쿐v=a[���v�2j�����$�99�|*��h��0Qe��ފ��1I�5�	ea0^��.��%l%�?�P�u�[J�	Ͻc9f
Y���6�N���:��!F�F���\I�P�糺���=I ��gFQ�S��i�-'c��S�]D��`v+���i���_yqS�E�?v[H���Q+m�R��`�;=l=��(t�������iJL�F܆�m�������'���[Ą��f7" �4�@�o;oHH�]��Iܤ�3��h��D�}��R�GK��ƺ���\Xh�'>��YT[>�I:85� �h�m��j��%��c8l��b�h=�m�����=�\���Q%{�Xؙ"E��l'�J�Ty*+��� X
�'7 WK�����-j	)RDe=�7Q�tCV+�AP���.2�����xr�*9{M����1��N����V̧�p
�������5�*N�0�6�+S��]���Ro]GY��v���wIJc��{ '�f� ������!;<��n�O�x-�G׬������Z�A�9���Y�	��x�%����3@OΔ<����i�5�E0�orY0�i�&R�P-O�_l9�-e.��M�ZK��UnA�a�B����{&,�4�vӁ���{|w	P�[pѵ�����,O,2ݺ�a~��k̔Ɗ78aWe;F��/���x\���G	0R��f�ɛe����}� �:xS'�5�	UH���CJ5OPJ6��l�!i'�<eEk�u=os���xBV��	˰a`C-jZ1P�A���FH���Yn�S�qB�_.����
W����#��r�M>=�8��n���� �Пxڪg}�������m~�����Q�Ǹ3dxK5-
�7\�,��������!eX��7����J�ghe`M�݃�h T�f�ͧ;��u:�or�uq��,���V�\�ݜ����I�GW�'�M�/-���ݜ�t�x��r���g�����20��ơ���lïuQ�mU*U����̠xJ�T~�M�ˈ`�g^��[�k�������ZJ\�\�����́��0��ŷze��g���
��N1OO�mb��q�r�&�ps�t�6��c
���3�L�/$0�8&M��d7�i���d������:�(��AL��ӂ(�l��U�\�&�ت�Qg��_�H��9g�������"~��^B�g�:w���C��H�z�q�_��Ą�K����C/����,�l%��P >
Wو�!&'˛q�!��A��,�er�����*�9���T�]�b�+����y���>y�CAk!%b{���\��R^[�_	�]��&�|�͙�Ӵr��W�I��x��-�n��.ȨDN��~�R�S�
$3�^���=��<��듵���6�3[���|~���V��ZV���A���d���[z��A@̹���(^o������S�τM�5 ���=�EF(>��_S��چCP͠�q�k@"�1�X�G ����xc�@�sW�� ���+��aM�X��;����4͞�J�אּ�<if�0�R _?�c����:�c�w�6��pv�+��ހx?�]Z���X���3���ez�Q��+�# �]U�f��;)o!��c��P� �؀�� ��p�(�b�A�����T�H�	{<Iĕv#
��f<P�FS���P|!���T�᝹P`���)}�ld�r=<-K���y�v�d���FƵ��)&��w�#(�u�\��Ki�<c9�0�)�+��aM�g]�``��<o��[�Ea!mȞ#e�$+s�MN��}x� aj��d�k=a=:L�8�V,���P��[oT����*vT����j+�� ��\�'��˽�Bl�H�F���:�.���6��0K� R_#���Za:6����މn�Ԕ��g-������tA�����������	�|h>�����mJݭP���QSG�d�� ǋ��ƵU��x����[�x�� �κ��>�kCd�+1���ޙ���8��T�D&���}G'�ɇ���������F�mG��%b�tX��ʅ�%R�1�TL@T����|�ߊ>��%�
��E����t���m��і���F�J�O/�)��.�+qu�#j�[ �^��s%�{-;��q��,��!RJ[�EjTp5ɦhi -�I U�x��;� �E�M��L��M�j0��ICjɅ���^� �Z��Ϛ��Ӽ�n�����v
�%�౶[�i�(+έ�6��f@�{���N4i����[�`:y��`<�b!|ڎ��6���X���#�ՠ�1^V�L\<T�hVu������H���c�o��U������b�'t���G��{�m߈����K��_6��-{i�2/����ՙ)oeqI�v݇�"�[�Lx@�6Ɯ��fZn6��g҇��<+l;{F,��<�����a��D��=��i{�20��9�u�N���#����d��y�pX���㌒L��lh]�i�O꽝�k������
�l����8r�A*�f^�v�0��'�mA���)vh9C��Hq�ʷ�d�oq#�w��m��EĀQZ�Ễ߁Ƽ�	�lkNil��HB&.�"�,ę�G20�
,���M�$�T��6��Z+Y�.P���gQ��h-^ٱ�/o*�BR�d�=���(�*�ye�T��PE0h� @8�m��$��x�w�m3�Þ>#Q&���9܍�\257t�(�!<%?W�%��&$�
��'���#��2�;�HpE���*S�y�`�|ׯ�/�X>j�� �������=Dty)��v�U�B m�u�AAU_o��p�}�]4T����u	?��:����:/��A����Ӄ¡Б�=ӟ�4����ft"����,]���y�/r�vaS������?W���P��xb<�g)���Nn��<��m��V��y�����JLnG~��(n�D��j�*&m���?�ݛ꾀�M��y�% fᴂ��j��J�h�=[2|収�>�O���q�L%�Rak?����0taU�^8q����I�O�����d�,�'���N�I���_�A��M��ع؆�N�a��&���R��_>�{�e�G{z��Bm�X��T�jk�^�����.�9kB�w�FG�>���/�d�[�%�f�C�Z5U0�b��_[vZ��e�)YN`�B��[N��4'�ݨ�w�P|F9��a�1G{�'[F�U�gĚ�YsLoq�(P�a8M�� �ą��pBujrA�vD�A��j!�)����o�Yc.��R�=@b��o�E��yN7:3�$�i�4DM�9y�an*�(�u	y����sK_d�Z)Z'��@GЫb�H�2�M�����ܑ��w-v�I�s)f(�C�`����89��1�a6WN8<U�r	���X�!�2�M�]�����+�E:���(Z��M�%R�T����LÌ���N�
k��̍�bK�_�hZ��l�T�?�q��6r�o6
z��^4W��h�~gg�n8p+`�߼�_]y_���l|M���6���{����.E?�<3�meHBy��R���	JB����E����ܾmD��ψD�D���s�bt�sA���B7�'�si?�R�2
�dYb���Gp�wuF�Z:˨ل�s4����(WQ��J��?�A�W$�{�k�0�7���E G�ܵ��l���eS1���{�	uD�y�=���{!�?���8tiu�]w������17*K|l`
�m��CX���l�ʞ���4Vw�%�\$�%.y�sҕ��O�E�����nw�u����	F
�<%yCB��2���Bq)���������#�c���nQh0{�ċ�ẒE~��h�!�<����V�y�vc^�P�`�*��l۱r*Vn&�\��8/���Nۘ�[:����M8��؉
o� i���-������s�i���-x���T����GL�XQwWJUL��Z�~��9$D$%��!��N�p�)ZI7B4r�2�������\l~>��R˜�����쉗ү��D�.�^�� ����u&]Ne�$Cu��~?*�ٻif;�d&� �&�$JaX�0a��|���X	?	���f������h�~�XBM�ݸSMm�c)X��z��������8�(�w �/��0(��-� ǿK�e�٪LC�
d���s�38�-;||��+D۬h�����'� i9`���r���Q4���bۜI�cU�;�����ԗP}���y�b���	�qA�80U#�fY
@���:�>�oՒ�9�h��[�͍"lK@n�:�{{�7L俵[���x?��x�����)��ɩ�=�b	aI�Is��̗ 	b|7��;57K;B�.��hg�DJ�Q�;��z�`�`�#�{�jB{�KX����^��2yx�@�N2�F�U��9�<�|�ZP����%��^�$�
��ݢ3F��*�B6V؅��D��Hu�b���V`�Ǜ�m�e�>���bq�4;���vV=SX�<�}kԞ�~�&������f.x1�'���s!�'�#%�B����wg��LDmkimG�jA6����*����V�1�)v�Je�?�	%؉?�����%��m���է��cxen�2J�B���3�/����D���Ei3���PgY��I�����a"W�~iU��^Ǔe�����8/c�	���3$!�	&?L�[O̷�֦��gp�?���V鿬�4�A�F�`ݼ�<��ߠ�4�=e��i����B��Ed��>�Kpꆅ·�|\c������\������$@�m�Vob�\�j��U��ũ^�v�A4�g�WD�w�����������~�T'��ȹf%p�B�B��&��:G
~ECP����`��sa8�D�D�z1� qO�#�ٮ%��"�Υw���-E��t�}$<6'ĥ�(i�9{���� ����o�_/�F��x1`jO�R�����l0'#+��t�rN2l�m0e�kgP����e_�G �e7����<����S)�(��\�r���b\�~uQ����sA8~�8ɬ���8
u[��$.�}�4�,�찦��8�o:I����e�j�?ə���e�����|8{�@���7�<V�n.���p���\{����#]�|~��ם�9Dc���ω��������'�a� �R�{@)���DH��i(���mr�@��	�#�w�\&�k�oB�P[# c_ND
Z4w^������b�k��:�kCB?[w���BrE�@��~,�p��V�S'?l�wNC�Mjf������,�
,�N�X�p
|���g�49���s�����RKBkr��H�v�_OЩ)1;㓵�IS���.��AO��r#+PQ�n>����tkUҲ���ͨ�G��(\[����M  �D�sq�|�f���������p��z:z�r-���� w�.���8��.U� ���u�n��y�~v��t���l9ۘg7�K�"�� �M9Xu;�9�ʽ���I��{�2�EYl����l٫��m�`vy#/�H�bj�?l�C���}jU�<{h�Bt��I��:@�E��3���|�n���K�� dj���X���OA���\���C�����S��`�p̸<�q�4v��00~/�9��f��yخ��	5c��15��G2�>o���Z�p�>@̘�|;�\��gt5j)��M�i*��kw�$δ���ч�I�����,��:�R	��3����?�A���Cd:|�[g�m7#���5��c>�P�[�\^��ƪY�����{X���У+m)��Fa����c�`�i��lRSe�U-��RM��P���@�!�C(�X8�3��F��pL�M�U�-"�{9>��j,�k�>����}o�~�l�����V�o1�o�:}����UZ=l��u�(�;�`մ{H�A^��|��Q(-�;e9c���m��V�#����ݠ�.��,:��LD�3�OXL	NF�>P�^�m蓵�I�ex�f�~m(�']�����Uq�I��s_������Is�;Sl{#n�r�D ;��{{���+]��˵�V����jC��O�>^Z��a�}1�n��ۯ�IW�h��}T����<y�X���+,�5h��s�4"��h�[�5:4�j�Q.�z�Zj-�Lz�?��{����z����Cn� �I���%K���bJ��� 0���4���n�33�z���_mé^�L#��4��"�o�	�,�=�i�k(C	\Sf�B,c7(	D�%?l	h��'�eК�͛�D��/�Yh�N����Oyӻ�>x��[ߙ�f0�b4J�hm$B�]I�L�c��6D��ٳ�e�b�ECux��]R]���z��B.���˅^8m�P�ܦ��1�����z����"�j��S�.��M� �mJ�"zX�0F���գfU!�%e���ި�yW�ȴ��	[�d��)h��"�����K �����̈́����GN�������d����pr���4|�C��x��܎�4)��w8⦱�ȄB��3i�:�:w
O���}_Ч��d��{�}��b����;�� (I�y��s��fg;ֶ�Q��\�W����T���GX��6���T䮾����3;�*�q@|���H�L8z"]�%�]��l&4�F��r���rаY��l��|޸��d���q�!f��[��0�hK�(o��t�}��T#\�����X���m�����W$J���Ѳ1v'�]~���4e|w��_+���G���V����{�������R�#�?@}��n���2_�Gx�'e7�kBz�O��%��&�����ې�z�S����Ȳ|9��1��ik�4S��< ��ڐ,.ѷn%�}x��Б,B@����/!�y�k�2b��P�V�{6���vZ'����G�8�߮���F�7�J�̹������b~��I�)��9R�Gx��d�H\�����?��UΜ������8�<���Ww���{��tY2No�؊��,�q�R�j0����.�(����͐ٝLk�ɶ������*����\�wN�~�0cJ���~�	{0��6�\`vDX�%bN��8xN&�k�y��ٷ��ȅ�FWZ��_Y��z#��n=�5�N#vLD����lR�����W:�v!mܰ�DBS��.Ć���>7qһm�7 ceu���B$����ec/<e`�
0v��u��I��� )Ӥs��6�0S*���-��rmVI�ӉgǸ��>Nw�~`TqT�����&l�',��`��"bWr�Łn�p��qC��õfSP��k�1LE>���4��Dߞ��"���S1j��ڼ˾��T�&��W"���X�X�~��T:��DY�1���H9>�$B�Y���rZ�x-v�����53=�Ͼ�|N�8��檨콠㉌�f�E@�: Z�5��4�R����ކ|1NH�:��=�$\@��`�{��*_N5�Og��wFɠ��V���n��O}����.>G���8N�tVϷ�\{�C��ؙ%�P�����5u������-��wWR�-�r���#j,��I��^����n�H('�V���;q�/�	aU��e�1P��@�o�J#2y�
�� �ǕV,?���癪v�)��g��Ɖ���.L��
�ʏ+��@��M�T_­@rA�<'iN����;��ݼ  K��W��V�v�v���T����7��^ب6g>�j����l��57O���	�q��e�kYOK����m��6މ���a�Y_'9��ᐒ;����^�����e,��P2b'O�&����Bϑ����Be�'{������P�{p���#����qh�b�g��!U��R}<ސ�-����H��Cad^mB����ޮ.��P��ũvc�ԇ�)������+�e!j�Wk��xu��d�ld��MmD�C]�hʷ)U���r'@�[����'�1��G�t�,H�5F�gh֯�i�A����"5�<�T"��{����{�7�Lb�r%�I�w�ʇ��X��笀l�֧Mb.�����6��Xl�}*)W$Z�1�a��6/C��(���Q�,�̏-���O+D���+$�@\H�P�W{e�=�?�q����;ͫ�mB[#	]���$�+�M���h�x�R]C)Y�&	�b��yaI7^�,��<`�
�)�Q J|A�|���f��s��T�0��-I7��L-�P..�Z �*v�/�Wl�����N���Ψ��H�?���#UH�����{f��4�hg��R"r�DǊ�"콸0m/a�~]0���_����dуdqN�#�=��h�]\Җ;�Vhl���R������U�-�b�l�l[���D�xB��ӛ��~2%����@{�7�����l$19�����j�����R�3���%|���s�����n;�'�l�iߟ�/��|%Q�9ܶ�8��k��O�Y�Z�����P�鵦�&T���/���R�y��!&je95D���{��f�}��۳*�B6q?L����d�%���
��>I��S<L�0�����m�3���a`��b�3����'�F��& |=�%k�Z64��TiX��]�/[���ɲb�;	����l�>]�������/:t/��DHOql1O�Y7��C.@��h�J��E�@� ��gNdk�C[����e�^/�h�X�&��\�V���<�������m�خ�/6��Cs<?���M{�����Z��1 $)���!	����׹����U�K��9��g��ql@�|_���0�Nj��Q.���GM��O�r���v%���u�mq��@Ky\',�6��fdi7��SɎ����d�5�P讚s3���u�Sǩ�����5��mwOd/�:�(���0���P��]���DT�4�j��ݾ.m�g��	o��_�7�ȩ��&z��2/{^����~��r������$���8/wQ��@30nv|��/����*V^b$�)�4DĀr^kG#���	7�-Fi~�"v��|c曟V�q��6��AY�J�;3zm/ƈjmҸ-��9ʉ��0ULw_t���W?��Hp�Vdl���)-r�߇�,i��ұ��:��?�^���h�k%]��#q.�T������A�����UAk���_��Jv��~z��&A:z�og�r��6�_eB��#�}VG"7������{Z�%�İ\U��\ΣR��eD�];{ߛE�(��l9Z73�@?s-B�����b���P����c7����t�ϲIF竝���QG���p��Ek�"�4�`:����t'Z{�? �+)_����B�a�ԔlVd�]#���r�>8e�UѾ�c�z[S�I���i:�ܔΤF��'<��=�z̦�tJ�d���bG{��g|�����e�D�dU�O4��J��f6��9�'Su����hX��5:_��	�g9O+K�P�4���A�^�y�y/��E�{z4�%�����z�R4F�FR~G�W��9�����ʅ�מ�0"��WD>2���	��l��
>Ł����c$72o|��.��
�ǆ�'v'$�i�|Z��~�����1�ZV6"�-�S]!��.,V�A�N��_"Q�N�z0�f<�Pb%)�K�� 7b�v�c�;2�^����g�zI��ݞt-!���e���s����2����������f�.�c�:S
��vbv|�z�%k�B%}�:�+�_9�K�~��\����Lt�~�^ٯCr�$�S��ь�(\��Wڄ�?eC��d���X��.�6���X���%'�#�ޫ=��qt5S)�=;��T�r
|�j���c��Tu�(�O_'�TG�J�.?ؓ2��KGn�`��1-[���A4F�LN����p(��$�g{��1��j>jx�8�8�����"����&��� 樴z�a9�W��3��B�U�5k�KM����I�Ux���$���mY�,��#p�����`|�@خF ������`g�f��d͏��U�N��B�>��F�����f���e�CG�_�&��β�s�f�C�X�A�7p$��,�E�ٻ����d�ˆ�.�4HZ��B�S[Aup�c��x��=�&�o��kF	���-^]�]���+'��~�Ҥ�r_�­Cm/YT|���a��h�ª����T٠(��;iV�Y�M�#[���^YKZ�^�\�
q�F�#���ԕˎ|~�\��gkYS�A�ٚW(Y���b�l�ȣ_	�@��n���qג�h[X�7k��b
��l�!�l�m���c�7,�n9+�M�xG��~����p��d	? ���\�9\"���}>�4{��I�N��;�(97�}j���}��\���1��b����~��ZG�A���y�6��W����2��۱n�I˶qb�	F�$��h�G�la�d؀��L�8�'K��`�<��SX~+a�{���u�$s�JNN^Uqr&�N������5�6��JP�����&O���f��-G`�vvog���X�L��,�zH��ǈ9�H��~Tɡ%��0�[�F���]0��&u����;��E�5�>�� ��I��<��1���o�W���N��Z�8��h(��?5ϧ�a���ƒ�'�V<2�9E�Yn� kЮ�UGPjw"�}���ԋ�+��!ߡ������K9�W{�5s:�t*�SY���է0�>���C
���'��z�9�����8/j0bh�`ptB	[�2�8�s����ʵ�5��Y�j�YMSp�y���8�����Mo+t�V�����,�%���	�^�%�m��{!҉"'��e/��(4�;2����ܻ�?9\�&X�RW]�8������?����zcY�w���gϟ=�����Rmڪ��^K=�ؐ�*�� �u/��Ffٽ�g����^�ZDB�=���,D���j����G��fe5��x�4%�.��a%*��-�B͟B��b�n�j��N�5:Crg�u��~�ȲT�
��},,�5������s�I%����8�X�>�ŕ�
 �S�#�Q����9:���-��N��/�B:�|P^�6����~%p9�<�RE*�p���&�L(
N�{ENh�|��FE��	�$�L�}��������+�>b��0��:X�-�)���6��鈹7h�2�4;H���(\�,��]4)���ș	Y%NQ�DO'��?*��69EG�N�����G�^xz!�������"��W���Y�5�4SIl��jۥ#ه(k[�����/Z�2����FiD��'��z���s��	�F��l+�jY^���V@�O@�C�P8)C1A�\/2C��o���4�+��f�������2�z���b3O���|�2�k�*� �>V��B�Dj�Mk䓚���E��\^����!GD�z���"RM}P2�³g�q&Ғ<X1%��wo�}�E�u0��S�[0%���m@���tW��d�f-�/�D�Px4�~��w�n5�4�$8������������\������ϊ)Ew̙��ڝG����N5���~G\�x s�7]P��}zJ��\�e�X�n��=0�xX1%��+�ո?>^�{\g.[.��3Eè|X��m"�}��}J<��|�N��T����S�>�H�
ꖵA3�����Μ-vx��`B��	�X-k�W	�jGh3�J��K���l��L�`cx��-p
��o�}^۷.�6r�^�\�u���wh��`���5K]�&��'�jpp�ۼك�3�xEk5��"g�����t}-���H�_Ju��M�{&�iO�a��N�]�w�7�Y�/��)��c
2*9��L�9�B-��G��c������1:E�����Q�-O
k���:�*�\�NT�͗�� R|��8��l���d�n4$��$װ^y�K���5�d�ε��tbր���:�J�{�;E�C�cVh���};��F��!rhc:؅�Q��+��r�A�q�fW�,.�����@.�
��=�y�լw�[F�;�eӃ�#�C���No[Uє1R^���6�Po�����ʎ��G|x+"���5�Ҧ�P�T�b{$�F6��<%�d���F*��G�����}�f0��JT�������O���w�I8��/'���<��Ԡ��>\v�7-��1�8����]Mt����-��Z��x[5�ѡ�W��/\\�9,��I���!Zh�rXfG����ѥ�N���~43ر������j@�]����2����X9�+uZ�(J~��j�F��jT0�9K��%���o����ج8���=c��N��w02�~���QL��D��0�gw����F8f'j3�[�ܙ���J*l���{�`���/i<�Rh�>�eډE����1�5'}���[�����N��%W�-�O�e:�����֦�Qd�f����Jd.Rm?�ѻ5�:��bZ�]�@y�t����zHP�И�O*G*�a�ޝ���� syĩ��E�/����w����b��78�����@�\��gc1�-.���ȬϯNU��I�ӮB%=��A|0�&��+i�'���z��䖥�c$+/8G�0��������_��;�M�ʗ�3%n�-GQ]	:���@V��~'\q�!�>�t��u���{�TG�i[�J�6�k?�"hg!��o����GQs[+�2���v�OVl�p����In�^c��I��Ebw%-<�>���E�=3��2x~���Ug��˺�Ӂ�19�PhS��(R|��[�$Y��@f�a��3b��h��$p�o�Nj=�kRh:_%�K)Ѣ�`�N� �*�~E�G��U�+`������g��ң�5z��������CHZ+p@����i�v|���%>��
p��Rc�])�R�_誛�d�J�<�'�=�zn�]!n��68aG�6��o� e�mWQ�W%�F
rs����Gʩ�M$�4^@=*�����OVW.�(
����Qc�'�F�Jx�q������}�����Bi����o�_�_aV���v�'F��1�!Oƺ�d��̺(0���H���*8'd�,����Kf�,6qcP��z�J9\�#�ӡk�`�٠�ĵ}P��X�|;]��y���|�_ߏFȊG߫����B`Y��b^, b-T��\�[#�H+��W�O$���#��4���K%�������s�Ag�~�5�PHq�Sb����2��L^��'��zt�4d�b]rz���	���`�Q��L���oc�����[�6F��CkiS�j8�oɽ���'�� ���.�ߍx�޻�;sN\�cw�)��������d�v�W1�9G�l���E�R�p�S-bBB�L)rv%`Qt�cY���y�/���w;�p�<	(�%)�m(h�'�A7�卥��u��#w͍�38�Ap�1�$�-���TUr.��>�������4�LA"�L��)˵�{]X*ֺ��I5�T�*���u �YY��Xeg1�̢>FI?�R.�~���c8�B��m�Q�G(aJ�|h�I�&<c��{!A*�L�ՉSN�f.|���U�9��F�J��	W)"C��Z><Uf�lV :%��r=M���}�2z}�(hw��Ď}E> `#��=���v'�Ӯ&���w�ŵ_�#��3L�3`-�ɽ6�a��-��O�3�<�	���7���IHR�:>��+�Nr�B!��2T��`iy���4SMI�!s�>�;��#�X�E��׮bi^wN�4雅��N���B;m�K��r{`!z$���ÿQ�\L�G��	�����ذrܴ��ĵ�c�4�H5���Ӄ�XSG:Z�
+B�,��/g��HIk��*A�Z�Y_�G���@n��PSIA���R�#�e'V��+`��e��dD��_�՚�/�1�%_8ũoR��u����EOe?rȸ8R���%�B��-�5�Vo���v��x�a�����Hq3�ao3JC4�u3H��'���-�B���y���_l��Q+�y��G�8Qbf�������r=�0L��eY���T�iJ�ˁ&�V�V��!����+�]�_5B���Q����azh4�IiHi�����L���-����|.�����jE���ٽ�/��ț�_�H�D�pʜ����}���hM�(p�d�q@�-�bй���ŦɛA�w[>C(�ww��|E?����E�^����+o�!N!�g,��^�����E��)^��L�u ���>vg�'kb���_N��j� �ZsMqŎ�[t�R�]�_�w���@7e�I	�Ί~��6�#��}����?�وq�X��T�^��.��s6_��<���zH؅S }yVk�ro�� �t��ig��D/�1�6��	�1�_�yb��iط�T��z�~�>����R�d��Dz��R'�Qo!&u@���[������륮�s�I�Zs�	R�H��?=�'!�����{iYo5Q���3\L>nd�cˁ��}0�e�KAU�&�ģbBW�QCG���Y���}TЗ��c{��ȕi6ړpػ.58ƚ�w�x�w���� ���U�i�3���X�+Ix�${�*71��y��D��x7��N\W;�S?�:wt�\;���m|;fW:[cՠ��5>�>5�^���V鐖��]������W��6�� [.{A���L�̆=�f�`7Ќ���/�( ��>�(JY�w|�� �
!~1!����OV[���>���ޢ�Kz/���? È�c#3��R؉摮�&��7Q͸�㋎��=^�D�x��p����o+:1[@)���ܱY�8�ݛ�,�e��sp4��qlw4��v�Z��']I�������*S�RD�0I�I�Y˦d���\0Q<RzMM��4�!@�(I0��lY�0w%�I$R`�ME��:��=AD��:|���H������FKrW �,��-d-N�pnw�����f��eg���gv���WlbÉ������B��8mP4 �ۆ#\��Fϭ!�J�A�>�z�S���y��O2n)�d)ާ3�qi"(�fG�'����������3�@��*n���W��T:V4.��E����y���1ƭ�c0=��G����V��w�|6v��ϸ�!d�-5;ai�d���5F�n�G��?9�����?�U����7�i�҂�ʼ�G���?�=UB.�+�g�&AV��Yk3�:��wT!-V�q���a�DF�x� �qQ�T�YZ���ׄG��B�FSfح�Z"̎�ڶ�* &�ÄJ���̨K�_E/>�����ۂm�m��M��}��An�*�z�R�O�����ٍKƙ��e��[.��~�xK^���w~��?�MB�$�<�nV~^F�1F��?=���R�Ht��3�-h�5�1��V���g�L��{�`ޡ4���gG��V�w����|v����G�����~�N��|�"-�����)��G/[��sҀWu�;,/�勺=�F�=t����ǵ5tY�m�"]�"��r$*���8 E��yƣx��c��>���q.��G�F����Ƽ�G,��	��no`�T�"�i�w-��e�O1���f��\�CW����r���pj������i>и��s��9��'�Vf�̼��_aB��|+R�޳z����4�«���Ա�GIHzn�, A����wyM҂Z:t�$b\�EBs
fk�h4�������e$�}�'���Gwq,�&|: ���ɪP'߁J�&,���́��T���!���곢����-\�u��9 /Y0�o�+ʍ<�C_ ����cKמ�]��]�?�ݿ���w%t�����<�E<j?���9o�|h3&��)��ni�<Zף5})C��酊㣖�[���}Z{�X�i�3?�aMpM54߃�t� DB�zA_�-�Vq��):���0�/6��^>]lT��rG��0���Pb$;1�ɠ�ܓ�v��h��W`Fܖ��X��_~����	� 8�_šF�H����Ɇ���9�a��rܭBt�g�5�+��4w���Tk^F3��"����-;&��8�V_�)P��CJ����Z�g����i���W{~mF'hD�����ͧl��c�q�[�~������f���b�5V�h��96�:Zz+q8��L!@B,tA�7Oi^�$X�&'O�
���5�����@��q�P\�{m9;�yF�s���^�a$3�-%��p�/�U��2&B��b�_i� ��vl�Kr2W��2]�".w`׶��`SYٜ�F�>Q���H�Fg�O}[t�r>_CcN�������3�K竞qC`u[a��!%�����b�9�[��ڋ�x'd�M�Gޭ�LE�6H6����p���W�O���:���+ȿ�%�>��
-��|�0��E�.��?�p�n�O�U+r^3�U�v $���-�)Fֽ���:�LS�q��9FaG����Y9�L2q !i�<�I�p��4���D�����"0r�zg�vV>
g��0�-�gP�0R�ڍ��!���)��Z���*��y�'�{ec	���s�x"#3M�#=9�@�ҿ�/)��~G��++������av��h~MN8�˓��a�����B�L���	$pD�B���z	D�����V{�1vݪ�g��| �d@� e���;l}Oww����$Q�Y}t��DP9�If%�8L��W� ���\�&��)M��}b��e���5��W�ߺ������q@5������*)B�q{ }�M�-J*cU�<�Yz�쒸�P�l�@_�0�;O�KB%���všoW�8���	g�5��ȗ�Bd]���HN{//r�stë{��	4*^ѭP��n*�G���;��[	��kP�)�Z�L�����ei�[@�� ��y2Z*�}ȗ�����1-�D*�zH �B��a��)4�ŨJf��Ӱ�A-s�����!��'�0��詀E=}�7C��;l�����Rڇ&el�H�m_������V�;�O��}݋1�4�٢�Q��ſ��x^�@=�h��nf�xa��+��2��dU,O��p�ŻtQ~w�'�g�{�c(l�,<�8J�S��WJL򑫑�S8و����:Y)��ݿ�]{���,�[a�SY5\(�����?�D� �ťր����wt|��;Ka���V�-γ���:�28�l4?��(�i��w}��#.G�(��_Er���Q��bƺ�Z^��O�k�"��A;�vZ��O�Q�ݍ��D'�P�����z���hzY���<�+%F���m`?�3��Tr`}!8��G��T9XTWn��������!E�t����[<��<dm�N����#�<�$�=�v��\���v��I��ȶ)�"�9M�Otm���ՇT�9)f=0s�KS��p�������'�W9�쑨qJ�a`���	h���V��Z��~W�#v�����w0P�F5��;	�PXi<�8'^�$�[�f�W.ʯ�����|rt�����W�>ع+H�D��4�J8��^���n�e�6�g�b߅��fg������+%����q���qX�:W�oйy�b��pD	��b�Ȧl�"b�'���"��١��m�/�a@w���Ky<<��N���1�P#������Y]��A720�wγV���/x�� �����|�>����EZu
7H�L�A]�SA䊛X
�∞����}�z�_�D��$f�6d�J�uu!Q�($p�|�̫�����V�(��~�VZ�_]]��n�+e��'���̣Z�~��c~��A���V�j���.՚~�������?�$�MC����?��v�09~m�p�);�fʴv���t���y�(!M�5������Ѐh�%�y+�[��K�(v؏h��B��>%z����ͷf0���e*�������SR������I��"�yG��N6��.ׇr��b9$�=p:>�A `/w��bo#�L�6S(O_������h�D��׍�ٔF��֥d,~��#m�%O���̲d��[�[.D�k���@�zO�'q)pdO�;JWz�Q�!�rc�u���~M�Eʕ����иl<�GF��k���1p;��?ob��#<(;R)���/�(�9��m�_�!ALh!���|9l���ʃK�W�o��]Y�l����%+�.�KT��Xa��\�"���ہ2�AJ�L�Z��c�� 8�
	�B���0s�e3����+b�MDMrE��m���H���fA(�z���T�qR����c��
��"R��.JH���w��� `O�=���,�|!7�Xt�',>���G&�[�r�oa��:�p���,���I�n�8��K'�y�Z�������EmR?}v�O`&D���xjϾ���Us��b��*�
~�M�]����1 ���VT&��^�J�s4Z���t\�Zk��(R���Ӻ�Waw�F"��u��3z-Xk��R�ղ�+Ѕt�Q.¢J�B�t�8��<��
u}&(��	�Z���W���!gl(u�~�8����~&� �֙r��Niy�S�`��x���`�픷*ڱ������k�E�)�b�܂�������~�l���lE�]j�~#+\�iKM�������&�=�wLAbt!�;����<��2��Us�fڍ-���f^���G�\*1�¾��&]i����ֳ�C��x��f� rN8c�,�;��,��3�I�̱#;���x8Pz��)��,�kw����H��#�����Kuɶ^Ox3]������aG�x��C��d��PeUf(�Y4�ԍ�8
����)��qK4u�����{w����S��i����d�{����v�4�dF|)������0���{j�w��}涷����?�Tf����7fT%�%'�>K��+�`$�c�e�ҍ�>�/������@ۆ"$��v'?���v
�����!RF��l����{i�	;�>}Kz:��#��N�ڇz���.��݃o�������_�O�e�k1Zoi��xz���f�ǁ%FA�*���5��3�ou����yf������TJ���Yb#:f�hW��#�I����jŰ/[�i�r������ ��u	��Gޏ;2�[h#�Cʋ	���L��7��Sʬ�st�F�]E1�'�3����S?��_L�U�k�!�i�MWD�"��t@ZH04cN��QMV��E"R�A�M~׆R$
m��%q�l,f�ы�(�/]0y��D�� �i̑�
�"��%|�;���r��t�m�w��U�����]��<4M��|�^Mg0�e��u~z���w	q�ϋ�%�֠X�H���#�
��h�ڤ���+P�'޽U�k���	���g���ѩs���: �^TG.Հ&=8t�ۛ"�\����8�L� �*'�"t;;^I�{��q'��r^~,�j��tj�@Ne�tIɗ�C"�:C��5���S!��0�_��K��.��LOP�7H��[^@��ސ-���N��$��[�`oUA�$���B�픫M�Qa-�Y�-�y��_���<1m�6����p���c�r �Q�ab��Oj���{u��fwG�Y�`�m����+;����4#��6p)���zwV�G�v�M<��o�qP�b�F_*�v� �6�ai�႘xgϵ���+hᓁ��������w��6d�$p�֘n^
��D�R�l�
��ϲ��)mB?G�"�NKs��n:'��^�j��i&0I����(Z��Ey�y�ɭJH>�=����J��s�y� �]yD��Yl��j2p˵Q�e6#�O�`�~��n�A�&f����ΐK�>����
N����_��C�=`���3) Dg���fE���������D	"�en��T���$Z*{�k�� RvI��Y���a�C���b>i&M�%����F��܋r��l��WK܋i��t�Ş���	!�港(XwLi.t�A2Rc�`��1h@�1�^�#�<���X|q�b[dr�Os�i�[t��{Z�psM,cr&�a�#�ubj�Փm����g9K�w_ ���қe�.���!e��Z ��-�^z�/ �Gw���uVuP��H#���?L�39Kl���H^��ܓ�T�D�8&_:�y�����I*;���(85�&�|�Ea���-Օ�S�o�z���e�*'֠�$ܪa�C4�[���D=m �_�n��=��Qv���FK���Dt
v�5��;��2q��أȜR�\!�+ ���R�M�9��@N�y��gv�e8]��~6Ux�i2���ŉB*`�E�b���G��c����ˆ{���&�D-�gw��("O�$1����؂T&��;���ʔ+��]�<���ؔZ)4�f�J�r��JK(p���K��:NͰ*/����۫!i�mfX�	!�=���䵞(`7����k�������b�f��[ [<mT�w}lA|(:ko�ǘw�A�Lc��@�ĩ���Ĺ�*n|�����ʃo,��7��E��ת�JEȑX��-��g[=�Xe��4]���=�O�`<'�%����l��R���o���2+�'	�]q���0չ�t�
Ԉ�ᵤh����G�0��f���^�ZUh�f1��8���iR�Ã���dG��ޑ���G�=F���d6�� �,h����>�^�G�6Lu��V2�@�ĕ>>��RpX4Zb�G��Y+��{��4PK=U2y0L�����}zb�:�t����9��K����1qh�z���ܯ�oϲc��4`�>��]��`z��>ȸ���xG�V�b�'b��y~��oA��Ɔ8�1��u ��G��~�Is�f;�����J�ș9�ɟ��#ΣSG4ߢ�ZX�[�g�U!��%��*r�3"X'T�� �zQZ�?7m���u�ġ�ŕX9 �l�X|,���4$_Pt�&30$��~���+I�����C�!��c�DҁS�M)ĸ��-j�>Tj�k��8���,�/�a�_�o��G�k��d���>��J,���Ff�G��t��h+���T���j��V(n%�WO��*���qz*�X��&>�Zpk��6�LS�f*_�:b�ug�ǖ$]�E����+\��:L��)hJМ�ބ����槌������0�ޫ@sx�L_N�c�=��z�mi9�_��{��W�9�d���k� 8�l��>I�)uE �wj�&INJ�� V;x#�d��[rM�����>}J$|�Q��L7���.QXd��Htu�u�b���;]D�:����S9'�:�����i6�V蓽�)]5�G�9=���*��x��#�wG�C@,��/� B��Q��	й"��wxs �M�yd���^9]���P�L�ȻheS衋u`Rpe�p��>�gV{»Wd��t�y��S��!��/�a*����.P��.�yא��oUj��``ߧ�� 9<S� �+!k�щ�Ltu��q��h "�BA¨91�a�Δ���9�h�K�LL�E~�'�R]���Y\C�*}=��C��z���/�G�G��4�|#R�����8�+���_��L��4 ��3�J%�[�_���YluX���m��͋�H�%�����o�u��wܫ1���Ą��3
�L!8�|�Ki�ʐ�����d�,DE1����f�1	�(�C��R�FR�c$��!���]��7�d���]�L%2�ȇH7���Ks��+�c�E���%bw�D�v�$0�U@YІ�9-=�R�<]�҇u��>���ꭜ�������&ҍk��)���H�q�qj1Y�$�`��/b�_Z��4&p*�Ҕ�q�}��,oj���ͨB*���->[��k�r��ߒ�X�x��`3����q�ğ��W�o�5�a`�f6�[L&�ra�EY��V����10�ʲ����m;�����z�7ΘN�!y^G���F��	�W$�F���ȳI�G�F4��M�D��;�����5��j�TU+�v��n��x@���p�\���I�E�����������C~��
��DM/�ȴ��G3	Yk�s��`�(����R�b�����^:�5A��4&�D<ƨ(��w�F���D7',�&�p(^����V�kr����ݲ?�� UK!Mw�U��6F�&���'ؗ^{��z�o���]��ޭ8��Z���i�.vg��6���]��ӝ��b���m�����޽���ߡd�!��d�u+{�z�YI�¤�M+�*���3���*L}~ڷ��(ϴ�~��x:�Dձ��m�ʅ��a����ؕ��:3N��
Ū�s��o
y�- �
��U�9'����DE��f.�<��Ѡ���&�3jt`ï(�He���a�����E�Ll�]�<��ZkY{{m]p$u�]�^��f�ݍ&!�p"��J6�e�]=��=QӋ��o�Xt� 6��d��6�o�!	í��>��di������Ӽ���ɔ��x�V��ƞk5S)���e �~@�@-C�d���җf�=# �v� '��&�rD���I̚$������k��Jm�9���	���C[&/�tG�|0&����&!O��wM>�'���m�'�jW�2���0�0�}�ֳ����w�(X���t9�a����9�xMm�R�^�{�oE�b(*��	�.7:G�#�pR��0��˄Ŗ�N'�wi͸��Y�ps"�L>}�	j.�{����w����s�T�NPy�(�!?9u�ώ����,��ݾ�&\��o
5?�'���q̎�ނ�!T/����r0&Ì'8�Y�J�-`v���  �;dRN&{TvQ)�g���RʲHU�M�F�=�0����w�R����}�lZ�2���{��]<Ia;j4�8D��|� �-v)O;�Ρ.՝$L��R��HB6*WU�P��AE�K��w!ޖ1%�����;�E��J���J��˜�\R%v����Q��%I�(��)�3��n���"��	�~�o���>��3�_���;Ȕ��rP+�9�<�U_r�I`G|F�TC�Sk~0�����W�/۳��fO8�D�h;`�$35e�4nƊ�a�n+D��O؈EB�B�U���R#$g*I�=�.5�,�A(����v����@o�<����]�~4�[���Es)��m�]6��G~5�-r=��)�Iz���*��o:֘橺�#�.��O�-�"�?�J�f����4�Q��/qc���Br<�`��m���3�����Ƴt�;5G� �u؀C�Y�o/s�*��Ovdd~!���\�����5e�}�%^��j��*�~�f�g�����
:���V�
)k�ڄ�H��uKB�<5�A@�W��*r���"6>���UG�j[a8� '��1�����������p�uM~����yT<�u/���DcLX���T
�~-T�*�);~OX������#�Rb�.�����D���p�;hׁ�ǹo���(i��83`];��L�B��Ș��9��y�U�ϩ�"`��N�dS�$7[ɝtjJ"F��D�Pn��{=(5�p'I�����6/���o�
ѧ�ޞ�� ����V�<�~���z��Yt�$sK٠N gS��j�7�(�?�~��b\v��,��Lf�Ӑ���<�����䳸o�BCڌ�BbR�7r���/S��SL���ą�wfz��� RA�,���ᆜ���(�6�X��j�x��{�};v����ݞ�I�_��ͮH6=��d�`K:����;ټRE�>�l�;�x����-�Q��+1���W ۩�@�Y���G��S����sV�"�2�,-2����&t�������V��Y���|g�hN�y���]?���4�������[�*��gX�~F�"ʪ��u&痈�Tt��!pzM"���`��*7#2V��/L�� ���E�<�ix�:���7���O"~pq�.�np�J�&��=�^Y���7��
H���+4F�Q+����d���c|Ʃ��}@��ÒK�MPO��S��[�B��\�ĵ>7)�f�����Q33�&�/5�@�y�e�J�_L׍{
�IZ�^�h]Vl���b�L9������sӇ!T�l��"���<n�^�B��A1"�\�n[RT�w`���uxҝ&�$�f��l'����FD�C�5�+T�t��D!߀9���iY/Cw^K��W��4����3�+ލS��4�@-jT?�J��D�ݓh���Ȅ��n�����^)xCh7|�_H ���t{�����b_v�]?b�(Wy��A�q2E�W9'��ޔ��[�= ��Mr/A�4�E�>��]P�Ǎ�C�W7��>�#d�	8�G<����"�M|J2�EX3q�Uq����)�`3	�$`����ƍ����Xt¯�Y�W8̽p$	�f!Aq"ǟ$Ee�9������,�{�k�T���C	�I�4<�羣H�(��#c����8�C���U��ɹ�1?�-�a�*�1��!n0)t3�D@������3�@͋' 8�l����,,� +�+C����[��f=Z������%d]�k<����Y�"�ꬾ<�.��p���g��^J	���_m���&��h�>cD16ѩ�~�Z���.W�+a�^Q��)H��I\C��Y�Ĥ���0RA�4�,��`}�+&� W���d]K��-�A�jGJ�S�m����H\O��gP��T�Fx7b��4@��`�r'���7����ø�$.'q#m��o��T����'�9����N���Hc��~Ε����\�����������b��$�,����A�X~x����l?���(���.F����=j��=�*R<G˘0R�c��sZ�$������Pa�-��X����ˠ��PS­�vS�gm�M]px���ؠ�O.�aG����qn=ߓ6k�BJ�Bv�y�Wlv��-ޔ5�*+��wUu~��R�1|4��GD�z ���e����L�y�Ro�]��99uK���I���=�J���_%0 �ތ�k1�8g��Q���č	콲`��i�i�yZ���gz�W��N=.��Β�j�.��:�%�����������1������B']��su��4�A�ء��SB�Q\�KK����B�_0�%���:�+��-&	VK.�םX3@��C\D��[fL�<O�N��9�2��vs��b��;�W��s��d���.����N� �M����YM�� ;Oko��yP�5n�>�r��$�DE,L�B�v��q M�d�N��q^��Aw�G�u^%�t�<�	�~MYbG���*�+ǂ�j�	;����HF�ĉ+}�s�~8#z��-'%K�6�Ѹ�eP7U��	G��(�~@)Nv�����-�=([�*����C���d�b1Ho����O	f���e�����A��헧��Lb���q��nang�l�)�z{�ܣQn\w$s�<"0��*��Ā���k�a��?](�j��x�975m����,'�Y�K��±�FL�L�+���L�Ѭ�2�k�#z��Vt��i��b#!J*�م��_unw�yq.�»�Kk8�$i�zP��:���?�z3,å�~��c0�H"?�{�WE ����`a�%i�<Ih��J/��ە��,p�E�*�=�D�o��{��>d.�)4��M�UL�|���be�h�<��:���M�F1��3�rv��2��+�BӤ&MM�J���/����V7�$C�;M��@�'*�O��z{��p��]�y�3��/����ӡ��n%D�Q�Y�0�r��sA�j.�L�&�;�����nω�b�C5c_hJ��{���}�v�U�S��6S�h��b��E¥����'4�	B�ɺ<f�k�;�@��R23���!Qe��r@��ӧG�<I������V�+���	�!ٲI�A����T���)K�>¦\�I'�i��Ε�������e��R�%_�b�>D��F������קM$6�T��^r5^[	����y��,���7R���;:����02���2�[���']�ُ�ёh�Z�!y��AF=���#����|���[I���]���+B(,��U�~��-NZ�41cT��]��D�)͈ű}���8����4_h�C����m-�6��Z�N��1�-z7]'�v]�oѫx7�P�MB�W+4�K�� �[9#�.߳�q�k�����aɓ`�9�]��f�>W�7�u:]sP&���e���a��f|=�ڔWq�f9.'���R7��ť�"AzKl�!j�u���& 7ĩ0g�f��ocDLq���.tLj�u���~L�\.�㲟��M����D�Eo´ڣ֛�'��(ߥ�gNB>�R��X���;��|H�#M�^g�P7���	�����6�&/$�ŧ��Z���7?:Ó��b,���9���k:��<c;L�����}?��+� �.�D>{l��-4��WB�`��LKui{�ݾ*��5�P�5��B���zPj��Y���_l��LC���+�Q�(�rq�� #q�9������Z��8����ϑ���������?Y%���+��X<*���R����G����ʜ��fv0�Ə���r0s�q̝፯t8� j�i}s�AҶg\�{���xm.���Q)0\�'zj3pzl�,z�\7�Ί�(�Z(0b�y�D�/�>��傣�a�7Vmʸ} �g�BihL��R�-["��ѹ���'��i�{�}��v�k��"��q�5g/��'d�@�|�]�纷���`��-|�y�4-�6���p{��)X!	��q�9��{>�L0�Q�a���^�[U���R�в�iQ�%���>`��N�\��j,A�c��@�wy%�UPٔ3������l�CԤ_cD(�����t7������Cܹ8%<�	<N���fB/e�C06�g�Bn�]&�9Ab���,�P�X��Œt�/��&�hW*�܄�P��0Ѩ-����?E`����W"�l�?��	u�z��Y�����j�Su9�v���ۤ�s�����<j����(�����Ή�p8ia�Lnǵ�R�Df�&����
D�ʄ.��ou�&���kch�|�s]��^�Hi���eˀe��޳E�XL5J�r�Mr�z)�lL�jt�jO��1��#1	D^f%�G����ܨ�I��i�܌XrJyukNK���Dx�=~���ӾT�X���3i�i�܅������=������4�)�U��˸��}y�H,�mJ'A;�����x��=��K����jqn�L9<݃AW�:]o�>E�I�#$��:�+V8f�f����~A%�Or�J���bD}��~��1�|N�1��Q�ڒ�4���ŉ����mV��dE�����Y�<�*�b���+���/:C6�*����x	��d<�J�����z�L׺2�+E����bM��b�C�4	,R��q! �X��0�߮0�*Ҵ�rg�|�t�����8,�x�_l>�mT��?T�!�4{�CG�E���*&{�ź������.�Z��{4�D+*,�C�%�KZw�ـeQ�G�����b8����>�
뤱n��z���F���ZZ.߼I�� ������_�1G���VA�����H����oQ�L��.�I�k���U-�e[�=\۲�aC�z0)�O������[{>ӡS`�n�iK�\gWݍ �7�!c\�v㻷�� 
0�������Ӿ8s��o���M�_^� �^��hM��t&F	�: ݻ���y^��<97����+��1��ب�گ�gd��OL)-�ii�8��L�����^Hh?yN!}74dD��8[�}j�:i$R'z�R�oxϕ����9���-ϱ|F�3��d�#�V�bgz1񪇙�]~o��w��/�?�&�ۙ(���x���_���.�j���)���xjۭ�=M�Λғ�� ����P�"^Zu�v�0�:ռU��I��]�v7Ϝ߸��-���}��,�F�}�^*Q:�xa��m~��&>�X��-,
�����r,c��1�ԟ�"#4%��,>�k|�s��U��fy��ŬMI�y��4�*�ˎ�z��\�i��o�P��8e��\�<J�h'�x�(���[� ΄��S��4�Y����q�3�W9o@�I��a��\���+��WyF�Ȟ�6~R[�S^dl6R)��/$�BT��|�"��ak2v�_��7���hĨ��X��p@B��ӛO%�ݿd��������(��K�DE�e<FZ~��&7	���}��KD5��
&�ah�y��U��I3ŋ����� �>SG���%7��oO)��:,�A�';�!�	�1�	��uі�Țf	AB��J��^��ûX�l�0���$K�9��M�^n��*�7��P�ez��9�`2I4��F�Ա�g;E2�c���O�]�h�٧qk��˻��苸r�{RԤp��h���͈��Ҁ��t������%��Ⳉ�
���G��#�ho��t\�6x���R���	��r�#�P��v)AU1�^���z2�<繪�#kFPP����r����L�E�7��Ij�Dg�s���u"��D=�G��T%9�#{��o�{�<ݻDV���;�W�{��7�T��9����Y�����!�ӥcFD���kx:@��z�g8�=^��+4��tqD7*��~����b���ŹT{���T�o8D����k0�ى���uz����|P��'���F�Ivm�3Ft�ݫ����!*���( n\���qɇ���a�#����i���R��֞}�����y^��&��9�y[X��\�F��evzڪ��bxef)���z[m�I�x#�+̖���9,E�!a�x2�C(
�šxX_�%U"�6��Anҵ�,?Z%�����O��x�5�b�H��!��Ĝi4��2j?�Y���7��C���B/���a�ǂ�qa�L���l�O�w�e��;��r�r@��o��w�5�����TE�=�Rt	���0��>9Jl|������L�����t���[t�3���u�'+�
����m�դfnA��������F��Vz�ȼ��aۂ�ѿq�upK0�����������a�U�^�[��l�|8�߯'8`�=\%�;D��@Ȗ]�Bx�1�F��U*���+���C]�K_K'�O�)�z�8�
h���|�E�m/�D���ף:<6��n�g=)����A#�~����U��~��(�[�M[E�(T�^���
���y�o+bi��C��6�h0�V�ӟ�1�̌��^��V|לSH4�:�7�#TܒԌe�ء߳��?F61a{�����JX�É����������!;�y�6�`,9�U\o��jus�� "�p��a��e��v��4!����t�4�1`�z*�1���!G��0,����k5���l軞��#���lZ{��w�}=��O��_$#�{�V�}����w,�!6[M
�V����:x�M-!bϸ��t��w������c�L�Z�Y�4Z p�K0Iuq�=k�R>�����T��س�q+��Q��S:6��믾�]�~�G{�2S��ɂ�I�YM�Mڵ!P�ú�0s���>Bj;�C[1�B��^���,R�1h�ė�y��:���5�@�q��>� ���]Oq:s ��8`{���� r�v�������pO�B��}�m[h�M�W��X�c����g/��l�qiҸ�qk��� ����	�0�ɷ�f�e�TZ1�r�~�3��� ��3)Z6O��~PD��j�	����N��V1̪na�wU�>�H��ۍ6:�F;$	�C�E�Q�����ؾ�>�SW�+�P5Gg�8�x�`.���N_�fV���U�G;��A�}�T4fut�\(�u��sH�|Y���*=5=%ٓA�����}꼓(�g��֕�7�&e��Y��4�v��y��@�JtM�f�Y��8�����l�(J��v�cIu^��k�(�m���y3,�*��)(Z�[���(�VRj[�H���`���)	nF#��&�3z�q�����ה�B�O�g3��Ģ`e�+0��U�����M�'�M�,��y	�g��~ϔ�X-��p��^/h
��k��]���k�ܭ+���X���Z"��>�p�M�f�h�jbF�n`��**]�iI�ȕ���#q!�0�M�>��
WܩQ�\?k�n.����u� �N6_�=�ږ��Dm$�d-�f��D�+�������[�Ҳu?:kMɹ��?&�
�:�z=�=�G�t_,�	�L���=~0V�~ZdН��,Q�5�q�l"ϒ���0u�@��xh�)�w���Sɳ(�!V��A�1@2��d��G"����$j�a�a� [�o~#�*�2�C@����"�E$\c�bޥ�;9W�m�e�U�R�?�BWW���f ہմ���_r����v�0�#x����ι�>R �h\����h�|\b��i�|�7=o�棼A|{�M!�)��3��Q/�}r����v����_�~i&$�`�y���Ka��'������^�UiXV�(��Y��v�mk��=x8�G6
�+h��j�?��p�f�d��]�2'a��X���>ٝ�]���e^�6�K6.�8��ˌ��=5���?|��8�:jNL��e獗�4��N��2q�7Pȍtb"�`�۔�0d�
j����9A��3Q��K+m��~C�� SkT
uc���q��g�lO؍�Y�:/��A��%%M>���U֚Z�:���L�[��OMg�GIE=�
������I�����=��jPFp '�4��(C��d��b4��4���� �QV2ۆ���AH�d=��은߾���YԎ���s"9u���M��9:��h�-'S����N������R�Į�_w�J`
4U�5�(3�� ]%(}�j�׭��;;�j������D�����C��T-D�Ω|q�lX�$���c����Ź%J���6�a��?ړ�~�/ļt1�Y
��؈��l�e5���lVB6�a_z��F���\g��J���?����׿�L�ܸ��H�j(��J0^7�m$���&�p�'^��%#$�J���������~�US��h�9���z���2�=W|��2|�^����ԶGC��]oI� ��X�.<�z=lLGx� t���ݫZ��ȩZqt�FU���M$��"�^��F����^�RCr5%��l,�ڴg���m�nv	u=�=�7E�F|� �@f��n0e���L���ҫt#�\��v�`�O|���q���t�9r܄A��!��IM��k%�^@�7@J�H sG�b�X����f;(�+bb)�0��H�B�A�)�������
ѿ]"\�ܬD|�A�g�����1�ϑ �4������L�5rF+
�4�I�'^F��<dPǣ������s�=��Y�n���>�U�_}��'sX�1�߾��h�G��k؉��V�
`;�����G:v�%09Tu,&�mŭ�G�!���3�(�5��3�
ݵ٪*���UE�O̒��-0�`'����L��p�}��`����)'�T/������ߩ��b�}W/����E����Nɓa��I�;��x.���F�􁓒�	����br-q ���'	�� �d?�2�iXB����V�k]E����`��m��T��\���֋ }��Ѭ���+����k�L�z ��[�I$|%HZK����?Z����XFb2})���`35�+�ZF�d3v��� 5a�� ��Ou������M�
V������㐎. �+~�����	����<�[���--s�y?��6@�d�M1@�H�H�UAϭV5�\�Ms���FF��)��R1�����Rz[�wy7��u����呼ƕQ�K�n��@�����F� EsÕ-e�1t��Yh�Ҫ��[J>�]�[$V	�U�Ҫ�A7�o�s�Z�b��, ��Řی�{f$d��Bӧ�p|���:��' �D�]��j�x�ЀCf�_�[��BTfD������V�Rͺ���Yhhc��
S�}rB���)�ƪʰ�zJ��1NɟjX���{8�&����r����0���Fq�\�1��q=��A������lS�6��u=N�Q�u�.Y$x�$P%HQ\��b�d��u��|�ؓ*� �eDv>v�M;�#�&Z��(;H̳V���j@��yd�$Lf�3J<_:[�����D�q��$)��se������L�d �믌�6ز�2b���w�:ѿ�	���;�D��k�.�a߇��T�˂�hq��ζ�6f �>}�(�� �+�߂���ˎ����՜�*��k�-?pp:K��z��� j�5U�V�ub�"��E8���E���t#9��ص��.�
�6w��2Bh��g5����r�yw�gR!9х����N���(�ѱ6Z�탦�E�z��T/F�^��x��8��si'���oh0��"�:�z�����;��@��4jԫUշ��+0�aQ����0$����@���#2�f�f���,�m�x�W78�N��p�ޱǏes�v�{�S6x~���a�{=�{�|+)�T{�(�PWYy�W,����=���_�4>(�1U!&ғ�k��Of�W8�?�l�߳��
�����`�%:Z���#@��D�C��)
C=�l�-�ۮ=���n}?3��ֶЫ%PA<)N��b�]�)u�|��7��i&K,���--��5	T��pB�Sj�C{@bڴS"#r�Q�k��}1X8��V>aG�=�y�Ȟ�����6Su:4����ҍ:�7ۯ_�=�І%B���⣅�t�L5��,?.U��ӎ�|����*W@BL}ˣ�pK��7���]�b>�b�����-d�B5n����9뾦na���q�5�Q���]u�kp�|�v[\p��M
ɠ=�a�fWK���G�*2G=�v�>��<Z^��i���[��5x�x1�ܮ�xx�9k��n^�h$���(��6ʦ�r6��U7��<�N��zN!IR��s���]�f�=KK"�y�^��/�����1�y�����[��y�S)� ���[9k{�HJ�*�߄��4;�2�夓��Ӏ^�Ј�E>��j����*D:E�f�]�fT�^��*�p)M$�����7Һ��ʊ�?���Ӎ#.�Bף.�h�+M$��	3r�d�B�YW+�T�	�䱦�P�޷����1`��}.�[��7{c��g)e���_u�K�  _&�C��8�!�����2L��g�/;�&\�w��j,Lx0�N���E�jv����$S��Z`jA���V_��P�f���E0�8Q�"Z㏍W�|I>z�h�IH�+韬�4I���'ʊ�����|��%/>WaV25�A������"=t�?�'�:��y��r�9����z1�rM9.C�NF|�Y�Z�T���,��W�g�L��w���dKu���|�������P-f]�0r�Y#�:��9��{򴶆_��7I}�'��U�0�n�\܄��Ȏ��ǝ" 5�>@�|'*�1]��CZ����s��e���^���H���a��$ ��e��q�iXD7�/<��2?(z$:��?�	ұ̹���� � ������BJ}��o0kO��`�R��a�4�2�-xǦ#��G%���X�O�H�bj؆�all���E�h����U�i���zǀ�W�L��.V~�C�5Y��=��ZUsK! ��P/>�Gc��'�FGy���=���5
�d��0�\\�6f���Y\ԏ��&�h�A1�Q�j�gM[�_���n��=��\W͗����_��}�����3~����c4���M0l�S������tl���v'�2c�z_�.:D�z?�� $�ȀH��~��nJ�+��9��o4�RZ�8�;Gd��S�3Qb���V��^���^N�Vw����,�ӻt�� _l+�sV���~�y&�l���u��9�,�'�~)�uB�[O��+�d�e7%���'G]�����2Ia/�eq�0�L�4	�+���̅|�Zu����g�<l2MͲV�"ݫ	^�E}꺭&�bL%��/�gjd��P�~ǹ[�z;n»?�n�}�%�M���-8s��f�||~绣��&���d���aI[�K�2(wUy��otX㼖�ҳ����5j.m������+�|D5'���,��Z�t��R��Ӈ�.^b��ޒ��msR�T��l��i9s�<\�����`�M��WW{�%ǱU�t1�˫�M�uiҖ�ܚZ���uu[i7Y�'l���`T]�c������&ܵ+%L�[��/T���~�g)���?��[O�x����r�:��nQUB;;,���C���Y4���´����!Sl;���筀����=Z�����5 �ܝO=�W��8z\�bE�t�,6T�j^�m/����M�7J�L%@�aw����5�A��Mx����<O��q�H��,$�n�Xl

xn�+�['�z�����O��p�B���ksd�K2}�['��g�ç'U����5��f7+�h$�4R�c�if^��,�ԫ�Wy����m�\)����u���t,�B��w��NQ���2Cag`�_y͑;o�����.�1h,�+"]�Ie����RX.SD�ڋJ�[D�x��zp5 B ?���*J��8�`����&FQ�?O�ᅪV��E��v�@x��S>�������a�m�!�RX��R�k�<8z��!�����;w7����q��ڕ�I�b0�M ����S����/^[ �`i#��u�B�Za��_�9t�=����Ey��FXJqp}����dvg���[����xd�-���iX�Ւʟ忩P�(�ѱ#iC9RqQ��x����g�L�(o]Ujǫ����Y�H�e���������r�mR��D4�V�����^7��Bp�&�q��UjA�Q�4N�ff�����i�J�H�,�l�4�c%�<��|#���8rK37����@�!By8���`~�~S#J�n�"Ѵ~$ە_�H����=f1��pv'sA�7�p��2��I�����( �J\j�*�@��8O?��J4�ٮJ�D�\#J�}G�z�S[|�����%T�G M���p���Sݹ��P��v..ά.%�|7b"��q���8����,���4*����o�`\wb��dYS^���H���dMD�C�-7����A�[Y�#���=�[Su�D^�e��~j��7<�~��2%��L��eHiQ��	G4N��w�~��q�I+�*!�W+I�l�=��U+��:����YW�f���T\2 9j�@7v�b�pj�!"¬�#믣!%�T���6�2���q�]&��̅��'���]���z�l3Bja�
:P�!B[?���Cc��Q����J�'�Ů)0a��X�_�Ȯ�&�* ��>���pL�y��U����6&���ۙ�TB�nBn	�婘�Em�������.ogꚱ��;�*Q�jeE{�fV�fɹ�����ZJyp}O,b<����j�f��s6{�*~��d)�r�7�Z�=��i�F"��:Iv��E\�'� �k[ֻ��ۣ�)Z�$�H�Vu��=��N���:�u�/��Ȗ�� �RA���Kp`�e'A��.J-ۅ���Y�7%<�a�\��;��az�x��L%T�0}mЯ����ЩP���G��b�M�!@i|��@ю����@��2п�ݧW��}�!eX{�M�4��K��uk�-s�.�4��j�L�?������gy����4��0P�GIŔ�G��N����Vy}?��.�&�K&�ڇ@�-0�ȥ���� ���5���� ����(�v#�m���������K�,�^/��q90��P����q6ҷaVD��yB��V���}t�&ѶA廩�41T�£�(�o+����`	�w]�{	ZOV�ZJ�E���_�C�M:�~BYMV�oN��L����&�
��\y�.vqf�Ì`���}��q�u�/��?��ē���l�9���@g#7=a��LW���&w��#��24�?o�����Z�U;$�*p$�ޔ����#]�K	f�'̒BY#IM��Uj�;��̈́�gL���LI�kp ��������F���q(U9o��FJ�>"�J0�;���e��;�w����9"L�ҕ�3�V�JQ1��i��)-�� ��Fg���ܼ��ͦ��OV��+�{�l� &�`P�����!.k���q���a�-��r6��=-!�*ػ\�[�UE����~7���X�}N:l[K�9��Q�_�Ц��;�����Z�omc�/M9�p��O�(�1?׹��H�}}v&�n#e��D�E�(o� P�̄�(�:��������DY��L>R�
(k��(��9�{.����A�xȽ҆�� �Q�PN"%C�N�n`g vY�'�6��r?  V�
{��ր�]����2Z��-�v�9j�ɚ�1��׈[����(�{}Ѽg��ٞ���6߄Ȫ��'����4��xBs�[J�Ŕ�}����trJ��J�N�!

��W� ���:*����˝�Q�!�D.2���G1nVS�ݡf��j�D���VM�_�bϺ?��4�+�]�Gx�@�wT*PL-Ȓ�jE�&��>�:8��.�L���	�������"�Ϝ[P�Ɛ����\�B�Qʘ%5vrT��W2h	��%ô�8���l->�P�'�[�C��D���'��d�����~MB�\R����$s�N����{�yV��D�{�p'A�h�'\�0���z&2����n$�G�@��E��"����8&ѻ�cLՆ��ɸ)cy�ǽ�@�/>�ѱ��d���]�t
U�:$©+,h�]6TY��?@�l/盧rMiF��J�RV�7>M�0���⻿�G�����$����
ob=�z�JT��|�m���p��t��9h�H�Ψ&8��z@��浜	� ��ί�-6+h�7(HLj_vVG����'.�T�<�:�߳'Hk��XuJn9ʎr�D�;���B�
�Uo��7��ZpEjn����[+V 
���h)g��ƿWx��&!���F���V;3;u8X�nM1�\D��ٶt=�4FwK���a���q<6O�<��l��WzD$�B�2r����`AXK(G�f~
��^��+��7l���bzz�CRy�sh}>��g�ٰ�-���-��m��U��㽴2F�v�	�3�>���=B-&Q��h��Pf-1|G�R��K#��{FK �x��|�N��d�,8;���ϰo{Ih"*��k�w_) Լ�$[e�i�W�2TYHY��31T��y��i|���Dnf(R���G�}C�� m��}�4a:�[��II�G��6O�<oF�*�e*n����@�S���}���3��{yJ��I`�e��&*@�8�l��m=���Q1����{H��!j����K������>�!F�8Ȣf�3��0�����2���zUPA�����p@)>n��<�U!�a�z4$��lE)�c�h"gQU�(��D���=	h�EN�0m������]}[��S����|���o����H����{�v����W�ێ���ȓ�����>�څ}�ȑ�Y�u�[���]���_��+(�ƍ2t0�}<�я6��ur���TAU����dc�H�.Z$��W!�Yu���〱�l� ��Qֻ�
��^~s�h"��7�a� C[���
�����?�?k��d��X�a(��$��9�#>-8`LU���Mh�_ ӎ �_-\h�܈esd��o(]?A���vvZ]8�;ԩ�ьY�Y�vV���|%Mú~s1#�<������9��T�K��l��K���9L��|A�Q� ��P]���;�ꙢH�b�e�5��b���
a{�$�<?L9g���PF�w���'�o���[��A�p��ruՋQLԫ�F��?�`<����ţA�B�#C3�ȗ�Ҋ(�t���Szش$;�l��0pK�_�.c{F��E��Fo�V!���Rd����$��Y� ��K1�w�V��M�������6�GN3�#i�G{
=���e��q ��������O:�pњ-�x��XȨ�Q6�e�c����S�-����L�n�����
x�*B���D	��+9�s�&Ԑ�ܽ3�� �{ �xh���Dn�ؙ�l��:>|���&BV�V���d/f��Moc䒽&��D�c|MQ�K\
���%�Ɨ5���ɻyU�Zn_�� ~O��Z��<<
�A�.ht�>�B��)�\BC�`�*��-��2�S(����K)�Y����� �;j�?+��t�%R�
�P������bQv[���n�J,}��Gg�fٴ)��9��Ӹ!i����[�IC�cL�2;��:��V�!�\�+f�H��nY� �2�g�4����ۜ8a�5=*�є�s��d�TK�C^��;&��F�-�_������$MB�2�yDG��A�O�p��ϴ�cH��8�Z&2�}�R���s(U�����2�BAS��Alס,9qv�Y�$|mݖ�΂����w�� ��'� �K|��V��M�'�m�,�Ǎ�>���y��.Zh�U�<�˂�6aS��!H:�ȩ��̊�6˖/��i���8	�-b�/{���N���
���<�djnl��;JTV�H+/�Y����$���:k�A@;\ئ��/�C�'2�����r.ke �#mJYZ=GEu�9`D��yak��@�gZynF�ܒ5j��h�p���@kY>�q��D*"� �������R���YϞv�� i�zf��o�iŴ�r�6�E$s��i ~R>��w�	N��2[A��`�������r	P�z���w%�@�Й�ܢ�������RI�Pnq����Q�� �U�����p����W��%^zD!�=�K_�S�Ԟ>�]Y߶m�Q��R��vu�ĊA4�[v;��S������F�4�Z��hL����t·S����C��u��r�)5��:��2&�]�6�=*�ޓ�zd��l �8�JMw��u��J�2��Е�.��rP����&m��f�m��}E7ׂ��A.�&�R�f�&�g��Ѿ�C���σ��������0�t�o�UIE�<���T��5�ɣ����`H�ׂY�FBGt�]�����+�1Ns5��)��Ҡ��}���	h�r�c��ڮ%j���1�낤�GPUe]��� ��LaJK�ʌ���F�Yɤ�b[ƮɮoA�Ok)c �y�3z��ɛ��(Pz�o��1�:(��i5c~<�<�Ed�����%�<�U�)���:�c�L�s�)k~]����rZ{�~N`?�!��L�{�|�1���\�X؝�j����|�#����b�:�:�d��n�=�,9]adփ���&��ӑ��	R Y�q��k����蝡��X͐�����n�[f�K�_�5:��mlgK+��	}:�j�4`�B��ǾGx6���?6T��p�z����������)�2N�G�)��G{sm�{4N�QvŘ�w�ݞT0�+�G0�}̈́�����`P4��   ��ٓ�U�ʺ�l�/)��)�{�d�C������ƽ�L����+#BM������X�~�(yj���B��M7_��?��dѲl�)P��IE�� ��h8��w�'s��Rs&�
.ت��Ɉ��p��MA��$qE�=����-��
���"Ӌ�=��Ar��2]H����bh���@v�%��� :4������~�OL��J#�$�p*՘�����Sl��U��F��JG�V퓓���
qF|M'KIZ��\m�8��܆\rgYyU��.���2��C�G9*q�q+D�N��@4�����)����M͓u�Τ9�ڄ'�I���h;����#��Cً2����3��Y�TRչ��'t�Sǰ��{�1��F8�������Ľ�̗L6�3�?JQS�GfM�8(Ɵ�8�n���P@�7��x0�κ����Y@�
Q)n��/��;�H���]�:�-��9�������Jvn�vbc���6#��t@�d�#xg��}%����.>j*ɧ�C����_�N�4Y�6�q,���l��J�V]p��n������g3n�0Jmz��BsA��L�z����405�ȡ<���b6e+�g��8:�k ��1�;-H�)T�Ў����i��&f��^Iĝ�	��_q�Q�7%��`%Z��{��^�Ko"�ꘜ���qð �V6e���k�Kn�@���뿑�_.CB��3�{��j83F�&DaӔo�j���<����ut&"
�}����7��Q)*l>���>)��2S���-UM���KC�K�-j/7o䥬Ŧ��*� ��Ӗ��?Q�bGCKx����� &�Af�~A�J.��la��԰3X\���
�1�������S�I�]ޓ[�w}W%�� &3�����F��trh�G�|�e>���·?\�#�� 	�;X�i�^�-�<Mi�(=�,��7.��\�զ�樳�)���=��z�N=@�����L��/�d@�gNj�5���1���. �Q<先b�>Wӱǭ%ɦ�>	��#�K�Ĳ�<�H�0�_�h���^��=`���r�U��"�Ԛ��LV͞#��6,Ë��;U�Xpv�0;���� �r�
���O�+CM��៲(�^�8j���_Uha���S^���73����^���7d�7�O�鉄��T���4���%����6�G��u˟���nQpyٿy�v~��!��Mr�NNDIF$R�/��s<AA$*���D,�t6�C�P��v�d��$t��E��Q�_�O+j�+0���S�gY`�I���8M֎���������"hi���PYu��mݲ�{�Y��n)�D�J��L�љQ��g�W�~��-�f:�)�9wR��!��C<ZC�`)5�+,+L1���QGl�Ib�DF���K̊�����mkm&xg��ع"�������,���f�Xx"��,[��D.�85I@Ӵ�����S���+�f6����)Tլ��s��Fv��?�`�d�]�%
�_lg�i���Gt�,�3>�0w����c�\F(�c��8e�"�m��_t_]�nE`��0����n.v0��!4�=�! ��J?R�f��N���JH�6�^�B4��<޳k�Ǎ?d_릉�&Y�����*����!��)�:��V��[�M������ZCPT�L׸�i���e@��	�4=$�|�cZ-h��x^��\[7��ѫ`�&��'wB�	��x�fVw>_���\\Lr�0���.D��j�܁H
�%�aa>=v}���UE����L2�E�Ț�
�TD�Q��{R���F*��NRR�D6\m��qQ���ԻF=l	��5H��X�@�~�i�i�;���bJM%IĻ���ʌ�5�M��#�r�ocp�݃q2X�u/�U,	��FWP�d�M�J�۟�C���5��7d�,Q?�5s{=���m�a���T^lW,���/7!N���֬��H����j}���④��)N�m�5D�M��'p�iT1���:J6�aT� �1�@?�y@"}Jn1f�sYa*�N��\h
�������lxc���y̏�V�
U-�ZT�L��b�q���&{<!�-���군�\~X4�Q'Cj>�}��kt�aȭL�X\(ɬj'^ˆ31ۓ2'xJ��ӢU���,b�s�Ơt{k^�3{c"g;*k����ʶq}�V�#V8�Ƹl`-NmD�+oA��'��䔐����(K�9�j��?��!�.�5`���i��c�nCrM0��Ak�Vc���$��:���a�]�&�JK��a[�z����G���T����N1V�z	9W�I{
7���ς�}����/M�y"�G)�vLYwTG��C-[�h�?'�/��O�C��H��NK�%?x瞔�3��
"I�m����f�0ag}�z��W3��Vdwx}i�(vz�ŝ�ڕ�B�A�lC9�m��R�~�JfN%Z�TViHk�y�).kӧ���|��+T��Eo�~#E=yJ�����zȝ�L�9$jϚ�"+L���ٰ��$5�+N�����k$���:egv2�ms`6��koG<<0=�u}�����#���� �(�
#����"�vO"˜��#b3��x�hΤ�s9H��Zo�]O�&�B_!�tɥ��UR,��]0��մ�L#��nIC��}=��G3��A<U�;�p�ʄd>m2D�f�El��+dZ�|�k.�@ib�]���/o�c��0!k1]�إ����~�Q����L%Wm��J�+�w��7�O��_f@&����x $�8lA!R�?�;3D�Ρ�10R��Q���LA��rgN��+�Z��`9�����C���k�q=�}�<�X��vt��QI�_P����($ ������t������by�!& ���kJ�*�Lx\��5�D�y��]P�m�փ� ���h�^�?��ѐb����{B�����[&�	F-j��_x�#�Q�)�Me2�����V��aCmz������e��k�E3�N���5d�
D��6���i&A��e�g&��u��RUA�ɱ=OG ���lF�<|9��Y��
Q�������%iCF�ܵ��9�c�`!MB�lԐ6���!���.�C�6r S"&�g��d6�uK��Q�9����|L�?��Y�l���59�����C����肠F�P��枥��G� �*~N�w#�7��H����@��Y�$��b������<��h}t���;�h����Z09��ק����8�Z��bV0?�l���œ"'>�.q�P���RǱ�����Hd\�$���D&��}mץ�*����)��r�!p�'	`�?;��pl�ž���8�faK������~
5'�j���@�Wny�A{+AT�j�y���!����W}��$f�9��{�/'��"�qҎUm;� �!�Z�|B	�>���s�,D-g�(�?OD|Y�5y�WH��>8^�w��5,�YD�I�f��2r|��DM42������ȱ�:�-M�)������F5B��$?��=���~+���z���p�=��������H�	��,g��_�Wj8N[ \ɢP&��OwN܍B��"�Z�K����}�6ٿf^o��V�6��M��얃2:t��~��k2��L�;�`0�'�&&�o�qK��؍�b���O�4e�A��������*@�����H٩8�\��Y��.�('�U:_<{%�ǳw �&=�y`o�Z���3-<�}G�0xx��F� �>�9~�����w���<�	,\$�jpCg��zײ�������ӟ9�}N/'����j9Xؠ��/��"�yWh�N$lt��0��I��,|�|>���$x�5	�о�?Y��?���v �W�1���<�q�o�OU�;o1��l�E!����7�)Sw��_�S��˴@f��Z�h�2�����L!�?ƃF}�yYçw�m��CՕs��zTW��'�w�Ƽ�m�O��$ �D�YJ|����S$�\�z��yg�<�@��5��z:S�G�@tj���<��/��7ff�í�do&�^��qGVF�ӏT@7�h� ��bg?���{��6��`�r�|�EŅ��(Nr�=������^��F���u=_�[d��^�yצrJ�P���Q�����+=����yKr9	B�3�����Cn���}������0^��O�$�YI��$�Yq��;N%<�-T�E��7��v׏�s.G`||x6{����dP*_d���l�ߝ��ʎDy����X�E�`�	��;��)���S��>q>��t!��*m0}���D���o�>0� ����.�2ѣ*�^���NdLe[F%���l��PT_�B�/<1�'�Kql�2G��`pz}���9§9�ũV�Dt��K�f'����j�>ø���ѫ��WHP*1۩:��wrKBw_m�碂�_`����S��}��ra�)�ki��u�a!l�\�j�U�>�Z���#��UN�*mۨ1�����uI���E�ࠊyq�
��f�)�jW�3�#��5�����x���rp�i#�ͧH���Z�6�U�m��f��[�&#�.��ڒ�x�P���m.�ڼ�#Wp{��f��{�~��z���G�E�/,�d�����L��S�o���n��zL�e�[K`�P �_�#@��C��29�G��Qw��X��� ����b���C�E:�lN��K1k�|�T[?�1�ў?�`����
#ΡE�V*�Z�"�rt��!#��@�@���B�;=�o7��3��m�J^��X�jK��z��}R���K�A�X��O�AIK��j^�栆��	�X�����Ɗ�z�R��{����.ފu;X3MXM��u#�`��B�)5�|��y��0���ɛ^�D�2K'
]{S���y������/�ӻ_�?����O��L�U����ӱymX����s�؈ġ���}�D}���e��v�ᥩ�n��Y�ם�2P�`g)7{��$�s�wɳ̽�:����-a1%����>��F�Q�=y3F>b��0�$����B�S5��Tu�����#����U��,�����@�]Aݗ�؛h���m"��jހ�K�����OF�?��ޕ0Z�d><�'��� S	+�{I�V��K/Wګ��<r4׼�� ����M:;�SBz@�_��ʎn��b@��Ȍ���wm�os��ʔW���i��^�V;�����;����9��>�F�R碱dU�5�~�/��[[�ga�o��/�K�<f����\'�Z��;
Ȁ8�P�Z��2(��'u������AG��F��:�<�Vޚ��O�g��$��G;���3�"���홛b�>�b,Vm~c{	���:�βA#���A�409���g݈�^�	"��x�8�QC�~�s �*#a�@�1r�+c�w.���8Ł��p?��/	��M����N���׾��j��������g���qt�6���F�t�R����']�$H�F!��q��@S,��5�i�H'ѡzJ�
Ǵ�UPq��/f�2Ф3D��O����j���W1_�iK�<�^F%��-v2����LrDy�ֈ����E�>o~����5���|�6���0u����@����3jo�|��!�v��d�'��ήs�8����ʭ����c��*@hǌ�r2U\���o��'�Ǽl�ma�2�f-g���]�����j-]�6��@��45�C>C��p��I��3X���s7O�̙�N'����������Ny��=|�d��iL-�)�F�o��4}��hb��ॳ,�
'
��t�>���~�ރCv��U~���腢E���+
t�S��u�W���|�L.݅���@���b�U���q�� E�
'�7���	���O�0o��qO`kt�R�G�^���J��,�q�k��d���V8�J��9%�9c (�߇K]lH�;�3x����c*�`I�S��yqd��(��p$�-�B���z����2�
3F<�â��㭾�\���64���V��t�����Cpw�k���w
yg�U���Z�����U��`�cO:���P��RA������,��2/��O��c�7��W�4
����7��N��t�L)�>DPI��*�}�J�[gh�Oۙ* �����`�%f�����T��޼/�������6�D�j;N2��H���h��QtL��U�ɕ����t��[_�j���5[W>J��p�f�Y'XvF'_��IN�!Y�_D���|OG(Ox��l��$4�]A+ȝ�16 C��)0O:�g�kM���o���G��uX{!�i����I�7{����z#1�|��~����lG� ��mt]�?�=��ș��a_�"�˭ް��e��F�Z(�H)M���?C䪬����r/��B.Sl/E��~U,�9Q[}+J(��T{<��GxKR�;���pd�?��B�osY~� �k)�5�`�w[�̼P�Đ�6�]���
��#|�s#ss���0�p���6�l��U<��C?o8�c��W( ݦ8T��hZ��&�K[35߁t)H&|�q���
����(W's�&�B'�.K-˶*C��f������
|	u�4�/w͉Uc`�.̋6�VU�Q�ml`hmc���VI=����S��3~�p�妧�����5����8N���>�ut$�=Wk�H%�T���$�@:�H�?�R���l���2U ]����
�C����8Q�n�>f��� w��P���7��Y�,�Q�+E��5y��C5�I�_
�����P�)���~���*�>���4_0*�>|+������51ы�Y��+�S�]�۔H-v�2��&A��-V�]Qk_+��U�~��E�8A�H�c��0alz�n�O�y�0(Mخ�V��z�y���8Sa{��й�d�RM>��3���<~���~-��t֒%�_������JS���Z��-�YU����>%��_�~�tj|X�b����J�(C�!.���� �	\���&L�2���uv���egZ؄�\R_��}�/�_�)�<�����v ?VW��,J��&@;��$���(@o7��B+��]uo��3U��%��H1�	����xu�q_#�
�U`�B2{y!��t�	���x�r���Fu�P�1��R�urC�c l����g����҄hYT�(�ۏ�+7-+saYQ/�c	���e����[��T��9��V��ʃ>D�[��?&9����[|��
������p��<b='$�G3t!�q��l��Z��ĳ<�ׅp���q`��)E��.x��G���˽���w���(�J��]�H ���_u�y�ik�6��}�cpC����T�,Y=~�Kj��^qӬ���cȠ{�4��&Cw�C���%B�?�8��񤆆 �|ުH���HX�%��^Q�����m���xq!W@�u94�6���{����%$����1�KDѠ������3�A�Q�7M/��9��Τ���Έ���Z�m�h�sj1�	��VC��bf�G 4��v��U5�үo�ud�u.���a��W��A	�����O��Wf�����k��ڨ��_���̪8A���Z���',��Ojh��?m�	+��*�F`"����乊���_~P���~݁�����y'��Qù#e!C_�=Qq�?�JӚPv�E�G�m��	�Ӓ�p��0M�%��#۳r�����_2;c��G�BCbMlY��׬�gi�1ew|J�L�J�tl��Y�v2�6=�Nl~�^���z�D?II!{$��a�}���Y�V�pV�	���tAv}�;�Gk�M�t0b��YcS�`�b����g�\l`@��W�D�w�F�!�wO"������4�y-�V��	��1� z1!^,�8�z��+2as�sv%S��t�Y5bo�����kiX��_/|TD�fgb÷� uSI��/d�*�O�fT���֓	�`����߬����(�tOe�+���Q�H��p-��kx��?�P[�-�
�&i&f�\k�a�zpr��{��,(�*�n����k=��j(����Y���n5���d{��M� e�1��%�$�����4�~~�20�f�Fg*�[f>_�<c	��e��MΖ3�J�8Z`���Y���ށ�rP�mOU\�":X�[���_W��J0�74��Xɧ��8�D�'��"x���;�#�ڔ�E-3k��=[j��C�u$��َv��X��YN�;@"&��%�'�R¹��J֭��-�nf0~��D�Wۄ^R��[.y٢ �s�?�"'C�x�`a��l^ڜ�8�>	�'���=R����2��x�Zq�w�ǃ�R��"[�mZƨ<��;�n��悢ET�[L�9(�6"5��M�b5��3�<�8��˙<Z�Q�?�C���H����HnO�����B���F|G)?���yI`����0�ρ���L���=~�\2��"��ѩ�����4
l M�4j�i�x�2&��m�Yg7�(�c�m���њ��y*�7�Ź�7k�%lp5�������ؼ��Ü�5����ߔ�oЯ0�f z*c�����!�d�W]��;�����%�!R4�w���A�ĥ�h��)�03�o�gY3���$򋎱�X�Q�5��}T��$:�ENi�����,$�>7г�yčw:EhW����������[e�ĈZ� vBJ!�u]l@i�k��[.+Am 0B�N�σ�h��N���(��ȓ�B��4Kޜ?=sv_�Y��a�Kc0I���k2hh$=/y��
��e�v�X�DD��� �R"�+i��P�Z��h������V�e�E2�����?��f��#��2����77�<'�6��hH<B�a!��a�rU����LvV�:[�~�`��	}x�p�HI�8��Ev�5���+.e�M�q��E��s@�0?=u>���~��P��<����[�]}��>��C��1����w�Z����肋w<3��|o�UӜ����$Aq2및|e�/���x@��
�����B	W���^Z�pd��AF�K�W�e�#,b))O�9���$
 ���̓�=85Q3MXH��)I��3���D���#	vU�@�OD�8w���,�Q5s툜M���DE5��`,�{�f�;�6$�}V��V�:�!Pi?:����ڮ�an�xD��fP�C"HѹR���-+�8A��S�l��?|�M&�, �M���1�t�0�e�O��lA|us����1�,{�-��boQ�`c�[!�P�O�GCn�׵��$r��U$���Oy�o~l���"��$�q�aTB���I�h�ǤUv�A�_�R0^�@[�`M��R��ܢ;�ޤ�i�5a��>&�1��ݕ�8bhJ4	�`�X���d2��D�H�\k]��y��\p':�X$��N��P��ڏ:���:��9?�n R/�K��s��%4�Ȓ����W&������6��c��;�O(!\6g�WQ�|qʹ�,J܆���s.mI(F�8���֜��h�!>��� {�+�#5�&+]�9U�2T���`�;��
�s�����kr�7΋�a����7�%']6� ̾�!Q�̎5��ՓV~G�c��-�WO�A!w2m��(C��Q�:g�LUӏ#K�}~��h�����A�ZH2t�H'�s\P1TH�:�p,�]vw�`�zy�7�`�=�����\�`Ē��4M��XK(	���;�x�����J���%�����bbn�wq {��3Ϣ�F}+fš�f��I8�&�C}��cs��Yݛ�>΂��z �n_�J��ɅPW7;��J�o�	��A�4X�����d����8��m�C�˂k�R���8� ���6&����а�^y�p'T������XNO����_�|+K���W�6j[*����_���J�H�K�zF�8�B�r��I�03��5�5��뿛�9�2Z0+�牴�O�e�*Bq��&����&�%�#{T
��0W�ƃL��,,h�ߚ����xgs9�ՈLH�%�[w`�P��_3q��'S�yh�IQc+�H�f�̧�ఖ!zdp7���B@0�^ҧeU��l��u����mg����+b|�m�gO\8�Vr
�܀��̬����N}�
��Q��pŶ��.��h��LEx抙�o�v7�Ao��m �1m��rr�Y�pPHG�\��a�>8V-�f�@��s�z�, �=rb,�hc�#&���0�o���H��Ba�� F�j}��m?]Ŀ�+���O�N�̀��1�"Ԥ��?�ɳ���'n�G}�z_�D���h��J�7^�M�/0kyteMM�涜��Dz��/�8���6�,��2u�7~�Y���=ҙL&.**~&��K���.\z-����	Y)�Z��F��S����nvf��!�a�V��{�6Z1k'���Z�0�F-�w����pYN|J�3���@�qt@B��R6H�˽	��f���3&$Lӊ��5�_�w��g���2�9�U��
��G���=�&������ŷ�9�[Y�]}n�l��Y�@#xߙ�9�2��TS
-��%ڦ����ps��_#1?qz�wP�1&�igY�e���Ӥz����?����1��u70	�W?&�8�+��p~C5�CF�BZԐ!F��U9v�qJ��kd_ �;�j��� ��|O�P/s(����å>0p�E�@�"!��i>,˭x.\�Ʊ5�M�2'zbm�+�@�z�Q1�3�%V���T�3@�g�`j���3�T�n��	o�,=���ʰ�C�6P'O;[�ir�r��2�	�a9'o���a�I'�w�F$ρ�@_�;x�����b?�߰��UO�c�+�;���I�+�9R�!�6�����2eQSY�4*lD��187�f��Pnc2��0>w��M�N�!;>T:��26y��@�ѐB�:�(�}����bjH�Hj����}�����1���J;m���� +*��P�v��:��T��Â��������q[�1@�u����L�'ʪ�T1ϫ�}Ĥ�0E���9(�	�3_�QM��<3��ڍ��@��ɀ�Nb.�]�OD98H����	�V3U��<�3}M96*�ՙ���3L RM��bW|�`+���(�k�O��D��]|(�(�j�����D��/�#�d��*��`�B�d`��h���.������3Q� W�sK2ZJ%����������
hX��:���⣢�q���3�����EUg�"基8O3�T�4k�͸�
�wC�Z������I�W���Yjn�߿";�e($��?W�>�8�q�6ɹ���24��Zw���q�@����}vЃ�|OX^r�_l���4*�$��y��т�����ʷ$�y=�P�긺������n��v�"5����+Ɣզd ��w��!ͼS��t:����f��p��0��d%d��]94Vf�H������+o�4P��r[7���T�w��6�k�������o;���<ew�����' s���fZ����ՠ�ӷE����/X.D�M{.w"�G��!�⾕��{&J�J*�7*B��-Ԉk��q21JO���)�,���sY߷jHK,�هN�m� R��dL�Z[n��盢�0f��:`f�[���� )<��$̑�f�0�����ސ�e��e��c7���k��������������d�z�Kr�i���d�`��_g�pג��a#�>��{�e��X�-x���#/�~��q*N�����Ni>�x��$K��!�S�H`� ��� ~��@z���:`"o_��̂?~2��:�}�vJ���N����R-S�q�Fˆ�a�Rp�e�;����ʶ�SQ��
}�)��4������g�X=ڔ�Q������@O�Ȭ�I���ô�ġ��-]MBCqjB�D]�wAMs����3��~_�&m�E;�{�Ȫ��������+G�/��ȝ��I�5#�ﹰ�$��2�@���+��r��r�NF�aU��\�*���GOO�q(�{�2�hp�:z����uu$_��f�N �8�Ӊ�]EQ�)��k6����
K����^��YI�j��n�:vG�JO�� �2`��Y�%Y��������y�U�H�zq'Ҍnd��!`$�A�-u�ݾ��屖�lO'�0����_@tu��&CE�
2��n0?�`F���G�[Ǭd5��*�ؗt�̃�v���O�5~�,�d�ne� i)�̬dq����;� ����b~�����L���/o~�[v ��b��-L�]����Qy"N�X���ݮ�zFs	d�v3f�>��!���xc��nCc�ϖ��o�5�r�P���.ҟ[���Iwߥ�x��K9�:��^��F?F�LM�z�t���K�c&����?d�y������eW���[�Tu�4�mJV>�����LZ�f@��T*�x�
۪/�/~2�
�U����gbW�u���S�5�6�7ŔH�/���3����n�kIť�KrMBdx� _ԑ�c��*Y��*:�^�M1*�&���ot��� ꯭�{�"K~_�K�6�I~���7����s�K�$�FV�K���h�h�\��dR^�kf��.p[GU��!>�ǃ*�$��d��y�[�+�5������2v��0[��@�U~b�!@��x{o>A1�Ϸ�
u����aW-T���\B6�LJK�t����/�ER��/����F'&֢�|���/\a��NQ R"d��T������0���#�|�s��_��^�Π'
k����\�굖}�SV���ȑ(�`+D��_䢎?�#�O4G?�_��9�*E���"0eFH�H-r"~?�i1���XS�^�#�v��T�O��o�C�d��ѰX��ۮ)\��龃i�o5��ʠ�(b��&RV�rnOģ���G�pU}�W������7�O��r]hh#x#��)j-�c��R�H%Wn\�`-�ǭ�!#�C�3��aJ�����4�N������#�H�e�^ ����ٕ����l���
I������'�Y������� �]�H�IoJP�w_MT�A�8�^�O����b�B�Hf1;����k��w/I�~S'�ָZ���X��>@��L�4{a!0eW���h3?���T�������oC�A}��t� 9�{Sm���8%b�y+�t�#
0�W�	zi�]�[��Z��+ ������◬h�#��4C�.B� �꟔�]� ���f���CvU�q�j1?�~��<�x�P/ϛ;
�'��`���8�-L^�w)���\��7ؓ1BGOnԷ^c���W��7����HA�F7��(��O��sxAet�F+��7�C��2�#I�~Z�U� ��獱V!4sr[^Q��WP����������8�9?�-$e6�'�����5�hQ��R����Bk@�I�*�џe�\[��Lt�SoQt
bK��9*��P�ϫ˖,�Yhvu{��.R�92�A�nhP��[%>�u%��鿖*j�P��Bo�Q:QR����K��9�ĩ��-���l/�Ɵ�K����;_@���&+��[��ЌK.)FȬ�!	�fy;Dt$Օ�8^L`h3b�׿p��{/�6��[���J��5�l�Rpq�>^��dS�3�X_I���.��qߓ[�,�<�+<4�Tl�����h��9=*��M@�u<��m����.������"V��N%lb���$A�G�6��b�p]@�_�g�\D�}6�\ć���!ٯ%�!ǃ`QG»�=;DS���up���hGN��ƧI<U ��*��r�h�J~������nM�S���l�g��s��$�����<n�W�o��g�FvD��5D�zJ)DA)�ߥAn����h�|4)��P䀶A�>���)�8�@j�K۪�%�Z�(��A���pZ�{UBK'_?�2���G�ZU�C��9�V~�������S[��2xhsq2���F�����O�tL��ߡ^Z@��,���;J��g�끣�q�e�����4���H]�F\tN��3/�4�O�]���i�J �����5w�Ŏ̌R}�-Z�C�sh��h��8�\�Y��&�X
�y��;�
S��3gf���H�g}�+�g�����G�u�/��"YZ�V�+�o��%㤣�ُzB�G��Q�P�P^Ft��z��К���M���v��H��@�wdf�'8�`1�?����l�w��������s�sw'�n�ݏ$s�4�4���`� �v��S�'p�d��ɐ=��*:�F��q��u�K�N��FXT�U��;{��+~hYR�h�����t��<�y��r���
���J*��['�s�V]�Ap2י���p_�����8�:����I�/������<1]�Ł�RU����!�F��
�߀Z��.`�OJ&�Њ���dd}p�vHNA�*��+�����992PQه4�6gI���{O�	�>y�`��#Sxq0";jZD$D%�@��$}�3�ș�|`�K�nD|$ޡ��H�n�U�"�w֕-��9Y�h�e�����Cj���;Ań��irp��gC^S}��h,�T,��rWm��9ae���8�H]�h�>�)��)���ɠ4b?�<��S�ޏU�a~�U$7�Bz�ש��駌`e�>��Tm�S
J��lA��&�&ɢ�|+~�G��:��Ή�L#�ڱ�-B��#'@�V��u1�� ⚐G+�q��ͬ�Z���L���Uß�PZ���ٹs���(�I���U���y+�� q�v~�3��[p7+�I�����PxI�N��u7�61V 9uƦv:�R��q��H�ϓ@ pe�q|c����\����)K;F:`�s�(��H$t�g+P�**���+-��F�����	#��*����$)h���Ц^�BYr�^�	�Yƺ����`_%�o���nM�ȍuN�b��<�C�d��O+f���-y��۞s�U�����M!���\�.�Xo~����9���;�h{���t<�2lc�\�"�ӒbE�t1�~=�4S=U
,�ڽ4��ܗ�g��u�7#��ر�����%�VT���K��� ���E���?�[j�hS~��1��I���H�-��܅��A���`�'�O&^�}$"��I�7f�(~��Q�䬋��S�T�ast�����̂����w3{���	L��8����hc5ut��ç�z��jg�bh�"��c��k������=V��/X)t�81�\�amY�y�+��O�z� YS!+S�.FQ��9�,�I��M#����������I*�HEI�s~3tF��c^�/��馎����|7�n�c�kH4G�6FL+\~3�*z[f_�{���R�a2�\�0G�n�1�}&>�b2����
�2 =�� �ZE����n�R�o���^����z�3�~���æ&�:�a#��=Ys����\x�����rЉM��[W� ��:v��wû��3��`?n8�zY�Ћ��=f˴4���h\�8[�s+�<E�?%+��G��s#��a�g_J2����5��EJ4�6_���*[�r��f4�RDP9�cػ���7Q�X)��K�����4��VK��u�؅�L5ݼII��̄��L֞��>L���f��.�"ݝHWJ	�]-]"�g߯�������'�f�P�qM�ű�a��iz�"���%|�~	!h��I�OFF L2����h�/�G��µ��h' �+V�08�i�%L5��@Q:�k�}`<�ɜ1���<����ˮQfĺY���V�^Z��g, �@�2�I�.�0ٜ��0���đ����y���::RJ�;e���I�m-�����S& �S#t� 7T=�'����F�@�J8:C۲>[�����@Y�xaFՌ���L�e�ں�#,MsY�(_I���|����&�#�u�����y���b��=��#@����b���ѕ�,m��u!l�|����/<��|a�p8b5Z��5��~�r��7���8��2���Kn�[����2�/��|�������.��(f�ʎ�wC�tP�TT�ai?@���#/'�C��ޒۨ�t!砩�E���s�5�:ɡw��rj����#���P
��T0ݴa�V��+�w���֢E�Ϗ���>l�g8�8;1Y<1|����m����V8T�|!��9'�����x�|"`�����)*��:��ݵU����H��1H鴀c�]�J-�dd"V捄i��UC.O{I?��ɓY�9?8�ks��D�������R2����/2C��� zh����(��T�,���$���.�R#�{v���+(���!�E|Q5�1�H�j6;͍
l}��a�dl��2_*O�7G^������]�{����:�E�F�<�;���F���[b�W���Tg4���w7�씄tSbdc�����$%�mj?	r�Y�fznғ;C	bu+-~*�-�v�j_��)'"Y�r\E�rc
����/��A��׀�5��� K��ȷTO)=���C���Br��p�i%n�z}ut��E���E���`K�D�� g��]�Fa�#c�9��}�;6�8�#{���x����NW���t�6��\(�2%��Wf��wP?O)�f��%޴$m��E�ʬY+#��M�#�zG\9�UY��7���;����zT�Z���˄0+,���O1��it�G��̓��L���*�?P��+9����X���̳o�4M��
�E��g�]]����ʹtc0�)�K	9���ý�R]�xUYhq��z�@CMY�'
��6h�M�f<!k�	��~��ŲC�O�݇1�r�i|{U�gQ�[I��,�#�IX�P��*<��6�R���g���s������?�e��Z�֝�y/����_DCCn��T�o���H`X?���;� �h#0 �0�9\~Y]	�6S�;����T�.M�r�OѼ?�����J��[�GY�$���L�=���l��AD�C�
�k��X�͌��j��v\�i3�����/yM�-��G�K���������h� ���T�����!e%,�oo}��3Q ��������N�3C��n�&ϻ�?�t��Q���s�_O��A~�;��gF\�B�(�%��b	Y�&G�Q��m��a8/b��3]v�$2�1��j2Yj<hܷ��oCzԫ�@e�(N8�A?j��dr[�����c��h���f8�`c��Yo���c��Q;l�S��g��*
�a���3�����1�1@U�P�}�T����vZ#Q�	��E/��1�_��'��� �`�h���J=���Hf������+�^U�9oɤ���ƸNvM̷��Ҭ��������]M�0l<��
%�j"f��]�1؛����6M:GV����<�����M�J9���KY����,����UP{9�2c>���cL�e�6�A��(����{#��Ny}�Đ4�L8�Q���������D��"�r:�9p@0uS�LP>��6��VKb�F�L�>y�f�q�^����o'�(>ɽ��ޮ��Ѵ��NN]�'��ӠFn��|�s�H|]2>"�n�Ŭ��[�>��Ϲ=�ϸ=jb�6��^���u/[�,��~�erEm�W��r:���4�}K�V>���
-��'��)�a~ .!{�^v�ڊ�נ
y���r���'Ô��Iɷ+���$y<�6�i; ���K�Ԇp�{�-�����*m�ŀ�r9 +�lz�e)��:è�SBN��3�x�gn�	��.%��hc��;~�C*{�U��LBn�X�@�C�qW1�|6�ܸ֩1v
�!g�K�J���{E�)a�#O�!p�]��mS���?�A�Rf{�����f�Ռ�8�O|qzޭ���/ʏ�^m�2��ɼ�b�Q,/��̕A/kX�Bn]�Hx�C��^/��^޴� /�m�"�.��x������T�QO���TD���5]��ֽzz�[�~׌Rp4��i����VX�l?Zr`WG;�IU�;�zO�͸�+���/��oWO�"��N��Nrjz𠳢�W	�X</B�w�IX�;D��܌��^�5=1�h}Bw��{�J�y+�K2R�ǝ�'�tQ;��X�O�+����UqnV���B�|v���|fܜ.^�u!6� �F��E���Y�(�Iu����_Q��`
�I��u]�'�����m�*�R ��}���f�;6E�Gy��Y��4���9�~zw1�B�nP���F�n1���0O-:+\����I~�J8�����|A.�v������G&�}[\�!EfȿȽ������ї����w������%"�4(��z��9(q��mkG~F��[g��Y)~��+s`�'o����p�7��D�RY��� -z�o���D$JJf�N���=��"7��d�ުP���A�4 �xoeFX�G=n�Dw?ҖS���W���Bl����^�ܒ7$�崾.��|)z�g����������=s�r�ZE�vug�D���i�؊)�4d������;}�`�+i#��X�~��~x�8����FgqAE�8e;��K*g�&��g�7iiX񲔃[3�0��XGO�l8� .�8��$B��@�P��\�ϩ���R�� c&�M�T\'K�Yx��)�qq����ª����QB��M��"g�u���ɇ��e�ݛ�y�A���K�bY@�K�;����a<S��}��ʺsQC��zj���1����PC�N��Fb��(��[ò}(4$A���1�����4� �kp!ſ�iN1�0U5�u�N|�T!V����о�����;�m��E�J��ѕ�Eͳ�{s���H����ゲ�%7G��z�ґ�p{1J�K�����x�^�l$h�goU��{�@��Qa�$�i�����ݻB���8���XűU�Y0�˧�pũL֡e��$��������c���D��Z���?��W� ��Ze���Ԏ��88�x<�G�U/�8@b�w�ϫ� &�`�\Ԧ�9H�w�l�f��v���8�6I�ﯮԆ�������Ul�3
T��/ze�g������m���$�>=AZ��UX��ٕ.5tb�� x�Nk�
;�y:��|&y�?bXg9���W�'8��~��vw!:_#��2~0ǳA����G��tw�4ig�c��:F��:l�
uMaQ����7?,$b����vu��k�|����w�Ǐ5�����N���`�Y9�O��C���N� ���"M�zHvm���_�����=��7x���H�_?�=+��I���%{dy;{�H�sMFWY>2��<�8�z�S+�������� "�:��
����:]սɕ�%�hd}�'0�p6>��7�܉��0�	�k4J�OJ�9O`B>��&�0ߔo�w��}��LO��,�v�z�x(=,�!&Og���F�q�Y;�����3Z &��QZ����ۂ��I�IyW��f=ѐ mA�~��4���ݠ��(�r1F(�`PD�!Њ�$uGc��NsK_f�{��0��*�f���r;N{�Sp�*����t��m;��mEr�S���l<��Vf�����qQP	 L��}�$�_���?8��S���8��]�8�:�3<������ӽ�3_�/H�c a�~O��`�5I8���=�M�^U���/z��G4>	V�����}��)����9QA��
�=�A���;���X���b7��a.�ˀ�dZ�e�����8,:8��6��+��d0��t]������}����#i�k���l��lŧ�}�礐��e�^/�0{�� �
�6�K��F��}{)Y����+T����_Eɾ B�+>�(<.�;��"0��l@��ߢ+d������ ���M����H����e�l�&�V���i�_�-E����+,�Km҄���yg��Rܖz��F��A�W�"l�+h9*��byزX��a�jgp�A���-��s�(���Ս�����"�"�`�fF���e"�03ً.!�LXt�#ʎbn��BHn��Z�&�5Yk�I�!��>�s�"�ρ�;�*1��O�)Hl�(/7�T��I���gA�\a���._���w���1����p���υ����&���Y����{�u�ޔ�7�|�����#"��}�V����ӎ����Ƈ("H�Ip�
߬t�]bT��|^dSn�넻�Z?٧�7�6ax���'�S�<� F7�H4|� u��j{��q\X�#�x�{چ�^S�h�$�8�Eځ��wy��Ɓ�G�Z��9�wF�������B�_���w/�M����'׶v�#&(���w��l2�l����ٶ�XNx`���n.���!���s��;d)�=��$y$�O��7��M�|/�����G�{T��g�f�F��r>�-���f��(r΂�}ʤ��׍�eH��u	6��'��;��ߗf��6�#���y�v�����е;�c_�0���2�T��I$�R��җG�r�ʈ7"!�6`X���C@lZ�(z4���a�9�|��9����U!+E�ɂ�ã�A��@����dB�=���F��rkY���X�j�K�}o�{\i��5 �
�DJ���]�}6�c���_+@d�$�L�]^k��֒?u��:Ľ�EX�eI1A#��J��"~ȝ�X�s��6��?����l-�T�� �| �p��I-�o[cҥ�i��Y�E�V��4�޿�{22�R��f�\-�E���@;��U����ǥ����b��jk� ���*Nfh�>�})����b�L.�	0�M�χ\+�<I�R�� �P��M���q��O,�5���ґL�7�.ѼG�w1w�RϏi_��:�r\��We��}y��ۅ�jk�ݑ]��
�nN��iAh��/�@Ǝ���6 ly�ǜ��D�}�d�܏�*��ri�ҹ�-(:���*-��燉���7������6v��\z�N�4!3!���\�U�&c͙�R��,�Ew#[e��8�9[�teB��\��O�%���k�Uz��ske��d����g�\Ş|cl�D��Y)&��X�����?	�c-i���}m$�=�
J�r�L�,�6K(�����!s�ُG_-��Ȟ�x�&��	_�42y
|���8�'D��iי�Q]�6O��bA��N٢����-&��ي�(�y�����ɝ/:j2�j������_���d�l.e�F�����w
1Ӛ��� �^>c~�l��6���~Ga�j:�������@NITb�k�U�+UlҞ�~=�D�c�c�|Pg�6�n��հж������$�M��K����ԟĆ1/e�����+��$zg�~�b)yO^<�������!Ad��yoq�ݚ��l��'#ٳ��hsb5Z<�W�����XUaVʱ��z�ܹ�/�.L�N�S�2dG�qcrd��T��0tU�61����`�b�;�z�DECh�+���d����
���(�$�㑥&`軙N�l�,H���Ք��p
oܩT;  Ƌ���٧�ғ�y��~$��D�i��	�R����@naք�b��G��4�j@Es0.�J�mn�
���G���.��^�P0���p+����V9�g��O��o��	RT � ��6�\p�<xy�w�q��gA�7"��y�n:�=���)u��|��Ƃ��+�.!�]f�@꧸��L1Vi���s�I��!�#��ksҨ:�����,<�(/�tWt�h���<�~(Q]��ݓ�T�6ˤ�0��GFך%z�yI*�-,2ZV暮�ƙM���ߞ��ؑ4ǯ�ʥ!*2m��X��/�g.ᷔyb�zk&��|t��r���<>GZ��J&�����NG��(������%�Rli��߽���[�T�r���O�~a)\O��g�pÎ0�qw=CiU��,�ER�iw��ߴ�
�!?һ���y�P�~T�m(S��*�aBF�՟0@�����1��N��=դ���||(x,�ħ�]q�3$	EX⁸���SF*[�	���:c��k�2���U���p���1`���G���ڕ�~1X������<��C�(�퍵��R/_0C'�uX!����:�.���~7�LTcIk��@v�TF�o6���N"�n��Թ���Hۦo��Ah�J6�|��>�l,���B�g�J�Mn&�ȵ<:!@g��B�S`w������/���jL�M����󴼁���GPRucS`���AH�ύY�z�>tT͒I(�mE����x�{W��W�˕=571۔­��Ɵv��n~�$�i3�L��D�D��N����~���0�`dw�B��q����C�1Fy���fu�bI���EdfGә�>Q18i_D��<�����	~�#�|�� 
��>��j�^�$�A8�F81�C�R�������I�}�y��K�%^�K�V�x㷈+�jJ����&�	��ȱq���w)��D\����]/��Sk��T�81kb��3�l�i���?�Cr9˘բ�L2�b+NWʀ0�e�:~��
��V2B���W;W1�����D�L��Fܾ3X�~A�V�<P-�Jv���9p[L�J��h#i�R�B�z����	�H��s�|���N����o@}�J4�}�:���Y5(��%�a��2�o1{"q���ѷ����>���d�I�'
�!f N�`|i�t�_��'� ���
4��t���#���c:̜ZG>�͆�.r��$C��!�Zgg�q�\AdqL�']N�`�[���
vz��,�5��j]D�]R�,	�f�����d-6{]��8̨�5�߸X
e�A Y�nd��2���*~����eV���m�(՛�u�$�TxK"����*�� s�9=�`[�5��{ծz]$�j�E'Ü��t���Pհ�-�[�n����&$]qg��]^O\  ]��:�LK����h�8t��7�m�PJ����FK^���}�Kp0�H��2f��>
p8�����%�	OԆy�Ё72��eϫ�\׭��;������_��'���?���H�kb]N�S۝3�Z9z�l�ŉ����RXy��Q�Of4~�av$�@������Ql3O�>ծ�h�}A�a�b.��T^��pID�sА�Ħ%��*�$7I�x�Ӫ�i��g ��;ɗq�^Q������,���8�y���n�e�Y�p;�tUYp��uyCG�y�qK�(�N~o��%9H�$՘���s�Њs6���̣8ԧ�*�����vɸ�+�&1��/Gջdjy��C��8^�3qsd��F���Υ
u��f&�[��2��m)�}�O20�v�ǙN'��q�#'(JX;�a� �o�7i��js����J[�&��0��D���sڞ ��r��Jl'�0���I���	o��6��|3���~�T�.o��y���F|��W��'�]��z�M_>x��g�V�[-�����)��߀��I� c�4�K�wA#.��P���˄�4�#��w�R��n<�? =ֻ�ٍY�ļn�ѳ�g�qi���B2�o���p����ɔ۽�)�mւ��W9���;FS�$܄�T������kq�ȏJ	���88�:�?Q�R��/�V7l�(>w�E���Zԕ��]~*�n��ymPK�\A����G>�������
�h��uis�VK8�n����-��WO&)^PK���X�|���������'�ǽ#�?�KI|t���3�ۂ�Z���N���]O��dK(���P�Br@ 4<�� W�{�v�3�i�LcL�Y=�S��+��M�ouX��}t>��A��sVw^c�)�l�Nnw�,��!��[r����)z�>��~:�=k�J�n9Z�-g0�6����Z��]���S���s.��mʑ���g	���CX�d19_O��.%PL+)�ۻl��e�����qCFĨ��g��/f�E3a����2"�?2�;3�}^�>�=]V�K1�xH�Øݢ���m��p��N"��C�E��;>lF:�)6��'�'�i�-у�o��]��Y��j�쒄�\K���
Z���� �F�aG(�2�%�o5�>�NhYg�@�趩0ZMhN�{.��h�fa�=��Pk&(I<_�K�ھ\��A�:�6��&R���|���� v@�$j������"���J�᭒�ZI,��eE],7��)%܋�7Ϥ�[i��
 ��GDN��9(����OR�� ��v���),T����`ۮQV�>s���G[o"?`!�����c\,��� %�ӝ5�%y�^�A��D�85n�x���H��|7�2n5��e�&��*��U�@�d��6�UiR��?'����~T�#|v�\�;s� �X�>�6��N%Bg�|f�������,pU���FVd�B�ë�cC��#h�p�DiB^�uLxf"�z���%�!	��6�^���{��ZJ!�<9k� 1�10�n�h�m�Q/i������P�F��ѳ�ѫzF����i�	�Xx��G�]s@�u�S��S��(�2�HM�ul�4�_�`���v��&�k�P雏hX���#X�fD�`�߱�sC6�v8�u>v��!�b �Arz�4��V9kb!We�^9,�~�[���&E��2*���'����|ؿ�1!�jB��{!sM�|��5ev��B���'�c�$�&��GãP�R/�+�S5N��-��T1P4j��f�I�����_-�-�[�q�vk|V8^]Ǥ��/�QE�Dާ��"4u]�`	��WqF04����윮w,����k�������,��E_��:�<�r,�df���@�����`�$ۯ^K��PwM�4[��yq�Z�C��J ��0O��Z���v�}�5���d�<������	���-�	���E{V5��~Y �t�l�F�y�Bd)~��$�D��َZ� �?����1� �l�*7O���v����!	&oZGk��Ҩ��=	ǖ$�Ie����TI{e#�����#�3ӱ��O�p�VP�^��������q�<n�����vN�l|t���߄����9.n��L�(�y�e�Q�/�y��,[O�lר}S����	�=�|�&(ݠ�)�8��B>��U˙��n��[�(��"j<N���y���Ķ櫇�E8-7a���u���v&N�&\@&R�V� �w�6�y�����I���?bB�y �P:����V�mX(&X�G��<��8Y��^��e����E4 ��V�؀���&ܙz����d�DP)�TcH�E�:��t������}'��VQ�w �昇bgߛm��-��܉,%��%�KN��G�r�.���A�Wpُ���Ӌ�����y���hC!%�(C6����5��l���
�`R��O�0���u�:�tm�q��Q\�oؙ���B�#%�ۡv�yBT��0vĨJ�eY��#��8�M���L��[h�6�J��oy��a.U����=�7�#l^o�#���X)j����q����"�F�r~[Ab�_	��!9�'�4"W�nKQ�'bA@�h�0���i��S��k�̪0���,.ɺ?�.b��kWƃ���&j�]7�i��d<z; ��;��s�(���� �E�J�J��w��(.IN|�mְ���Y����	$�NpČ)5��׈���O<�*�%�F/�������1�8������tl%��J����������)S��q��{�"�!�6zS��lX��+��8���$ۤh �D��O����Tл�t��`S�ع�'h���Bs�t ���d��	;!q���,���b9TN�ˋ��3�ݨ�/#�W���/O�#���9,��F�P�!���h���|V�|��+K�B���*~�Plz�9
e;�B*]����J��D���s��,ņ�naJ��:R��Ef'غ�`��4O�"�x��d�����c��y-<<�[ʬ���<�^������X3��',�~�D�a)���<�Ȑ���43Gq�S�;Y��/Q���_�c��־�zyd�w\Sgca-!�n�D��Qvڦ=^�YX�q�Fْ<h��+��#@�q
TU N����h�����ȓ1���Q�P�������v���`	�Wog�&�fj�6����&@����� t"����#��W%l�7zo꿹�I5>�y�VxPQU� ' �3��\�>�� w>�k������;K �� &W�|�4ѿׁ웗R,��3��D��XE���Ҏ<��J�9=h6{���w0����$�E�4Ժ����@�taҤ�lE�h,By\����%×qMW9B�=��
sxhx22Z
T1zr�?F% �/��p���Ѕ��+,d�v" ���br$�������>�0�f'���$$�d�� V��λcEZ`��Q�~$�v%&�a�'��f�'�p�"C*|Gz4GqlN}N̓���_M�HM�=��z�)��,���@.J�;�%9M��`��D���$?����������F��+�7Bv����V�Ne4Kg�>=���]KC�T�O�p���Љ�D�VZ?N��e�>��3#�j����ǵQ��r�2�Y�OM͜��[���H��>#&�-�l�1��L��EXRCs������ �C����U2�$@!#�Zk�k���h|6�1/�dE�f���7,�ŋ�eN�'όM�]�uDM?���.�_v0#[n����[��!g5��$>�YrP�=,�ֲI�����#Da����Ro,@s��C���č5�sP(��{����c�K�����O���h���S������uN@;Y��
K�����D��o�����@o�cd��7����<$�G�Yx{i�j ���%�өYHp��Q�q�﹣4Q��z������n��T�D�3���OU��$6�}�h�-ѭ/���y_mA:�@9Z�v��n�}�=�ǂ&*QxTCnp"j��[Λ��B�
Yb�ԕ��X�L����6�BA����W���� =
w�A��jg��o�
}�rl������2��H`�M\�&^�䇻�֩ U㇁��1��6QȌ��J��!��&���%÷�G���J��T�&���,���\Gē��E�6Ke{�v�{����:����Ӻ!�t�F����^�1�G�>�[Ԧ�H�+Dk)z�B�p(�NA=·��
���H���A���{g5��y�q��m2MVZ�K��qkG�=b��D쨮i�Z��L���$���
<�vE����Ԏ+����#�V��q$0�ҭe5�����V��zf|2�Ou�t�8\k�F;Ƴ�A��ӨL�_z7�rO_���uGc�����"���Y��Z�������m�?*g�hS��SM�P�9x(�꜊ܗG�.7/q&ҝ��z@  lNm�{�i]�?�*v�Vj֑�0�l݀��.^J����+��*u1��;M����~n&<�!n�:�����܉�9�X5ݱ#�9�1���ȸC Iq�?�b�)M}���jd#�ǾH,zNHM;���,qA�:|�4J:�ےʧtjTy�TH<�,�zʍG7�-r꪿��[��:s;�$k�Aʰ��LU*<���vm"�7㺎���Z���?��Q&���\����2m���0��tT) rJ}�>5q݁����+���ׇ��d
�i�q`Fe��@�)	C�m��G��}ͪ(��H��<�U*Y�Y�	��~�'�H��%��cl�{A�H�m�d|m�'��>i�� ����D'�rj~{9��i��U]]N���nC��aj�(H�e��d�L�\���M~�Y� �Xa�E)ʐ��B��"C���6?������zF����'�i�Ƙ-nr�+x�����,ߍq{��g��8t�90�C}��F~�R���*h�~B�:��K�8;R��{*�ͧ�D�+�u��E���XqpbxqièY=���v����g�}�֍:}Je�$�X�gٽca�2M��D���\[F_��4SX6�0l�"���,'���{�h�-Le1��9U�Q�;� ������-�5]@�)Ȏ��/L�H�8�>�o)A�g�5iO5�.5r���	i�PH��DV-W�b NM���{�[*W򙛀jOlf�����;�D�Q)�H��4A�Y�hι�L�<'���Y�ҍ��#���ٲ�c2�J��<���h����b�ʁI�>����@3{�OH��K#p���,��ݰ4�)�:1�ԇ��l�'ɾG���ћ��6����o;����ۗ�me�R��<jHh^�v� �u)�ߑ(~��z�shOa�h������O6�T����>U�6s"|������vG�D��"�L:� ��Ǽ�Z���X�Jߊ�o��/�=P��v"j��an���]����]9����Mg� ҕ|������b�,���+�G5���]��-���\�^�r��a�l��+�I�6tV���?
��9���S��Ώ�z���:��t�㝹=�d��?џY��������(��e'V�p��q���_j}��@6�C�sōZ �Ǵq�����k�&aN磤��f�V��	@�?^<�1�i\9F�:
o��3IM��A���`|�	e�:��x��x��HѨ�P���7��cO�����zh���BV�؆��,��q�,�H͖ Fu��r*
�<��j)�1v���QV?0�Y9�� ?��{H��<� sF��)($bB;��;llGH,b#*�v:�?�|��4@?Y�������#�7ml��&!"��U��gp�,O6��sjJ|����l�E��ז=�.tY��݆�ɖ�Lcil��2�
�uӖ��G/�~K�Me��~շ��cA�>������M�!���\Bi��$� ���|��I����WaYF�AZF�S�7	�Dl�Bqa���}ْ�J�����(�U��XΣ!?����+x)p�9��3��;���h�Hv��7�j�Zo *�C���M���b�ܥ�K>��=A,Cӡ�t2��[����i1+ �6� �F�
��N�s3X�Q����r4BUl���kt��+�@�q/�� ��4�X|t�s�$��D^qB�m��ovˇ?	����.��e���ڤ�3WVd��D�+�q�w�B�q�t�e�f�
l"٦��	���l�D���w.dVe��r�z�4���~4�7nnrʻ��WJ?���v6�c�=�-,�X���p�q�{�tcE|_���9��>�W/�I;�t��肍Xh<��ŗ[΋'߉��iD�~J�X@�Wz� �2���]#@��L�
�b*7�b9���L���`�C&���gڳ��_�������zqusT]��vYN1Ö{��a��0q�+slHw�0P�K���F��0��q}Ve�Ϝi=�su��d2����^�q�|�
��f��ǘ��C�^���}BK�`h�j�nJq�$"�RԐ�b��l��þ�%����Մ��z�l
>��P�2�-��s���8h��	�D!���iw���=^h!��\�!��5� N�ɄƊ�˙z���pK1���[��u�� ��G�T&�%Tt�5���ȴ�PЈ;/|�i@�^����ć�Ԉ�_�C%ZQN��*�H;����x=O�RdxQ�V^B����'A�%uU�u��~DDl1�������
�f�"]Z�����&� F�j�U����W)k���]��̆�q���f{������pDhXA�&Dԯ����[��~���h�_>\4>���є��4��9������dyO"�����*���]'#G
6%�S8��߇�!l���9�T#S����ɺZ[��bD�-�㺎�m��������z3mF[��U~h_��_k�q�u����ш{�W��םd����r����q���ZJ��dWe5��%&�9XuׇK�+��E�T���b-=q;0.�,jn��~�-�' �-U741�4�.�.�]k�'o�� �wU�`��uL��7� �)yH�g��$��d,iq+*<�௧1n\Z��CM�w��toG�����)N��Z�(�Q4Y��0���:/Qe���ŕ���C&����t
D�\$�)U���.�y���U�����oڳe�Ҝ�P� jn�J@TE|7]K�Tժ�ړ�nO�Y��R'��۝�v�R�N���)R�z�)�rQ��-����]¤��4����,1�����zq��a��Ž\7�����De�*N=i��|L���]�F#�H* ���8���M���9]��g�2v����~���r�"�_���]���E�i�G�]Z��m��ڄd��o;�cނ������b��n����K�Z<���Ӏ3s������_�5&Νz�ƙX��8�\��uZ��k]!J��#�*�ov�.����ОT�:�u���`t_{�P�n�̟���6x�~��<���U��J�F�w�r/��'D#����	z��ȰA2l-W���XKd���w���l~���9v/�!�O<cA���N�O��{��fo�v��`�|���o��U�� Y>�}g=q�O�F�&5��]��Vg)�ChS�/�����817��$� ���o��w�X��|��=���l���_:P�<2p��/�ap|c�D�w��:N�!z�a��8�>�5'�˿5fr҆�}�)�W츌�4DX&�1���{)��ŘcH=:2`o�(MF��V�?g��p�fl�u1���N,�J�Я9�iM���"�����r�U�d-�Z�鰓i�(	t��47*��6�ai�+r���9l0B�*h�-�'W{�%��b=*��B��	Sq�H���Ƥ�|��0$I%�ډWGD�ĩ�X[�0	ls`�l��l�ƃ�yu�76\P��v�{����g)��-�̀��#�t,�.�� ��d� �o(���v��U��![}�X/`�gJܦ���{8nya���f�r��Ab�)��pI<�D bd�Ֆ}���~��ۡap��L����H���i���L8��<
wC�?�B�B��rr��U�'���נ��o,m��NXB��䪇�1݃�WC���V�A�Ӂ���������:nϙp�-&���Q>�t��	�X#��\q��8y
e7 t^���Ew����d�/�k�~�����@�ܧC����Dљ���h�Q���Z�#��U$J3�T�)Vf�&���j�q�R�������s�&A���ȑL=&U�����f�.�Vy�9K��t$��18���CU�F`���m̺�[_حK�
���4z2��L���	��қ��$E�	��U6�x*
W�x_7W�ƽ.�*���v<뗞CzPʻ�K�)��2�ġ�3��dY�����P��MY��L�x��8�$rH������y�wգvDR9�C9��������*�����U��B�VEp�mChw䕔�A��؜��o�p�Ļu�>ѩV"šI~�$���>�m���)NV�9��Dj���Aª���Է]��幘�_��[�h�֝e�
(�����Jb�r<"��Mһk��A��~\��q��\D�L��6�܏�%d�����v�/��睦�8��&�&��;Z�L�
$vu0�i�l���2Bu�mw����q�G`Ue�܇�7T@�;P�7؀���[�`���q��`@��Ⲃ�rd6��l�k�dZS�װl>Dn4��Y�����n����d��&_���>�|L�a7%������}Y'�V����t��rۗ
C����͘�m���uL���+���M�y�9E+Š��A�p��L�``H֍T��c`p%clGF����	c~2>q�������к<�a�o��1Eg��J�z��I��]|�8�N��WX�4AS���<o�~��hv��e�]�#�q�_��2�2$�/U�_ Xx����8��LJKϺ�N�%�1D�cU��0��t�0���[��Z���BQ���W�v��:pP���h�x����� t�����4�4���(��A:0�}eL>X~�g;A����ؖަ�f:Z�]MM	�B�}����&�J�iyf�s|!�|"۔�]�JqI��|�[�,�k	
t���d������~�O�~��ݮ*����]�H�� �G������u/Iȇ���������2ʐm����֭Z��D���jȌ��v��U�{f$�����k�
y��xYo��Lv>�fޢ��=�������"p�f�ݺ���(��b��K蠉���2�r��(�g��	/�62��%��e��Po09v��-)��YT7�!t��M6�7�O��Q��)]����� �9?޸ �/B��p��Y��W��b�w��$�����)��J�qU+��@��z���?; .��қ�"��!�O�G�=��~Z�o�H��Ĳ�,��o4Hc�)�υ3|,8�X��:�a���4v*o� q�����"ͷ�@�`d4t����D�K�-���:\��E������»���g��H��pZOcx����ŊV)^[DXC�뷕�&�s�Ǖ���R1iLC(����23��G��2��ӟ=6��?�"���k��}X�"C��!ퟔ(QR�x�F�(��i��JDP}���J��.N>c8���J��hw27R�e<$m���8��S����`!zj��D[�=Z$ihy�d݊�$�>��]9�X�;�Rʿ�5�%D�I�� (�N���x�r�"�+P��;Z5McZ.z����8DN�
ɉj���4=�_��6`6V
��%�hdA�wO���e����Y�q����]!�R�,���|�M�HpQw��Z?�$�-��Hȹ5��*/�R@%{�4�Q��D�Z�Ħ?���q��yrI����?�����+ó�zTY������%��g��0lFϻ���s�!��>��W)��edЕ�!6�WvTǇK���z����lI�m:��ư��+ۜ�Q�k� ͎�v��vŴ�Ȍ/�EU��x�*/c
�'�S+��Z�y_nuf`Y#F�#��Mds�oz/ȠU?�B��A]{P�Y>�2�x�̬��w�;�)7�9����;h�#T�~����+xl��9ݚfI+yҾ���͘���q�KR���8,$��#�?}���KK�R`��s}��GL���sF��%蘛�,L�i'�|��"ܐ���@lHc��q�I&���t����T�3���W�a '��l��D��U���!!Y(���X��BIL������n�h�[V3�t�.wRm�i�KR��Ad'����O��������/���؞;=U�\-�KK�|V��N�/��W���W:�v�*T���,*�l���b�4J �!���{�R,ͦٴ�ӗl���x�G�v�n�������,��Ԣ/�!9�A�u�q,�`i/!�����+�Be�h���a��\8�IZ	uh��\��:����ڳLl ��sr݉��Į���-r�U8��[�C�dI.S3��S�S#N\�y��K����$�s{	o�Y��:Lũ��\�ߕȉ�#X�7?��Pڵjy�*���{h#�_����ZZM���k������n�L3��N�OJw �����Њ�;;U��)1+�3 z���:�(�4Z�.��@���Fs�Y�����p"�~�}�w �����t�O/���hq�ϥt���Xr4����Y�)�395~l>���4���<��g���@��XUfb��NOq�c�$�R�e@�P�ڪ�H�hBF_�4��a�⦍a��O�d�D�8*1vBFԐ�
�l39��<��ƥ�����(a��Q��;I ydH�&&a�b}I������������.{hGW�[����+����!��%Kj֌:�˧�Yd s�K�@a�H���9��M��cfZ�(���g����M��&ت�T���s�[2�MƸ\*b;�T;}b��>��a[��5@C��#�%�R+.�:��>���V%��.�I��k���12���	BZ���\f朚����tT9��v+3��2�d8��Ŭ"6"��������)bov$�ۀ�bb6VNv[�@<t��]��H���'Ip���?w�T�S*�ɮc��������$P�:_&�Ͽ�Q5�Q�����/S�P3���\hꁫ�\��]�gK_�IZ��%gw&uX���p�
x�����+��t���/X���l�`H�Z��Vp0HQ�K�T������"���8w�~a|0��Dg���e�w�b��*�<�M���5	�٬�Q$�"��{de�.�����V{,���sw��[
�v�e��;C��~�����lyX���++AΗ}��'��;��jc>U� �}U�@�N�_���Af��א�g��򔋊O@]��c?�	m��bM���j��r�p��b�&��9��1���H|�ą�
���}4$Ӏ�GB�x�@H�$�I��YĴX����E���'Z��Q���t�㸌����#և���0e�U��0�H�N���'��O��X����m�]�9w����<t�c����֥�fL�^�������������P5M�����x��5.ۡ:g*��X�4�y��d"ڪ����ꌼg��o�Zc5"Q�l��0l�� w�	���ӄ.���|�����|���A�e�ȴ��HP'��W�f`.��Q�M?�ϊ��R�O��k��9yEr�a A���e�6@���`Ϗ��0��;bJ���Lؾvc��(?f�<|�7�"�_��Ȋ�|f��������&&�=L%�u�{��h�)��I���c�/E�&g?��#Q�G\���ː��s�n��Db{�^�+��q�,�؇G|�H��ﰱ=O��Z�\�+�"9֒�+�M~�o������ӕ�D��Fb�(w?u�ߕ��V��#�5�3UbB@?�����pT���<5���C*<%�� ���چ���3�J�EѼ�̲�a9����z���M�R�%
��w3�P-����*q-MZ����ƞZ�MmU w�W�:�(�(f7����)�+EdtwO��{m�	�0�l�b���y'����n��qrj�0�wtKpHWoT�E[K$Ia�P���������;��85�i���^���I� ms��
T�V��Y���p$�Q�H�,4��Y6Kvh��n���hq���A�������F+EE�f�13�AKti�j�D<t���w�g��
�%_8'��A��g4�}%cP�������y�v��5���p�p���(��Y*_��my����a��mK���@���;�����0$&\����	��&2�f.�/���x�S�E����J������"SQ~��T�@�B���h�S�'H���O�W����V�&�֤��S�F��9�������8�۾ç?GWZ�؎}�0w\O�~_"����Z�x۸1�>�K+n��� �Mf�"!�Ϛ1���I ���������r�$�0k.���	
q�h��d	���&\��>�����~ ��E�g9���c�M;)��$a)�C��B�}��/���EH��.�M���E'�Ĝ/y��a��۲�#\�
%���$4{:���R&�,<���c�wN:�P�u����b�����l���C�ުW�O� O[��U� /]���|�'Q������`�Bq��^���#6�V4qU�0y]V�����M^��a������Z��
��ϛ�	��
�N:w���|��d��?gW�)����L8�FB�w=���7��ǘchkޅ�U=�K����Js��j�gH���3�NN�..V#��r�q>du��}i�|���G._X6�;�El��s��3{w�/�!��+7y� ².V���p��>����"���&��T-��^X���7�� �^G>���K�Yn¢�vFA�A�F�7�G"N�mܿӟ�נ�0O��z����H��6q�c�p���e��|��1]d�/L¾
~�z���7-DTȳ�ױ����h��ʞ��JV��t�l�8�7�&b%���<q�����,�гv����8F�����E�F-+����Ak6��m���@�	�D?Z�z��}]��KB���DEo����Κ�Rr~��)B�c�̫tS�^"mPK߄h�,��V�|ylf�Y�9Q	4_�<6���x��׿�_o �
�ye���q�.��=cW�LH��cqW��V��|L��.d,§w^�L�.�ק2�������u��Gjo� �y9]ŉ�� 1���@�L� (��T�����;Å�Pb�nY�Oܺ*�uAB��|_r�^<�Sۄh�ȎFy�}������H�M7��k�T*��0{|ᐕ�~�Wji¢�Fl��~��}��V��[�!x:܊�_h�Ċwqsm�ٌ�p���C1�M����q�H*�����?����� �p1�����7"�c7[�O���P�"m�t!V3�}�H���.������D��n��k۟渕!�Y(6GH9k�otP>ӳVܹ�ʷ4�Y���0��*��`�QQ�I����`��@*,�����UE�fjǘth{�?�jS�q���my�3�-��IZv>;MK7e���tP+�p���~Y�s��M.�1�rF� ]@��&.b^­0��R@aE�	�9�*���XG�2�ÝƋ*��wju"��⿶14NH N�{V�^L�&���ӏ�jG�Ǡ�x"oͣ1�0.�-��k�&���),4:��jQ�e�i�� 4M�Zin����G�ٖ7	Q���v�bl(X�����%����#�؅{&HH6��u�6G)��Es�Z���X_��˵{By��=�5Q�Z=,j��y4Ǐ�P�ep�Pb]�����Ͳ�,���b&p�)�`���-���c��ަX�l�V&�s�C��ʡ��o$���R7�s�#��$��7�ٚ�,����[�s:���&����Y�d�|_b��`e ��F���b-��7G��/�~�n�)�)��y��M�>h�r/�c1��R��@p����P��䣈��	�1�>k�D
�F��˱��M�4�`6�ߵ�T���ŗRʝB��Y;ͭ������/��A�{MoQ���S)�PK�ș����)������>r����P4���:���z�=b;;u-��=�vD�h��.Cp�����H�ZQPd�̘�Ӯ��ҐeW���I©��,sN�ㅾ�~YvX1���l]M��e���J@�O��Ʊ[ O"�Eq�Sk�\l۶��4�x5�K��C�e�~b���[�^4��xv�k�{c�~�F�ґ��-�'F�x�����fht�#.d?zx'�=�痑����"��P#>�p�x��М��
� ��������;''��vU�t�m"����+7��q�����ƛ�����`�k�ͣM�Ow�Ȑ; ������Ӥ�\��;љ���4�B,�@�l��8�2��w`����G���a|���y�=̉Q��Z��Ma��Pv�e��?3Fs���9�wx�b�K���Ы#�wQ���XU{�z�Ч�8�$�ͽ6����y)�Ž�tl��
>�~�I�:A6����G��:�oɒ��:J{�YM�p.��ڽ�#�����Y���,����2�[�����=&���=�Υkx�9^E�ς����r�k]�'�H���S�T�7��cڀ�����l������_���U�/* l`�<�����U�q�-/Y6;X[��� 
L��8y7���wV�_�]G:����ї����� C?�4���$R��	�ؼɶ�ה�2oVҋC�_e+6�R�+@ͽ�`��Sf0f��dS������W�n�|vdZ�����@h�_h���ta����@�#9�/�+Ɲ^n�H~B)% }� D�v��zB���@���lff�y�7e�6���7�p�@�w<_��F�I�(���<0�����s�L��-�i���!�t#w��+�r�JQˏ�j#S��O'�$���}B;�'x}ߓ{���4Tq�o ഡ��>y��l�:��#���
B�},y6�gD'i���o��x9Mb Ff�	�i�NL�3�g@�g:�����`r�� f_L1��_���|0�oW�Cˌ쟱�^��Z+XթaZ����y��|</�Y��Pӥ�
��|̉�q�0�
;��X%�L�q��f<���	p�+A#[Ftm�k���{vfv:]�Q�̠ϡ$O�z�HO�ːK��މ�F�w��;+�*����>�����L���Ac!��̲7�j�Y'�u�{����`A�d���N�D�QA|e��#��r���?gba�jH��-�A���CMd]j^�5���©��(s��vo�D�E��KX?S���<K���(rUz��"�:$��}P /��VU
��Q�w@:�BN�nec��|?o�%%�=�������%���Y
pԷ��9�_/���?+�^S�4�gh(\/	���M�\}!|Q	2~H��N��]� Pe���|��n��F�d���<gom\�`s���{`	֞��܀��ϾSd[+�ur�S�+rIz��3D�ʙM��Ns�Vۈ�1�8 ���1�TCiqS�I�3?]5�b�l#�]и�&�(�l�Z ��3��ݤwϦ� 	Zk����z����`��ശKb51tH$��aZ*�3�E������g[0�������d��:/s^=���w��'�#�2��m�>D6�����t-Ot�W[���o���m\C~���cz���u�8���4���?"��1����cUu6�%��\#���D��xK�$���owL@��ih];P�p�,��95b��;0���)��(�Q�f�u\s𔷮i�f�&����'�>��8U��s�Kc��"�7�{���R<�#h��+D�kCs������,��>/��W_ft��6�:Ջ�X�H��{�c�Iꔉ� ���{䬅�}EhZ�J���7�K�~w��f<E=?Ǘ��I�O@u���jXcO�%G:	�[��f%l���V�V�/��L9��h��K�
~���_�t�]�_K|u��6
�
�S����h�C�_�ڙ1��N�7�q͵����^��p*�(Y��}v&��"S���d�.]�8�w ɦy��a��,T�Um ����  Bڇ����!鼋�8s��QM?R�o�oh)5N�*���������)[��qo�[�������x��GY	TB螰���� �?BM�pϵO��'�����-yÒ[�C9��!�H��V�D�~dg����z�+�c^\�B%|��r/e9[��*Dа���?�#Yz��t�U�P��7�<Z�'<��|	OO0��@���*�'��i/	���:[v��.�5��B��X�/��hN[1�߻I�1�s�a�5Zwx��J��M i˥�1	�Ӆ��!W[���3�G�V�v��M�`\�׆��^k�ȁ֣���P!��!叛�׋`�j6$��1<�|�!���wO	�j/r��o5�F�L^����Ck��FF���4�Om���g=��>#ՙ.
~���(�I?3���3J��n3A�����c��!(䞓tD_��9n���c����ɝ7�_��0��-�+���{+�A짦����[ ����#r��G&�ԝ)va�C�T";Ad2p��I��Q��b��� YL_�C�UԀ`�
k�T�%ؔ�w���1CI0�L�9��8�[�WwU\����-�\C�Մ���,�U��e�|3���)/���G�E��+w�Sc�|V%����h���1Y�@:DUB,�.��^�%���|*�Ҫsun�*0��c�q��g����L�D���o�ܰm'�0��sn�5�kI��;����SI�(�.s��6^���%N��"T����H㦞�e��]?�'�j�r$1�'%\!D�{�Q�;���v��}��Ќ�Gܵ:�j�:�uP�<����S�2Gڧ�Cf(w���t�"��T�/�,�o�����O����&l
�Y�ӯB��&rK��)ḃ�P�Ju��Q߄�pN!�����T٢�L-b@F��*H5d9��f�b���^����zx���Ǌ;SR�{)e@��>����U{�XL,�\���2)�E��� B�k�ٕ����;:�Z/@��}�J�L������ ��Y�?tP��2 Ѧ���O�-�ՀO�}�YP�p�\��a����N��jB�����ou��]��&%�E��w���~�U�.�fG�;�_g5CF`^8�FT�8ť���p�m�'٭���7��UI0G����XV��*HI);i�=mO��o����WsHT��"��Ⱔ�4�T8T���˵�Ӱ4���D�]��d�x��L��9��)FU�9K�t�)!7�uDk�S��0���+"	�R���q�в�!�V������f��2���k���˕������\���!}�i�����}�y��.S�	��,W�.���b=$E�s@���:#V�am�q��&S�.J�=]Y�	"�zV��ړV\���W�Q�o�yP  ��؂�(����I���\���"�.�>L�eFo�'f�l5�,�}���๽��eS{6-���L���~�C�3We`�7�3q[	�d�Z��7;�:K��S��*xn=�c�E��xqɿ(l���鐯��H1��������A ���ٷ(�Z�R������˕(��&��a���{�wB�,�� ��F�� �0�a,���~ѻN�Hu4��о>���R��(��Æ��ɰ3o���0�q۞E�!2yw5v�PC�{��jP�k9�p�CV.V���N���"����~km��Is�sL�}ɴ�-|)�0�g��5��Cw���#�E��֟� Y��)���mOns^��\�4�F������%xĿ

Xu�;N~� �`��F�@��\n5z�H@���[�jE��[P<j��ټ�y �r�3%�/���S�g�t���=6^���X3�����T8E��臭	�u����#�J� �����<X3�[%��jc���Cl���c�!���O`6���X?~&�[�}�-;n�eu@ń�]W���Am���m���]�)�"OZ��������-��5/'K5R�}�t�~m�T������O8;'�N[ԙ��%n}��Y��Ao}>�X#��DE��n5o	�8<�i��ַm/`�s3E1e�p1�Y�FM:�{�_̃IJ����Q�/OW�I��'X����3�	������i���s���^�T'���������6���,���!Q���m�ؤ��/5�μ�״�E����\Jh[���|���I�9��t�y���$�P�J�?1�n���t%�(/���uG�0�Ac�!j��$�ͨ&�+���Z�A���<I�X�j�5r�er����2g0����a�Mve�>09�P������<��S�@
��צ�l �*���Z�qYbTA^DR�0�鳁�9L�gr�D����c��o�2�����I;U@�/�k_��M�i���>�Xs���l}>��y����U���^	�7��7�2�9��$b�I�7![!�T��LxU�����>T�'�Ȁ�`��l���zK|��������-.B-T�)j��8�w��/��C�9��:��KEϱ����FF��d��G���$�_a#cͶ��B��J�d�F���J���)U�B1�TE�e�pS�V8�#5��.8Ky��rU%��ǯ!1`�����M4a��
n�Tp�ð�M�Мw����&W$��<���N,�C'#�=(2����k�!k>o&�W��眿v4Tn�r-p��=R��$n���$�{{jWc泦�O z>������~�p_���t� �?��
��H�ӱ�\i�������RL�E������8"�+7�a��n}L8�@x�����>B�ʷ	%��a9�*���ϻ�I���1��I�"��;jU4��W��k���{,���~W`M��a[��#sc���^JB�C%g�ˉ>w��d�ϴ�-@�B��K�;_�c��!|M�0��jWCɬ���y@P��R���cd%��řL�Ѡ��>���5����+�nv�
�?�uO&����@��"�C�*��܅���F���eIgk঑���.}F�`������vy�v���푐H�$v=���Ah?�a�,��V�g��_xg��6�P/%�>��],��i:1�����f�E��QX6��t��Q������3pE�k0�Ğ���n W�L�����ձR�(1��*P#��ęA`�����b��l1T���MT�z@�T1T�|�vjvw(<�@X�-m��@^B��A����6kƪ2���5�R��H-L�X����}�^[ĵ����?B�GPU.��]����W���S��A[�JJȤ7Uŧ+N���E�t�>D�b�O�;�Z�e|D���߉��q�>����D@W�r0��p"��/FO��P�P`/�=�|FHpJ�$����!��O8AW坠9J�4�����J���`�6�ݽL
�`3hn�97[0L):rC\zv:�\ǥ\o�+xq	�ά_��[�ｬ#5T�׭��b`�Č�I���8�'�R	�;0���W�r_wn��^��"�	�ۋ��a��Ͱ�yQ]A�:g!:��ޙ����D��߯�*���t���=,f 0yn�D�i+i%�V^ge{U�!���@[��VJ9?۸����R<�?����C��������QMM�����v&��1��`D-����
�Gi���CG��+���m�ӣ9p�\�'y�O���WΡ�2�Z�h�	�����%1���Z}�Zd��r�C�=R�k	5]�b�� �h��K�����������=HE�U�%T�XۤvE y���bN��O�Xe`i���p�|����-�����l��B����#i��� ?��`�3��S��⻩�ʺj[�yy�,w#T��fe/���{����?5i�6Wx,�+���^�+�:�/��T��K��crZ#����(q3�"��H�;W'�/}���j	߿��TŤxN�8�˝6�6�z�����O�`�F��I8+t���2����vL���P�u�+gUR�F�� ��2p���i�)�m\C�Cf��pԲ���X-����X�f��z�nJ��$X��At�,�0��~�v�9���o��z+U�Àщh���{ډ��u�t�-�怵��aL��ȭ�)�P_�-��������\pv�jѹҀ�N�� ��-a� WVCN9 n>��޹i��z��HD�\b������C{�u�$T8��k��'t��m���֭rY�V���{��b��w~�Oz6.¢�W[��_�ڂ������孰����5�n�X%�)����B��r��m�R����k<|�,$�\sñ��~^}�g���h�ȑ;�H�	�7M�%Y�l�I��"�`ta�:��S��4�Tv�p{���;��vw��}��F�V�����E4*Kd��1�[Ծ���'���O��lJ�����?�#tqdZ�ϊW.�F�&t`��W��l�T~!	��B��<n��:��v�oP�����/߂e"6�q�8B"Z�E"뮅�e)��+�{�R��u���o�6�S���R�ؚ}��a��	��[�/N�Y�[9]yá{vji�t�J�o@XPJD{>���V�l��S���9���ӽ��oQ}�QS�O<ϙGwPn���(D�t"��@�&;s8��qJ�%�}U�r���͚�o�
�P!.7�ې��dTt�+o�-�\Ŵ�2ŭe]QNh�b�*��M��ui3�K@5;�����I��ĳ�܋�0���J�<�W��C6�d\c��N�n����!�)�G�ŋ�	�2
��!4�@6�U�Q���S*�nS�,����Ͼ���	��	��@��ɮ�e$$H�������k���<�(ֱ=vRv�0���VW5�&>��}�hJ�\��(p���pyԱD����2�)|��K�;�;����1��1Te�h���Gc�FKg��_?���lK��M��a��`��lpI'�S����r��ͧx�}̜�@RU&��H�t�ن�-�Rp����g��U�tZ,�]�MkO�3j^����.S`�s#��Ǐc5�ʭ�X�������VY-HB��st<�z�2E��j�h���\�$��YY;ǡ3\w!;LyV^v�Q/�?ٲ�@:o�+�K1_�ـ{$D��ɸQ��"���2׀���fSF��hۅ+�+��Ή#[
p�M�w"Hr�q{��Ю�FKC�{\]}��/u_�í��+��x���/�ڷ��gS'E���%��៖$j�A�b�6MjK͇rO��A��e�;%Q���fg�^L�6��V��O7"��&i/Ǹ���@!E@���_����+�;����x#H�?>G��;���F~/E9�wB�2�COT�!g�(����	8�Y�d�\T�R��MEk�����{�E
��2$.g|�F;<�If�őz3�%�Plx׳��q��,����K��|���,d=U�i��D��PD���Y�c��d9a��P��XVh'�,�L׳��l{�q���[X�}��}<�-��g4|V���؜��^�QB$		�#����鉘P[��)3"�<B�z�$J��`���eU��T��O��{�_�2�2[k�_�a'ąN��G�`�YY$�<
$/O��Q�RR�uΌ}��#���v���.�Hbx���-x�dpcst$�#�����3+����?��ߝ�c�#|�ۅ�Q�/x�jI�Z��5e@p5|<�
{ƢRE9�5 �|��])�������s�(�lL9�	�r��q�d(�bZӁ��'ak��溠��)�@��O�.3�Dy���O����f`�t����^cB��hO �؋�$tg�%����#]��eb=GS4��%���/��Mc>��E��a�
��Qӡ��d9�Sҳ���kO��徚�D��7O�]��?{��_�X�w!�W��*��TAZ�G�)��c+�ö�	�{ꓧ=縄����ˑ�#��wo~KX� sO۬.�l{,�[�9�-�����t$uԪ�^���e��,?z$z�7���8xY��qŴ�m޷�DLh��	�HBd�`{^� -�:�����,��-i�0X��H�hÜ}B�:3n̷�&�-B���E*�Dm\$m�Q��
��Y(�FG�:��s4́A��dT��9�$s�s��۬%6�cxf��N�b-rNA��)p���5�S�yd5�;Q?�3�I�bg�܏"N|\��ޝ����G���,�`��C8�1���b�L����S�����zDu*�c�d�pi�Fɷ����������VOQ���Lq�!$��(7;w[����,hU֝ �"�� �n*
N7�y�Ȅn��$=�X��$�*�%�RȜ���Ӱn1���ߨ�������q�_�����\�,+7�Ǹ�-U��s@�"Q��[F?������e2ذ-5�V�Y�7�Y�M���������Ϋ��ņ9u�y$���j�t=u��+uZ��}��B%�6�-t-�y_RM~��H��y���{��̸���E�q���kp󍪇�$2R�^՝Ý����LC�^=��i�j�>�oQ[��]S�^
��ȰK9�J�Q�{zT?���wMT����OafN,��o�B��wAc ����GLi�|j0���eCX<�� &;}�p�3�1��Q��3�圬���Rk���q�6(�(����d��`9_����)83���쌕����|S]��X�T=2�'�]b4�m�!�\5zP k �gg�n��~����ϋ��4��<�g���X��<C��k�J��S��U(�����x��
�W�$�VÇ#�=�Ѩf~hT�����Gr�R���=U=�z��gy�ć�lÔ���J#�n��؅��7�����6m8����=c��]=���WG��5��a3-�`���r�+��kG��X��Ba�Y��s�*H�C�Ñ�7o���<?Q�:K2��]�?+�^a�n�����&��=j�w&�s�<����辁���z���U�5��Sߞ$-ei���w��}��aQW+�a�/�kI�s��jD��+ˈ"��	S41&Q���" ��\���`if�k�?/t\�s�LP�k�&�5�y���i@T�K>����b�3��z~����jX�2ﰫ�"N���q�m\�^X�V9
3��Q�lZn�����A����ebZ�5�e�6�<b���~�imi!{�z��LLI�0v$u����P�4�N@wH�2���J�}vZ��Y���Hi�@�AQ�;��(���aupĤ��F����Yn����L��,l�-p!}3�6etdn�V�B� ���}`�`��|��٣�{
ɎM�:#1Q�G_$���U^����(N������(}q�
�~�y���/8"���avǝ�+��U��(i1�(`(��HGw:��l�L;���z�������F\5NV���%���2�MI������m��\���ñ���w]o�@J3qړ�sR���NX�m���v�6r9���}Q��<T9RA���7R#Ir��C��Μ˂��&`3�KV�r���fuD`S;�C�ρ �X9%A<(���7B��CG�C��H����RGhӴ��w��,>>��G��4-���D�"����C�n�69��IV��Wu�*G-��ݖY��\ɴF]����n���-�����t��A��<����͕Hx�K�;h^����`r��=���m�՗'�S�J'�4�( oip�u�ǣ�kD��Y*:���1��0�8N�a(����R��q����$��vD�����7�,���'K[�<�ɬ���4�`��8)�a"䪾���Է�u��:���m�,5�+��}�P��#SWI�I�^�ܱE��M����J�Q�8.(J��w�Id���4!�;�O8�M�U���x��f�q�P��T|�3������`A<roGw��#?�rLs�x��L�En�R���tz���7U����	�IBȐ��Mg����u����ew@�-�b�[7^��a��V�UŤF���R(�Ta��K|u}LY$��j\�v����m�c�'��w�iNG$�S��]��x �dǮ�5��᱁��R��5��U���>�[��83'�9 ��kS���o���Q-��R?4�>Y&ߜ��j3�O��j/���l2!�4���Ǆ%v��qr���3�u�^�23^"����[M��̆���m�j=��w�2�/xCi�;J7)��'X��6[�-�~� �o�co�����w��,��(�>1j=�9�a���s���B3��)8";hX\�\��D9Z��	�}q֧��'�U�c7*��3����Y<#o���\���W}{Z���EW=;�rL�T���i���� �@�:���`@�c�#� M���k����<�]n0��i��i :�ܡ,���̴��C����=�j'���p���v:���q�W��E��:��*˒%��V��l�m��?Լȝ�8��y-]�}�T
��j2jH^v'�Ö��S\ܢ)Z�`<E3�ZШ��Vy仄0WAhd��.J�����.mM0�{#�$���5!D3DH��u�q�륳�0�F�:U&�?�6���N��?#�L��@��)��2��~�jkAT"p}���쿿F.��>��'�U��V].�L|JpN�m:��M��k�ɑA(�5�H����!�1���D��sH���1jcP�\�2|� Ϩ��΀"�_Y%��(�`%qYc���ec�˔V�G�ef�� ���P5����i��/!��!@�iz_/�5���H
C%��_\�Pj�fɝ4�s��%�%u��L��c2p@�:�QCK��K�����{O����y?*┳��k��D ��Lj�p��\�߂�Exm�S
?����w��G3;w]�Zf�P�:-��h����˦1�u���H�2ƕ,�G�����mG�t����෈*D�}��]Ym���9�����#���W�� �9H��%���i�ɶ����z���/�#P��<��ʱ�vl�6��=�c�R��¨�g�~F�W��Ro��t�M~S����: �0|-�Lٷ���:xMI]�kupv�k�	\)�Q_]��%v>����mI��{�&�_�4�W$�E�P0�����rNŻs� �V{t�Ξ�����Gq�0:O���g)��hA#�@p��Z�)����q���kJn
C#
$�i~� ���K�x`x��%���������r�Wve��&w���ј���굵 � �C��fw4v�������5"$:�F5~��R4�q=�0��{9��H�2�ɿ4.�P�tA�m��g��6WSvMƧU���^��;�y"�o������G]2��Fg[s��S�h��֜d�&� k%�_�[�%�E��o5�[T����zh�U-�.�����WڛΌ�G�3�DF��`��0>��﷞��J���h�zP����V�T��ݱv�����M�MW�y�(�d4Z:]}���I�.� @@�roe�w�F�*��K����:}Z�+�M_H���C7��:�6�͕-ph�Զy&�>})T7ɨ���պ�{�{�{J���V_}�w� }��1�x���_�����)"��d"4'�r�T��hT���ZxP��}���{uɼ!�F<9�.$��o�	i&
���p�Pb�*��T�^��G#*�+���ūHJ���Uێ`Y�QZ���J�n�d�V�6F�"FͲ	Ļ�v�i����٫W?���j��9ݐ""����"��6R�F��: �0 ��=�arU�G��]�q��\��Z�&�9[}�v
0�h���Nu�,A��P�kw���J�Q+Z<�s��:3��Nq!��E]mù����5T
;��7��6 *3g� �'��;o���q��`�b�R糬>�(� k���Iq��*���lU�%��ȇ�� �q��'A؇}6��G0z�]xx�A?#�"z�H3�V��i�ϟ�R����:]F�H��ޣa
�G�>yC%v���QKx��H���8��F\��9�3���GrS��h
��Hh=矀޹3�ef��.i?�{�X �=r����せ��C�<� �Y|��m�[��d�g�����	f�y�;!Iǥ�� �0�!���l�(Ơ	T�p�L�S�F���b�^��B��V�g�	J��S�rז�����L;]�u��@"��������_�pn�Qc�����ߥ�ޕ���d���n���=��^7	�"�X�J[}K�N�� �Z���[.��yZWCj�ٶ��ײ1$������Q7����)i-P��%��b��,�2���\�����6����x�<� *!����߾�01�z8T����'��N�P��O���-�L������=!����nk!&ܤo̫���<��������YA�I�v��}*a�N��{QaYȘK�?��nR,=���IW1ʏ��R�����]�,�#`���.��H���)�F�S�-�>�do��t���9ji�Z��J�;R���d�yʮ��OF�+!��@��h3])�*�L�O/a��l0�ЍᝬA�R|c��u2��g
ʯ�U�:�'R��Ǥ�+��� �6�����m6B���0���@��A���AjV�̹V�1�/h�#����A��4u�&0�/���1���vz|[���%,�d�u����RFO��
i���?�>�`�C��ƾ
��˓�/���:��m�;�~iT�|zAw�i���~?Y?]��k��g-��x z�0C&s�/��2�ƶ�O�Tx�@oI(�mnTa^@����9/wF>��9r�k`��g��w�3�B�������ĩ��=_�% ��$�Ł��0�p�S%���T NMoL���lH��~�����[��Ck�Y�]�o��ɓ�E�g�X�,�/#a��"����_!�)�� /�� ���nHa��0@N}X�M=}��^�K��PI�QUwv�qyFb_>�I�f��°
9�����F�@4Q�s[�ef{����A��b�ѝ��J'��t��2��Rr�Һ�� I����ҝ!�� `�#U�͹��3�n�`!��9���x��IT>�iE�܃�Cϯ6 �����:�`�
�
�29l^��T�`��n���N��,�����1>���0� �fO7��^J�jCI/��_��2^H�7�E�qg��ݢn�P�'��j�����n-p�_4������`�O�9bJgf�2��%�ñRˌm���m��V���Q���8?���`s���_�E+"w��5'��M/*�II9w��4��IdЗ.
9�&�6�r+uI9E�˜iMi�a���������)jBG)�E)�b�6�*w�x2�5���\otV�������oe��~�	�l�[�nZj���!sz�\\�)*�;w���G�=҃S���xI���Hrj��������((�R�Tg,�z���G�EL5*M��M�(��>!��A*�Ur��M�3��Xl�^_�q�x �x@�7��0pt-�
ok�$s6���?�pi�+-<-фF�W�#'���o�������<� �  �(S�S4Y�����C����3@CPfA ���C�
z�Y7D_9Sc~Y`����A㲏����s�R+�;��Q᤟�$���$/� �w_9Wvإr�o�]��˧1x�JՑ`(I�>���]
���
P~G��Ow�yE��V�%]�")�u�������g�ȗ�aG\l������	��%��bEVB+/Kq�ϛ;ed�(;�V��󣘇�9�OH�,�^E����Z�g�4�l�m��/y���,^]:�	�[�^��|2�F���s#u	ܙD.aa��Z�A�#�م'E�׾��b���ێ9��I���4ґOEJ��5Gf'%��g[���tJV5����~���xw�x��$�2�È��WrIn	�n4�­M���,�=�u��#�����{�W��~�S؂����D{�|8��z�X���,lb�\�����v�ݑ�e:��>��{	&�8Ӕ�V�A�*{C-x���9���i���\<)��:����.�� �G��f���Ll� �"Tk���c��ܞvetI���	Rdw��Ͱ�y����P�.:�;z_2��5L���u[���݀�W������J�\6��x|"o���VN���x�(�4��b=�-��(���o��>�,"���}��N����O��7�s�[J-<A�g�[�U�\�[<�H�\��T5��Y�^�#��L���>a�h�p��"fI y3͎w�A;�'y�=c9�^�&�#܇\.�r4c	q�*g��޽�cj	������ 
x����]U�d7I�SayP�+�>r��2HZ�����|Z{\��/��hD/,�"Z�хv�y�R�;�*�U��nh��$�V���:4'�GI�4tO��9xD����*� �����u5�h�#¨q�i(�9��@�޷{]��Bt���1�7'렜!u5�N/����T��4�[ߩt-���AOp�o濜Ы�Hy����Sy��I>����d3?Q��������K�>pC�2%N�ԍ8�>{���7��A��%\޿U���|M�Kj�%\1t�+V\{�0���FW��"W�p��e|�����`O�{�z󟆸�?c����i��C0kxj���E��7���$�k,�[E���,��ݸ%�f`��*w�E��Dܣ�����U����Xc�Zl<k������zhp����<1����ؼj˴0� 1��n�:�{HFx��}	0�.gǷ}�̣�]E�j�O�J�$��*�0N��㨞����*���c¸^�u�[M�T*�X�ϚO�~d�j����p"��ہB4�L~�Mα��?�W����農o/LC�G{�H�B~v�
E�%����+()���d#�M�[f�y�xݎ~��C��aT����d�yv���k���Mo��ó!���]o�1���Ӏ"X�ߐ����86�]�30xoJ����,P\�q�]2�)��xE���f��P�}��Ȼ@�SC�(\-'qR��`�r��a1��M���]$��[�GO����0�w}�U������
�@n9�=T�nZ�`�~����߬����ӭo��bU���+�g�[�cwٮH*����GZ��D BS|�d!�+B�^KνfRNН�]�7�Y>��<C� NXr��h��j ��̨�O�|4�YU����M����
-��n�rb����$O |�{��e:56�W�7h-�Snڧ�E(�O�[(*���6�F���$�I@w@�����pN��{#q�-�?�h��GaۍiE#�vs��˴h�P&ߙ~nb5���f��K��sJ}I�y�����~��b�݊o�kE2�z��e`��0��b��Z�����"�~>kfB�W
�g��"�Ԙ[Z�P�z�L�>�q˓��N�b�	u%�Q�,��~ ��[�@H��n0?����=�	lrd|���s_�%y����Lg] ��E��U�<(�pX�ЭOy���d&�xi�+IJ�P��Ȫ;X.{�vu��@c$>D�I3��C�T�������1@
�����V��(��N�&���s�п���%>k+el��bD�-KZ�.YR��B�) �R$����M���uC�Z
4LL�,����w�
����H5`��[��6�k�Zs#����	�䝩���?�k�(Y!�9L+��y���h}P�����f�ȐtH*J��ڂ/�����5��W��x�����wJv��Q{�z�R��*$���ϕK��
d�=Œ7(�xf�k�\)�/���٣�"m����w�Ԅ����g�����m���'����QI���W�	�A���=�ğ�(l<����">�6����s3Z�4�c0��Z�r�?��5��E��.��i��=�v��w����� j=�˖	T�ݗ���o��k|e�!���#Ny>ZW o ������}@9T:$��k)[�Ԧg7�y��Me#Do�ڀZ�E�wS[���$������'W6���?|^��P�`+"|��&������NܛՆC��.���W��-W��g4Q����-�$k˧wP^�`99h���'�q�$ןx��b��R���lw%	 X��L܌X��ʥ�~��(�aA;�c~����_�W����%'wd+�:�ګ�j�K�����n�L!=񤒼_�m4�+���aB���Ǖ���G�;ad���f��?K!T��T�ngO]ЙD�"�K�>�ɫ/�&�f/��	��m|	�>S�D`�m�D�����G|Vz�wxJL'	�wWgX���~U���h�H���B~G���-ir��:�l��ي��sD�r�e��4#2~��`�ϳ[*A�vk��ߙ,��aqh��U�z4�Z�?m�e=E屆)NqwE�Z�)K,���2���d��=Q4��L$��)3�̊���Q�#�$7LR*� �<��Q=�Ќ����Z��_���-�_��UE|��cH��l^+�w��!��Tc��ѱRF����ۻ.ȱ��Y��!�#�@c����c��=O�+�EL�V�&֑;�5ic ��}z4
�H�82�#	�S���� �F���3���I��*{bG�+teQ!$�u'�����������T稜�̴���`�c���&p���b�_��C��' �J5C
�"D�����f����ኺ�B!�4[�m�6�r'j�(��⻓5^铢�Gu�Y_j�������o��Za����9#N��^��=Hӎ^�\L�;�'M�,|��s>\x�KHi�S���qt���.t��!9@��xp��9�*H�Y@�.��T՚�W���&���q��.Wo��X e�B�cv:�� @���m'8������d&]�oBɄJ�_�>N��:ZrH�$�CE!�IWl|	�_�,��|���v���6�d7�"��
���2��/���)'�U���&}mY����
���e:���q.o�@�;r]t�ec_"qtb�n�����A}��a�r�����.��56Zwǀ�:��]78a%�wC���$|�2�c�@/+z�-<A�>���>�je�I��$��c^Ȅ~߽l����D�:R�ԍȞA����y�����@�w�k��t��?����(A��/le|B$%�X�X"����� ��[3qm:���
}�ZW��9~-���}vk��. N�!����O.���=�Um_��P�����5S�X#�|7��.�n����%F���h�����|0W��O[k����y��'�|&R抐J�.�.wG�,�߃ڕ�g�-�m��2��gh�A�0<�g��q�)����t}+�4�(a}�+��]p��;=��'3Y�%>6؍|�ZM� �Mjَ�ҩ�Ȩ ��|� �5��{�� �p��3����G��Ȓoݲ������'y�����
q8+�f�_G�S��V�p��BǱXy���:K�M�i�!�v㊡`���}+���U�dY;R��D���*�����GL}vLo�Ve���*�@lA�1�ߒ���+WC�mU=�e��Oi��������1CUz��"��浛Btx�,<�c��)-���C3�cn����;��a�Mn�&������@��c�tQ��u�V�
�w_g���n���|���L�Ykf���*v���$����2�_�+5A�
U�v5��e�X�r��g6�=_@6�XB!p}�5G�� j�?�MKKba���FG3�^ ^�y��}�yPj/@��`���k^��	�j�:�}M~�'S����'l�$��� ƪÜ{ג�ۢk��}�
���a�e�d��}���Y ���b�$��g�I��Ll����	n�����:��kް��i@�M��YEn�h�ly�-�_�U�e@�vM!kk${�\��$��6!*U;gMq�bڪ��T�XD�,�΍g����2��D|_G^��(����� �繷��8u�z���6��壾3'-��&F���ϬP�	a����%�F�P��� ?�S -Z����)�����Ĕ�� �����f���A���(��k��j)Z=�K�	�rF8m��4������G����b����Á�oZ�b�a /(�L ՟$M� �,�g��l�`�l�͔2L���o��ƹ�}�bz��;�P"���&U
��a���6e�g���f��_1���`uT�p\��w ��۟!{5-���Z���)� �g���ƨ��X	�?}6#�h�3	�z��)�g��c^��9�e�����$�@L���F��t�{T����q�j��*���4ځ�^���5��+��V�
�9w-���+h�l�|���(���ZVʅ����FjS�1j�\���Q�{Hɥ?G!�]�I��w�I_�c;���w�����ͭt�ο��
k��2|��H�̈�([�D�*J����Z��������iF�����y�/�ɨgl����R7��+�x��E &�R��"�Tdq��os�c'�hch�Fxߪ�T�G1�2�w��B�5��{g�/�s������5Osxo�b�i�]V�����h~/�� ��τ�Rm0�R�BګT��F�\w��P|�]!�{/�5�us2i�������}m}1����!�{7zK6A�/��:,����%b���[ſ�ШP��௤94��FP�xeL3�s�+&	X��?��a5QqRG�H,��~��
�b*��h�E~e^�7H��9����ҫe�oV��������K��2�h�USY{ ��<��5?��l���ȷ�k�|UY�̉�rv�7�R�C�N��h����<���pޮ������֭�a�ؕ@�uos�h�2��^ʠ��9�5�q��#
���	1\��x�m�r��>�"@��������{���]��Kio��'�W�-�:��8;�@����(&\���XAz����;���h��rGB�)�;����	��
��켹0���"���kg���#:,d!1iӕ��ca8o�@�=Y=Lo��4�-�pc��,�T�à�֧w7��/�ex�"����K�nw%���ɽ�:��\�j�� ��z�JX��d~$��CgL��W:��i� S6��=���y�����K�!A�
�ߏj�.�T7��]�zNm=��}`5�u�3�o��p��^�Ǽ�����3��s}"
?�Q�J��o���d8R,��$���w�M(�Q���.1&���8[��2�s�f��q��KRRN�����i{P�����Q�k0��A8��U�x��4[v$d��[����m��-��0)� �o�ոJV�w���0i�t�myp֩9�<��*'������E����.r�r���;;H�`��/�6.��*,(d��k��c�o��F�<�&Wr��պ�n����*ǅ���&����}}�AVk'�8����[6w��.�2h����[(n ��0T�)9
<�L5k�:J߬e�pn::�`���+�5M���3FQ�$c	�J`�Z�(ɹ�>�i�lQ7��!���{4`C�Q���B�0��lP�殴6��EH����|�=�
�X����i��H!W;�a�������t9��!F�O���1Vj���Z�料p�)�ym9p�i�1P�Cx���)U�6�XVe:��� �v����S�ەY��6�vf�z9pwO�����T�ߍ���嵦�,\�R�u��/��ʎKA���|���1�VR�g�=���l<�Ҕs�U�--CT�C���L@f�� �G��������V�D�d����:F��68�\L�֮b��E���a�{���M��:=�zm�p��y���l���yDqp唫�g1���iEֻ6l��?»��p^;n�͢MM���)u��#@˱3M�q���eŉ�)����X���0V�(F<��}�=��Z#8�d�����u��x��=>��p�$%�-wK��S��U���\}x��ih��-�F�IN�yH9�x���%U�9B��IWd�$���;PΪj���K�Ytly���hq��.q!��Ú{�(��&��7ʠ�!-��KP �֊�����F���kI@�C�C>�a'�j�7Y=L�+j�K_^$u ��� �p�������	�^�/�Έ��)<>r�� q�������,nh�&�V��j	?��j��;$<x��C
��J7&M3����=��wrӼ�|v�EU���@nu��D�]�b *M���{��0/XɃlV�^y{�)��FYu�I����1(7J�.Xn����c\rNڸ�����m_����m"Λ^�<��o�!�(#�RX���`�����_�����/�:�h�c1!yW���ƪ�����z̛B4����]`�d�X��:(����iZ���Ec��Z�uDQ
��$l�7�.�3�$�ʗ�T��)pמ?[T=Z_����cٺ�<�����tRY��!�¬'�\ĕ�ٲ�
Y�p?d��b?e��(dF�`b�Ċ"1����g��p�����XȏU*��$�u衚��7p���VN�n��s�J E��Q;{m����j���V�Op�(Ň�d�_������h��ũ�ugx�6|K2 ���Ͷ���{��}��S�xk3�� ��p:����D�C������햢gQC�ě���l8 A:I�:a��M��?���xt��6!4�u{M��2k��'2��t�� 2gD�`/���)�+��h1���j�Q4tB��/aoZ&���Uh����7|��9Āui]�b���k���b�s~0��w,h<��C��8-�[f������U�v�p�N���%��"Cu�qf�S�ϲ��3
�Ov����Cp��o�����?�Ȋ[�J7:H��k�粛�dj¿�7p�Bn�:qo�6�}�W�ߨU���"�쑼��4�ie�)�(n���B���D3�qM�	��%�z��G���l��}Ў{�b]�`���{�. �q1`��ͼl5�W�=�*#��Xb
�����[�m�b �L���:xA�����i�������n�]㽤�+�)RZ_��X���s0�/_~����K״���f�[�p+L�?���Gg�L��r�8�Ǽ�q�`&�JZ-%N��$.�C٧��%s�&	,av�+#��_w)Z���x|����� Qq���8�N�tZ��Q�G��@��8ݢ��y��Fm��ٝ�i�5X0\����̝���zgugM�O�),C��w�����1c,�W�m��\�+�}E��gv��:��u�"ccC�LyD�\��d����np�棛ץ'8�{�Ϲp����������,O#�/K�G��!d2a.�ב3@S��:�UiRX���
J�����.���ݵXB���4h,+2HSR��#~ub���˜qm�Rj�8o���w���,��BTf���sYg*��Z��8:�ۆ�PO[���!��2�������J6���y�0�G�c��T���	{�B�s�T�ӌ�o��}U�J�O����dW��R�,�!���l~����!����u�=�ۙԫ��>�` �y��&i6��U�*iN5���������I�N���l�XE�7����%�{�D��NkI��;�B�b`��!7�c�i?"���RjO2 �\�LU+Hp#ۯ�U�[���5�Z��(j��m��[�K��%��<T�NOA �����4��ٍ���U�05Y��\��7�Iw<�*��J(�؈M�2�rn}�u.���3S����ի����_!0s��U�g=�ɠ����&�\\�-� �U��c=q
��zk=�5 ���#�9t.�0	��h�w��y�w��;�"W���D�E��^Qp�>)=��V���(
X`��Z��`�F$�651n"j���E0}�����q��y��/�ޮ���Bq��ZI�4)�i+Ielb�Y�D���98�����	����He����饽��
R�@ErS��&W�(+����E�>8^�1X�q��G��v���&�Q G�LFr�(�duORh���fM&%���T-v1Hz��yn�[$d��Fw��{ �}������%;PTа��}��ϑI��R1��{�����[E �D����qe�` 4�����~$ZM�zD]��e�"|��d���e%��I|������e?��+��Ҹ����\�s5 k�0!ytꝌR�5� ��VfmJ�n\L@�n�C����FY\3iQ���J�ҩ��醵V2�vf����8��s ��>�Şs�f�J��zl<U�A��L�p�ao�_�K��3�B��d��vMߩ��'tdmn��k���J/��q���#�� 
=�:�$>�W��L���/�H3<&:��jn���0�R'E��k��l�x��WKz6��\K���~g\��S"A@n��?��dp�^��ȅ�M��@Ӟ��i
��rEJފ�ǹ"�}A5X燦i	-BHjbA=��	�C��~�<�_a9Q����* iHN�%�E�L5{�ޔ�D-Z⥘YՎ4���t������Ѹ��ֹޯI:q�����pCb
Q�WJԌJ���E/#����Z���UΥy5Ũ-�{lWUWc�j?IqE]|��aM�m��x���
�
[l�l|,/��U܊�է�H�P0B)��z`O�OQ�?ϐ2o������ހ
癏/����o�K�Sb14I�*
�@{��P�����W�`:c_j��ͺ�%��
#4�����<�Z?�0`ˋ��yo�����e��m�+vD�|�����VB5D�"V����)ߧl�[m�jj�˱�����c�_X�F��N}��8��;�zL�fE�( ��RH����Fƌ���y��