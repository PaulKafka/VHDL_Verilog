��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ��>�(Ŗ�6�eQ�d*e��!i�v�4G[�\)C��S� y3�Xv��XcϷ�z���B�}��uE�Oz��q��̷s��n~܌W2����C�x��.ם:��˂S	�J�����ڐ�
�^ �	s�'�%���gM7�� �7���8�߻�So����@��>#�wiE�]�Da\E�ʙψ"�՘~z�X��)�f��D�y&�-��8R}qI���=-@Z.�������&�B�p4Z��q��M��c���j�R���AFW��\�T�Ɏbof�#<Y�^��c�=�|Xi�/7��� �#F�	Z�om�&��0�{��Ph۟p��_��s�-�|3�b����߻Ș�2���U�L�g�'Ň�&����!q�4bs!�V�#6��F���BGo�f�y�IU�o-(ޡ���W@�B��,��T%�*�a�i���jӄm�������H�C����ޟ���u2�g��'�Tf 4x��7�c
�^�N� �rR��/�7����n�U����'��b(�|��*U`�%�U�m�EQ����n���8���!*�O���0��3:�q��D:	�]a��N��^�Sk�9o᥅�l�SP��&������<��a~��+���CO߿EI��M�	*���tQ��SP��s:�[hl��_q�1��Qcp�?u�W!L��ႲW�Nïy&`�;KrS�6��5m���I#���^$o��0]�mE�FH.I]p���K3҇4���R\�7�^��	���
�E��7�w�,�$˱����eΨ���ow!9�����y8@�l��۷��7�:#.�A
�/G�e��+g"���BT�w�W���s�x�jgW'욦����/��@g�}�F2��w(Kzg�؃ba���*���������u����h�`]8x�#2jx�I�Ɨ�
�����: ����t���4NU?�S\�>g�q���3�=���Y��%X��D�F_�{�u����u���� ��v^���p���5Bp³�"�
u������W�N�����.�;`��+�ߴ�-;,2��jRQ���� Ȳ-I	&9��w�������W$���%^�mwEA��&=�˷���WEx�2��#`PJ��U߷7��gA(�)�D��X��M�9Ap9x-\�͇Y�&cbc�X+V�'+3���S+)�';���f�k�T����ir-�IA����ϑ�%�3.�{�SI@*>ϖS��!ԯ�k��=-���,�^Z_6�B�z+,-=�� ]!�L����g��!���<��~v�=cz;Z�Ո7��-5�;f툃� ��w�~,]p� Qn!�����F����=�C�yɀ�e_B�����2#�:�%��xMi� �sT�=�Z��CWy�cv.����xF��5�$�K�˘6ᖷp-W��T�8�����n����U����[���e74Q��:�:va����y����~9k虯�h�
�Cܳ%/dR�-�ͼ�����Ş����� �)���&W�*�u��#��[�i����7���C���&�X�lT�����Fх)�z�a���\��S�R�6���}]��m#��B��l��Ҿ.����o�FrZ9�٨�K��n^��Z�EFGx,ht�+65�&�b*ǂI�׆��"�X��O)��M�#VV��C?6��T��� .Ԍ�R����_C�e˲C1w͖#��g�u��n��x̖�{�[��t]�s�q�D^��h�soȃ`�V�췴��^P�����I5c9c�Gg�B3��4�q���ĩ
���;h�:�%\��琮�����E�v�����{���q~��,l���<��K��P���WL<��+~�e>N)R&ɷ%.Yˬf�`?L��IC@�֜�L�zM�Gu�4w�ҥn�?5_{�hG\��\d��qB�Ac_�>���zFAW�GpGL�a��L�Ÿl���y1�q$c �k�����}��
yo��e��=A���4�*G�r*w��m:�6<�X�T�I�s��L�#��-׎D�~4��2�Ye_ܸD��J�Z�3�"�L�(�%kr26��
�]W53L&Ѡ���6/�\=��/��7-�$�t+�}��M"��{��D���F�r���̱R�S��e� 8|'��CM������q��c:TKq�Dx�IV	(��
V\9����26��+��ب�db�U>T��ĮQxڒ��Z{<�㒩�o؝�N'�/�$\���7�F�w�R��3c�nw�,4%�A�Y;# y����H��j���T,�ЩW-~�G���s���ɑ��*�]�6w# ��>t�Ў�Sؐ�*�#���y�G�	~�ߌ8���b�@�ƥ�j�I��&��Gb��l�]���ZA\��|i�p:J�R��\��>��ˉ�y�Ϣ�P�<Z^I⢸e�tM�1���J��K����"}*���]��������f�d"��Z��1��r�E�aۄ��Y��T� ��g4K�Q�=D�&�\�uV�.�qɪ�xJ�#w��f0/g۞d1�i'-Qb��~���8r�H*��W�V��;*��Mt��_�@�H�e�F� ix�s4��ύj�۞��1��FU��C�,(q��+�	��J�UFtڞ�Ih	��ݻ7S-�-��Uv,�I4f!N�pc0+�@��X�K�n�S�lf >l�Y���̀ǈ3��eazʥ�c�˾��ɮ� �L�&f,���53D�'�����ׯ�N��8ߊj3J[23ɲ!�]F#�f�x��`ȥ���B��jg$8���F��b���N���c@��n�o��c6Maq[)��ݗ�,T��z��͋�<��Y����=ť��ɹzbw��I�3���x��}�D�Dz�w͊w�-���˼��mG��#����A6�i���`���1��)6��c迪�s���9k��1I�H�G�i(����oh\/b<5s�4��/e�pŷFQ� ꁱ+�ȖA��CƁ5̶���}�V���k�|�艛��eH�4NXl	$SL��9c�8�侶��4��w⟰�WUW��ol�9eS��H�"Q��g�1j(�U�$?�oW \�MO6�:o��|�=x'㜑�X�C�{rU"����B��iJ�|�*�cŝ�(�31ٶu��E �X4q�*�Ymٵ�a�(d}l̺����u�#"ny�"
W a��>ͦ_�./�nUhO6ʙ��[k����q�x��z�Ώ�,��(B��0r���k.��-�.��ΪI�"Ֆ�\Mjpy�˹\�\�ޭT�Ք� 3�NE�]��y�
�+e��ue�P����L�rkR��_��%�A���Vr7y��{�XWd���1����a��X���F���O�9�?4�+�֐b��C�eȈ��'���g��3#'K�u�Ic�����L.먖	�6��0[�J��bzb��q�1�T2�&�~tI�s�:���P���F����!���y�;����O�)��vvse��u:�g��T�V��TX���dza��2o��h
����5ʅՇI�b���&������P�38`E`V�_-,l�M��٫��n4Th���d���*�����S�'�%zeO��'��J���Z߶3�ZHi�+6�G�j')�%{�{b�7[�]ёdo�v���!�1}�S'^���L���"փ�5�TIhb}&���7���'N�Z��?�	���+�8�QE3�rz��-$��Bl���/q;d�V�$�d�?� Vtw�j���<6VT	��H��iQ�60Qlj,�FV�Xxrnc��#)1I�0?"�����1�@d��A>�֧ ?��o�'�8hr�q�l�8ո���2����}!h�S����xT���=M��������q�%���a3q�bA���#g��}n�
ዷ�p��w2l�o8�}8iZ� 5���<x�5��:*A���ξ(�bi��Ӛ�� ��e=�E���G�qh���2�=�1*ǥ�Q�ռ	ΖV�e��;{�ĸ�P
g��q�[����J�-x>xs���ۘ�:$�}���'0��/cL��H�xO\y�ý�K6,�9�����@�%�U��h���;���U���t��n��>I�£�����1ϵ�GH��7�v�k�©o��,R"�M���v�Z��\�� �u���#��h^�p�6R<j�	s�}�W��CA~/4�.���M��1k.|x#����j��6��>��.�>|-�=رN?|;����K�;��H�BC��U����怒�H�H�3.J6oػ���3y�j=����VIIF�@ѕ��oܐs�!��]Yґ��9����s�9;��jc�.���|\��
,u���Y��:I�s9��*ykf�oG�HoO_H��å+�A4���6	*�[5!o����4:6����(<�5ڨ���Ao��T��cs�HE�I-a�	a���^H��a<ot��������t0�V�P�{>�w�5�[���<>1r3M�{g[��
	�2�/΀�!�Dr�f��M4Q`}]���u���M�>Tw˭��s���$�<����V*�OGd8.���`[]y+K.��|i^�oT�mɝRD^�ci�$D�2E�B]�����l�	�
�we�O�AS.sIb�@Q���9��#����z�qR�9_T$�OaVT�^&Q�w�@݆��՟�?�)b���g^ ��	ԗx��8-�K8��`(	j�*��J�P�)��D�j�֒I����𥮵 �cqD�W��k��x�#G�4A�o�ym=UT[���E�'�Ƈ�$�7���f��Z2�P�'�v䘺5�/	��^�=~���8J�p���.#�� ��B������T��pF�u������cG���uZ
Ls1�/%�`����(����Dl����Y��r�nY������� �k���N�@K��Y\/�q
�8�M�~������!-��7��|�cDW�x�@��(�*���y��1�U�FY�(剛�����ٕ�z3�@-��ho�>h�R)�L��s���R(���KS�A����t�J8:��,u\��x����T��N��N�\��UU���]H��u�1"�F1��J���?M��!pd��F�D#�R�5ˡ2;�jA����B��j������{?`-ּ�a-qN�lF���c�m�-m���{�՗e�K´��3����
��xF���Y~h��䳽xQ��ѳ���l�9"xc�񰎋m&��O����Fk��?�U};^ׇ����(���؉
�������2�Q��Wu�g���}2���B�+'�r(3�UG#Ğ�Ǻ���
ckC��g		���^�hk4�/l�"_�oI��ҋ�b���굣��^�4�6�D]O����x8������ϐ�F�>�4)�C_��S�����K�3z�P�����r��a���?�؀:�ʨ	 |n���#y��3�N�z"�����:���l�]����:G���Ą*hDc�隸4�̍�c�B��%���}-���/�|���/Mxi���XI���=.f�@���
1Z�ҙ�FA�ƪ�r4m<#�_9�S�o�eF@0�~����p����޽uﳫ����u��aD+L�@�9&My���V(~���h���7+�t�ާ��s.�8�+c1��E��� Qg����W >3��%�*��0 ����0���}�o/
�1��d��B�ޚ#���څ���S}"U�@�U������ U���`�y�����!Z���_���5em��,������u�%��Vԫq�ɩ��Y."V
JC}C��͂�a
-H�RҔn�e%`=up0���� ��ܫ��RQ�9w\����� |�;���L�_ZW�qX�ehw%E�L�04�Ř-��rF��� ��ڭ"���ߥ&J=7��`�;e�8H�&H<�\�	���9�$���+�9�_^���V��0aw�K���mk��z�����s��?�Q��MI�71����@q[�ph³��s��ZU;O��_�B�!h�r���π~�l6�T �� ��x����Z�IT�C'�_0�c���$9�\T4E�?�6�j9�r�s��H�K=/p-U��*�*��o ���.��N��c}�
�� ��X�k�K����Z����5y��:�옴3j�Fi7��[0M8���'`����I/H �������LI"����RI��ȓ#�0;k{�n� ���|�R��~�M�q0PcW@��k�6��$��Uې����;�vr�r�+��bl�i�5����&�����!�{K��V4���:}���+��0S��^kW$vإ�]��	��C���ؒ-wg�w�L��J���wFR�XUA1h��{R���{x�_�˵m��L��db� պ�,Δ�d��z?E9S�ø*�3)�s�/7��	��{��Y��U��f�Yw��aD"�<��p0O�WT���E&�x����e�Eaܲ��|F˫G�ů��('�+�vj<����)'u9x�z�x=��k.�)>�cx�"�WrˋBS������h2�����5n�x���q�����*׍D�`w��M�n#�x2����g�ا4��;"�]5����F"g%)U������7]�@3�¥;���h��H����5+�\l�q�B#����S��Ko��+����LA��d���8��N��%�\�ڑ� �&��
X��<�M�@��� �C;&��GlW��1a|Ni��^�cV5�bgu5������iߊe&�4Mޒ�:�=b�F�Ǝ3���,�K#n��ڼu�#�Ӻ�M/�|G�������ꣷ��,��ӟ�`�X�r�[R	8��iR�Y���&�r��X�ʲ�NV��k3�X
�4w��Q�j�}gb���sޘ.mh�*�k��7����T�(6���6�PWG0Ufė,=���?�zJʢ�gǤ�K�!/]�A���L������5T�XL���/�S���N�"�z6�#R4I��� ���x�@��ȳJG���ԙ��L�t����f�'�>eg枎�Nw��A>�ؿ��D� �ӏ�"�O%45�n�C�6Rճc���5��9{���M��2J�"g�
ɚ�%jt�&|�zzJ|�ߓ���<ɐ��������V�U��,N$T9��V��OK$q�5��eq�A���x�_�B˚h=/��%C��!#9�����2����!��,��)�� �0�u<�Á��Z�8ֱѨ���생�`���Ьꇆ*z։5 ��*���2��'�÷�:�0B����(�$$��؏�OJ3��U:/bûl�+��_O�y�y�F��{�I8�^����05�㦢|Ҫ�.�򖓝��mr��Q�84ƙ�ꉦ�4����s�Eur���K�~]t0����'���9O�=�y���յI�9N��m4���Zxs0q��7cOG�~յ&�φ�!��ƨ�\�ì�Q���(��H��K���̟��a���'5�$� ��"<�uΥ5;Pm�����&w��,�Į�K��}��D�S4HG��-�j�2}�V�5۾�ʠ��toc�Q^.���!.���������G�HdX���A]	�=���Gb���&ky�޹�L��<�T�4�9��k�I0̞o�;	�#���*��޺@��;�m��\� m'"򧵇�/�%�N,�4���R�cN�H��`C=��5�%&OQ��V��@f#m�a�2�Z�2�� �B�ղ5h��k!ѓ͖����TL	�]�gh^/M��F��D�|�{@'��U�U<Jp�6		.������D
�����@��:F��avSk.�j&*D2+*e+I��C��5�!:F�c1���Ҳ=�:r��&��R���4����֏"m�	��r����q��-�W ��g�0oI��"��ot�l,�x��0-���V{� bgژ�-�&&��������AR����ί;��~c���z%K? � �lo��_�N�V��<%yF�:�:TF-����cx�z�3���t?RXA��බ�:|��e5C*�Wbr��RxP��˒���O�3}�)A�Yq����<-$
e)�]��+��vUg��LPs�| *�������
��F��+,�`���C���@�,
�� @uD��q_��Ě���̩�D�ًo'+e�8p&����JmF��y�%��-	ܖ��G���\��l=�f� ����L�f�]$��r\�ʬ:�3C�l}��\�� ��z�G�!Y$�aEs��̳��
'�Vf,�^�+�����u�?�(�'����b�ʊcG���>�A�ءs��?h�S�6]��}E?;"�*I�����������ϒO�xӜdٔo��Թ"��@�3���ܷ^ɂ��k� ��`�yv�SJt$#n���$�@����>*~��;.vìݹ�Oh���s�mLk4]���n�VҘ7n�P/�Hm
'��+;yV�:4(Am��G�Hߊ]�]�8 Ezo�C7JK�=��,O�PJ[�j�7rQc<ǟ�~�Dȏ��sC3!��o�,>� ��Y�Ň�CR�峏H�G*�ǁB��W�ܐ���܃$4�޸U0��1����]��l,�6݆."R��ܒ;.�+8���X N>/0�;��'��05�B5�h����'B-�����x����\Z;
��OU��i���P�A��O�;34���V��e�����H�^4�q�Jum�ه�;.�m�x'A�^�q}��;���M�3R�=W:�{�2�,|!� ��I�� ���	s�c՜v�!�L�-N�JO�=���!�P�JMd�Ob�g��9�i5
Ju]}��HU������AB�E�a��R�!�~56���dkh=y^ߢ��T&5�XT7�w�/�����E��0KXW��_�'�j6��ϭ6��*�';�S��������g(M>F���̗��'��0��1T�&�Ɔ8I���Z�	�����	�_��il��w��tm�i��э��mD���s�F�S�i4}�vfI���p톇]��>�q����[l��HzFlD�1��5!���/ʇѣ�O��b��W.��<��؀0۱�'1X_f��<o��MS.�z�зZ�����&�x@����)�Zj��^���w�8�����3�~-���������1�J�S���W��Q�X^��	�Kvm�o�`cbk���bs��8�AA�xϊnO��p�A�!���'�W����{4Mَ�&�n��'�s�9��2��a�n}�d���O��o�}B�!ad�(�9����-�.��)��Ɛ'��[=��oO(��Y�8hL� $����~��N?�H�#|/�H�%^��Z�v�Ӆ��,�"��a�`�� Ҝ��"�*�j��$\:���:�e���<�|�w��\��D˕*�:�	���Q�/Q־)��	��IH-P���	e��T��^�w'B�+���~��A�}���%��S����ٖ٩�L���O�?���~<�6��@�K¬�$pÇ@*�ns�M�r<$h}
�mi� �h1h�iMG(�6���w٦�'~WMʳ<�.�WypRB2VD����
1j �����z�8���W�K���bOr���!�'����6x���Hm#�O�*�_��I����z9��Z�F�J��EMJ�]ڣ�_�1N����A-�ӄw��|=00w"�	u��C8k}LȸE�v���,pLx�Hſ�(���	j��P3M
(M���3��<�@�0N����B��Q,��._�~��iW����\)�!a��/��/��d�+�.ΰ_���P)P��N"�����h<؜�|8���/�2WB�p���.��|�D��Z���|��@�pD�ԫ�67-�E������ A���8���q�Wȱ(&H�T�����MV�	�$��1j����B+?,y�胖g>�� cj�9n�$���tэ�Sߏ���}:X��V�����$�,q��D0�)��G�O�WCóui1�
;��C�^�!�����ˇj�|������ZI�ۋ�A Q9͞��o��(~��x�ʰA��:���r:."t���	���YZ�C4F�w!�>/��c�����c�E��j�������:�l�����Yxi���)�Vf��r����[�0��5���k
1��^�<k��W�D���T#�q�'u���9JH���u�r268&�:~|��Y7~}y�����W&�i���_�.*x�`yV�sM{u%q`W{�q�t�Wi*�
I��wd������s��u�fo�
eO*0�e�I�ޅx��)MFv��������s�(�&���#�J���jn���̑}B���tG4�}=�񨖰�T*���ʰR�D���Or+�4p����� �G�'3ɾ��E�-�.׈�Hv�7P���*$h�o�u���c��������4��W��H�jNѝs�֩���{)}���[%��>�/� Rls�:d=��P���Ha�5�"�1܎*t�΅{y��&��X,g�MVM��s�C�A�4�fO~N�S.lӕ3Y����A����c��̢D��C��Bc��_g&�,5!��Ě��V��aL>y��7(���`�swt�pd���x捺�<�i�G�1x������&��NU����*
���V��S�p�>H7��	�O�<5 ��R��&*�2{
HJI��?�ԵW`�}��9�� .� �Ե��������'n��;c�`UYU�Hћ�D��(ntr�y*�W���3Bf켢{��q�@l���ژQyZ|���h{�7+`�VJ|H�W���?��%��G � �<�Mw{~��V
E�õr+�����{˧�A�e)�� ǣ��u]�h ��c1@k����/�L ?i���]�yX�~<�FL�	?4��R�-�������R���4�u�҅ ��$E'M����	V�4U_�#�?�\ym7uo	n�bx�Fp�]�û;Z��b߻�63'Jj���@T�U�ya������^lg��8"�kv8�|.�C*-4_��b�/G�=����$�>x�&:��\։�OAEl��b�A.h���R}����Bo��G�����HuR-d���m��X�wj2%�u �Fb����6�xͧ��[��!�,�(SyN�y"��!��&#���?�?�jL� ��g0��.7j�C�h�0��S	�m����W�C�3͛n��쯷D�ϒ�1�{�ò�m:��������i������g� �Za�I����/7g�Y�t�����Ybe"F9N�^�.�����h�aq!�-���p�&��q����u$.�EG�"=3I��!vG5U3�נ�;x��=�P�Ŭ�ЩAz
�X	ܠ3�����T�
"�Q�!�spcɻ�'D^�R;Pֲ��ED�Sw>�+2t3�[��u$-�Tm]��9#�!㟖�*��@T��T���v�ν�J����=s�ݰ���9����&��5<�>+�+J�ZH�3bF+���*&��O
��^���������&�Cg�v�Zc��X��?�58�FP��w�v�+� ����ՉX��jB0�V�{�E�����x�-ӿ��c�6zý��Y���}_����� tH�@�[j�AA����������6v���ۥ��Ilr��k�Q��>C���F_dv���[˶ɧ�nþ�,����ay�!���ׂr:�+=��rr���E�˒5y�MF`��0�tĖ�7����n?������%j��E%g�yc@�0m����բk�\pPr������Ŭ�ly�G)���%����V�ן���W��bB�z�#K�鳦�8�K<����i�� 3��)� �?2<���Cٷ���$���c�?�t
���,ck��D$Ɲ��bWj1�Qp��xW�/JF�@.�0S��@���ow��?�f��Ak�Rʒ[BZ�����5Wk��K��.�n�yD��W���<�(he��Q�aIЀy�}|�t�b�Ћ��)�b��pʻ̲|�H��Gk�<�@�m�O˨�O~�|bꕜ��Wgd�F��~~�jC��֒���(��)� ��QOv�-o�Л2K�*��uC�b�2#��
�>�o6*٨���{*��(�hsjʢ��+���1c?C�������~X0r��x� ��MTc���C%�5𢒒ٓt׽a(I�+��Y͘7��w�I&���P�ꭠ�o�.w�f��NE����C��Q��џiGM���z;:�yZ ��tcZ��;�?J/��&'h�cA�fJѺ��ޟV���.�noQ"�����qx�k�+�Q���3�� yu���f�?�z��]!�vv	�1[���Vù��v���z�6ʲ�*��!�\-ΧG�]9��ڸ�P��dH��ֿ�����j��&��N��Ͽ�mb�N>�A$t�����C��m����~�R'f�8��bN: I�r���� ��&��:i�\]������?�/��7�]����G�z��TЖ���墔Z�r�F�Z�Ӯ�T�l�?�*��?��1�|a����̽�#\�C��Z�p�2-���9�vT2A`�5�1�� !����,D�?�K#^EPJ�o�B�J�EG%�`�\����͢�q���)Ó��C��w�V"v1Qr �{�J���3�T]�;Y��J5�'��:�k�΋P�ڸ����A3���o�+�_i1��$[P�gh|��i�����������Ŏ��]�>���brH$yW���.��Z�Y���*�b�����!Sf U�����O�LB�Eh��N���>��ߋ��ZPNˋ�diƴ�z@9� :��wOS�����8iեW�a���-'�[�I ���s=/w2����J�]�ܗf�D�t� u�1?Qw�;�a���Dt�ŭ�Xgͷ4���)w�"�/2kW\�yP��{��!����'+=l���7��,�.�}�u>���)�ǵ��� ������T|5oLZ�2s������Yn�BH�W�-T��#�es"6������5�I����|;-jA��.C�6'*�;��ۃP�iz�i�I�K�[�w�_V���{�i��:��,�߽m�.l�6��oZ�t���)�b+�Ggr/������8�+*c��CĖ3�����ĸ�X�&LM�pN�ڹ�5��<0�A�aQpz@�k*���!��(&W�ƌ�a�sXT���}��/T)�8rRQ�[$�J���:��R�.܄3H �j9���O<5�W�h'��)���8����.��B�[D��N�^�Ѿ���0	KY,��/)�!�/��p<I �ݭ���|��Nt=�v��S,M�����m��Y���W���ou*֜������ ̷y��	z�^���%W�\R;q�ƃc=�����r��W'�����`�#�{����}���i]йx%�;�� �u� [��%r�!{U����']�r���(��~�~�?�4]�J���@"���$T�\��7决��i��_̿�� �>���D�S�h1���cAo	��B�� ����GV�ܼu�XnI�R�q��U|;L�g;ӄ^B�z	�_T(l,��k��W���-l\�)�"˯�^V�NbE ƈ?�Bh$��!/����rI#��ʇ=����*M\���(��&�.\t|*r��}�����U����6K�~�7X��Ȧ�Tt x�f��,�& �X��;F��J���A�)s���K�e�S��{ۅ
@h +��_��$
�iל^ �3B�<'� �*�_Λ�~���%�m�H�Y���f��i5�oDtkky�}�۱���A�R����}���n���=�
�`uH �T׍�+�L�3�Q]��>�����C"$��]�޸K��uz��;���W��ݼ�d�FVc��f�IǮ*_E��/��z�}*�L�Ͷã4}X�$o�%'}�z<�t��m��L'"�}���P�o��g�_��A�FNW��3M1�l>`���v$o���j��j�8Y�� ���jٶk5o��c�,I�FR�d��ϲ
8�|�s�,f9ބ�^��m�nL]��YL���W�w`ߪn�P^�敁Mm�0䍚��T?�ݝ������uA�����k���>>��WH�߃��bQ�Q�`=�݊k�<���]m�i�����Ӕ����,a҈
�3�*�"�?u�=�Q��'7�����IC+��V����͗�>�i�4�R)'�/=��5`��ѥ�G�,�7�ƺ�?�$J��swl�o�.9��Jh���3˘.x�N���Ͽ�����Ye�V�<ٮL��s��Y���VB>e;���z3l�b��������5�/
f��蝶�*��A�&�&0p�쫞�dđBWxV�&��U�` ����Bm��
p���6��y�&�-B�J,���s�G��z�����&
c�G>1���*7E���<�L�Jk}���l�u��
�.ȣ�>qtkh��8��u�������}�1�DD|�����-�)����R�6j����o~�~C�b�UJH�"�b`{��eB����Tгo���oU�9u�M��c���b_z�iP���%F���ۼ�~H��~����*� hb�3�6�^k���1A^�����JKo�sj �>/��`9�*�Dig��LĮ��w����.�����i;w����q?�,�ay��K����km��T�3��I�>�<���V�3숊p-�RIwF�A����@,�e�@����PKC�B廻$y��%k��;��a��M�Ѝ���EY.-E�QM��`��m-�\�U~�R�86�5o�1�Â��O�a�p�}H_B�����7rI����}�)��MV�.Ҭ�桁x����>��gZ���(�N������{D���Ǔ}���� 3ƁN����}�v�r��
���"�D	&�th�<L�(,� ����j�1�c���J% ����dXF���s&����n��!�������mj��D��U<(�]�ga�gLb_�����/�za4
|(\Ҳ�ns�Z�k��m6J�jC�r^�/�EB�F2���c@0h��m�/k}����{�K�{C�{κ!�n}��`�9@s��O��w�L�9���-Dy"��J����8��?�q�
����o��|Vא�n��o�}k�1�̞�x]s����r���}(P�Վ�Z�vh��������ࠎA�Ή	��Oa���tNS�p��.�gۨ�,/��v3mR�c�($4"Rl,�&4�{��X:,���*c�o.L���([�I��5��`�k�`ل����>Hh&���K���%��uٗ�in�"4�q�r�1٫&��h$�����l���ӜX�: �T�X�_kъ���I�']߃θ�P�e�����T��6�f���}]7!;K�XBR�O�Ri�8���,�3��h���1V�tVR��h�ٸe�%8�$ѧ�q/���,<CNz��HL�1zC�����תY�7L��t�t��RwD�A��QW�����F��ȐI��5!wI�[�j��R0�QY�8>5���)�5�b/���zPi���:z�:�TC���B��q{�'��|�g��i4���7�+f����!�7�J~u���KH���}����mc��<w��D�F��{JTP(Q�B�`���.q���X�5��y��W�C�l}he��Fu���=`�J=t��t�]Sn�ے�wm3Pe�1��0��8�SU��t�+��07�d��F~��9�<�~`x^ŧ�Bp��ң*�i>7�N�h��0�]��G�m�����R���p�6St1��͛�6NXYu�e�������2�B���ʍd�?D�Kj������V�	�)�p�w���?]ٜ:5TQ�6�Jv{�n�����7��8�yH�o2H���̺T �T�i��?��Q�!:1���7כ#�����q!�>���j�g4�+��=Љ�I"8�g��	oh'L�S�XS�'p�����L���>B��߀U�dP.nK'lӠ���(	,p�,��{�"�۩	�Dn
�I6@-�^�Kn�}�x�릷^�?]a{�Z�^�苜���^Q�Qi�LdԭŭQ�<�s����x��/�3�f�<.���[e>��˽"��{H��@��/d��@}P��"UoG���E�Pk��ͽ�������o��ɩ�1�@��JL���k����ޟB'�=�9�y8�9'	�Q�SQ�&���q���#ф0��O�
OFa�r8R��LB o�~�Ґ~�u%lQhWn('��#��aP���&Y��.&ا��N��#DcWlQ��e�K��o�.F?]\[�q.��O��E���]1)φm˺�|0��%�[�*��RU�����q�i��e��	��s�˽Kq�_o	����� tlL���;%�O]�Ѧ�#\�{��>��>y}B]�T/���д�R��{^�Pt�P�TO�@�n�-�����vl��h 7�	�_z$Y3��InҖ5�FlU�i�$uHuk�6&�����!�� �Ŀ�Fd���t2�,$��3i����%Gw�eC��~f>o�Vاpʨ�p�,�>�O��Y-�(��ڟ0yK��PtOv�,^w��۫� �y�S�~�yQ�r����\[1���Il�Aݦ_�B�%AZL��%�)Wq�jAEm\	�1;]�a�vj1����d<x	m|l�q RSQ�����>��O���� <X� �l��E�"׵�Ġ�e21���Ne��JB�)� �$�����e�b�)��1@�{H}bC+�݄V:�y������$�<�M��_�*t��4(��(<%�)�r�l#�n����lfx+��U�s��RY��@l�鉵YQπ��lu,F�DY�����W��.�V]�/U�/I��(b�j6�hs�B�!$�(�9e�(�pX���{(��r6��+t��#�r�Hjt�7�$�?����t��t�07d�U�̈́�]�R[i���6z�GZ	O�x����9����Q�t�J_�F�F�y��	}��X�U��|���_Ց}o�����g
;J��fv�!E�ڕ��AjzҒI���3O9O$���W�:�6�Ir�S,d_&$e��k�>�U��0��k}�<z
R/��l�N{��:Y���I3���Μ�H�I��py�a*ߤ��B/D
�F���OD�|��Z�nV�'���ژ%қi$���ډ4�:�2��j��璈C�@V�����K���Zj�cb��)ȴB������(��z�Eq�ݱ��];p	I�*��*�Y�炂�@���W��Mnq�^�z���rJB�M2f
��h��4:�Ԯ�*�N��5M'�F�~)�`YQ�v�S�����(�H�v���M�p�m���?����\􆇫�{����{htU��9<�F��m7@k������{�%N�aziB���SW` 'VV�A���bW^�������������\�L85���e���J�AF/��u۳AX��ڒ�h}g}���4��Y���i����]�X8�>���7Bͼ2xo��@~-��RQ������8d��.j�����'�")����˒�~��+��V|�4��!w_�HX��]�:,@lg����\��! |�'��LώS�[�2�=C~F�H
zY�7�1q��$���A�) f���r��eQ�Kɹ�j�FK]�f:#�>�@�_ܙ��;���+ȼ׋n�p�s��q>O��t���E�U�0]����Nժ+��{?�?i&������������e�d\����0���+��W���_���D#�E@�*Lk$X%z?|�{C�9V��9 \��Uذ���m�M֞;�	KhJ���z#�^�Uը�U��[�rVi@�8o��+���좕|���"������2�L�F�b� ��y�% ��r�)�,u�����z&C8�܋���|T�G����>W,�Y� ������BMF�F,�30LO��}�?�Ǖ���R/Z��X�*�3?"�/ �E8���6��x��3��'Q`1<~�y�0��R�v���(���g�=6�W}o����a�i������[���G���c�/���\�r!t�7�-���q���HH�f@'���#�?؞o�$�pn�_�x*���>���4%�h��p�����UP��S���N�:ѡ��4c2��Y��.Y���	Z�ڀxjO��yn��kYw[r@:#+��e;�?Ҟ��30�3�q���1Y�(+�uʂ�VU{�y7("3m�G��z�a�b�ҽ�4<�
|kc�{�<�N-(!�Q:��J��;gS՝��s>��[H@�0OM����ȃ=0jeN��	����@��6�Ne߿�,zBS�Ks@t���k|V�x�%�}��Cѓ>�edD}�Z�WK�ua8%���ă8!*�%pF��TV��Dv��1�sBb�]w�����j�76��}Q����0��U4 �e�+f��|�
�fkj�o�� U�ز�`��ϙ#�&�i��-	��_r7�6�D�J���w�5L���k�AzG�N�E��UjQq&4Q�;oX9�<���
�MQ�/6��9<r�qG��触]JK_1��hj.3j.$�P懇������we��E����B�+���a�������/)4�5q��q��14�)��\q݋�zO	V���Z:���a��S����)线X6WϬO�V�}>��@Z@�Q �gBB���!H #:ZI��[#׈��-��� ��6�� �����8�I�t8�$�s�^�%yAtɦ_Ga68��fz����E{��x];�3e�>-�,��O�b8�}�)P���ْ]*�S�9Zam$� �f���X♔�<&���(Ii�`�#jq��`v<�a �$�C�hv�Q:6��{��ѰI��$`��ݪ���v3s�����,�ig��HZ�D��0�.d�N*�=��ρH���`�&���{�z�A�4����X/p3�����k���䌏_(��J�Ʋ�
,;z����X�k
��r,�H�'n�(�J���08�,�&Qli^�����K*�o��-��-~�㉥��moi�W�U0�M�kp�d��=4��Ȟ���^o�]�ԡ�|,�< �~���.��v����l�������=��c�l�Xߔ�7ٰ��Ӆ:D��Z)p�d/�?"����m�����?]����I:��o~�.��V퓮,k˫�J�KId5�M��X\?ɬ� fb����-��u�0�A,��#�{h+�[�F�8��U� z�<g��e��ǋ>�Kwr}�(�u�Ma��tb9
�@��c�������N���̂�����N�x�z:i~�9�N�O�
S_��>� ܍vAw�3�Գ���ܾ��KM���@���`|~�{���qo�h���C��sDh4cW�y8T$��g�#�\M����`xjߕ\D���0�Ioc�;Fs���'�`�7��gR�>'ykm�h���_y�i����I� �;4�T�"6�f��0!y����V�

1�;iąV.,�n������)���j�5�c�x��p��iŗ�<$��)3�.�֬|ġe�Eك	�&_��a������?����p�R���̖n�&�EOZ�}�R3�+wѴ�\�ϟL�p
�?鯼a5���{x/P%�ʨPR�p��O�m.���g���1[��(bH6P8�x�f�+��v��E�U/zV+�(�g`
B�C=8]1~w�0�8������ʇ@�o��4�V�������Z�hX�A�?���1QA��)5kʕA�N��*LW�
s�+���Qz@���M@��U���l"b)�
����'s˘'�n��AX�Vkf�1�횞��0�C�O� V�S�{���U�.� .�~yH�]E�,v�v���6f	$�H������wR�H��\�>V��J��q��ērW ��ʊ�w�n��3��� Qd'�g�Y+߬�,OF�
O��7[ ^YRj����IH�9�#u6$��FX/�<c�;��~�3ė�x�P��~�8ռc��^��r�;"��Pɲ�eU�D��r8�e�,���Ə�%<+�1����Wy����zW�ze�Ǥ�1�dV�����l��Sx��K`���@<�{�'���φ����^z���T]�5�H�0����K��X�J#`3����3�u\)��TH��E�A�Hn�.��v��+�����ŋ~�[ڀl�6=�,�}ڔ��.7��;~�Dچl���h�M�-�l&\;�x�g�H���Eu_PP��JqE˃L�$���K�� +f�.�'[���J�)7�u��?�R����%+^�%+{t�+��F�iN I<�����"@�|u'�I���P:�p!?���*��9v�د��Q�&ԫZ<q!+.*�t� I�M���3ʤ濇�'��+�.'>ڶ-��c8���B�gP�~�.X�S��I[t´f�	��w��}���T"�f��\�B��vZ������2��4��ݩ�yZ�(5xy�x5�z�Q{��B��",
������`�� �m$�D���BQ�}�W>���b���������6sW���D�8��/�E��I��->�$`�p�"YO^1��0�P�>��w*���ޔ�O��f� �*1h8 ߢR��V �Y�k�Q�Ls�Ѻ����\��b>��U�Z#�u5Y���q�������w���`� ț΋8Z��t#�p��R�,y�
lm**�(��j>�?*�3G��o�����=-'S8��Y�o|tt $���9����& �|���g�u�Ij�A��$#b�;���]g�_�g���'�u���Ls��_y@X.�I�e�`gc(��}��J���;�v��I��cć���a���JQ���&oݴ��IH����
za�M��J��k҂jB�gzU��\���g��/w�6����<�f���Uȥ���3�p�*�;�ⶵW����l}�{��WZ��"]q6��t��6x
��Tu�\J��x�
�j�!����	�S����<�nbN��w~4i���PM�L��TS��?��+�������-��$�I�]j\�'bg�h5\��b�Wn�I,�<��4Q��EU�Mx�
�3p�Ģ{i#{]��}��_���-6�U�;��.ԗM���*�����P]=��ZJ<�~y�\c3�̚�v#��6�%^�� R�	���8?���Ɂ�*�r�����`�_z*�V�x��\��BT_��{fғ�EӋZ��ti��S�q�H�C�a-cF���6S�&�C��~���r1B���T�$�	'��P?/5-ZO�|&��`���� ��#��x*h�O�<�PZ=�F�? �"0؆D��8�������f��?~�(���T�@��k���'bA�$`�Kg��2�I����5zK:�~k����`�-�R0��e3�SU�T�x�+x ,�H{����N����_U��d�ִK�;U�1��ws��* �&�[�\QDh�z��4��zY/Q4��7��k�X����9.j�����n�3w�\���{�qLYbS�H�Ý[�v^��� ��B�w�M1���>�ʳ���<�W�:=��{��I'��?�}ˁY��=R��H1|l3�(�^�L���Xl�-���N�]-�н����4%�ӟ���cj��:
M��*� �"�2���)��«Ys��J�XT&���� s�/u�U���R��1�~Ar��uB�:������(��Ld�r:���xd�C�d�y8
���r&�~U(�4��2o	��>y� ��){ke{!�ɑk���jk��(���h�II�EWABMc7R��>\	D<�K�b���5nFe'=e���?�dE<2(4���C곦����$�ֵ���}U�uDp���_Z�$�)�L]����^u8�4R$fe�g�W*����=��=����W��"j0J`�薎����R>0�T��^��m��B	�X:r�=eOa���U@9�/c]�U�����f��K`�@v�$&\�j1��� �*���D��T0Mb1��5{�)�n��]D1 ��fJ *{��4�  w#Q���X/c�Y�'�G�*�f�h(Yn��ڤ�N�?N���h�I���,�Zv&����q�>�9:���]N6m�f4U�؟b��Eɷ��6!�Wt��~��6�����׆���v^��5]��x�2��?N�֏�{�:�(�}�<��_�h_�QXFz��}����4�6Ϋ=����e�mY�x.�$/'�R�͍f1��y�},V`�z� ����p�H�
�#�����hΨ#�.���,�Ŕd�«1�M(���߂���'%��C��Z��a����Ȯ�����g�rbn�@��<��toq�sU]dxe��Q��v����@���b��X�4���is<@��+`"	���5�M��{�Y�~�Ǟ
�u�`�_ݽ��j�~��\��,R�f�:�� �:}����;O�E��ԥdG�6���O
��ڀ�n^����D�1���R����}
p
f��`TlyJ71v7�'%q����Eȕ)^�Ⳛ_���$��0��6�� ���^SP��iw��5ۅU�hO��]�E��
S��0hv[�d؃V�d����:NѻJያH���H@����&�3�D^��令f���~y�!�P�j�bwbN��
���X�j=��}�V�Z>MVY8�v����1��q�c���ٚB�ŧ�p��"��-_�+ؐq��ٝ�!^\>��z�U��Bx��Y�y�7���+&�	�X��m&|���[���]�A^��!|*H���_���������[4�N2!2�[�>8ʨ��
��J�Qɯ�;u)�x�ls��6�0z�Ad����7�I�N�vsܶk��~�b�R�H2
�0a&{��K�Ľ��7&2��&v��F[���i��������1];�>A�{��k9"����]a�ޡ��m���8f����'��_��g��@�sloy#��p�'�������C�\��IyX�+�Ȧ�\nq�I���N��!��[P᝝�X	��$C���:�����t������5��{��h���&M��X⽝ ��zyU�<$-%� ��`��;-7�/�;6T�ʚo���9�dk�� f���T?ҪǽQ}��wB����G�dl 3a2>��~R�ڌ��5��bc5(S�%�9Y l�!R��-N:<^ Ԇ���o���oD��&��ci�qg���<�l�r�fEB1D�4�a�T޿��]n�3,��{�;�i���%�ibߛּ�Zm�u�֫ ���q�zZ�+;I�F����@(��IP���4,���W6��Bm�p?Rf�R��!Х�'�0&����%���7�e)kX�z��0�DfPE��8`X�*Ձ���@�.�0��>��f�DaAe8� F��	�(l��$�"D8�g��V"B�N(��ŘZDkr��{�ן�,_�f�� @��Y[ċ wP��5��=��� �w3�֊n��ʸ;�!� �I2es�r�icE#L��r)�m^:=M������w�!�r��ٿ�KҌF�O�Y��Hʒ���DP�H���HqH�}]2��5R}�r,�*H�e����9�8���ښRڏƚ�j�fy��;j����M��e�Z�T/���$��Y���*v50n��}�'����Ң�HA�!}�b+���8�2\ѧgy�����3Ǐ�hk�|}��K�Oq��=�s�]c)�~�lO@����l�e~F��W�8��*d�+�����^�y����"����@��1-���-����4���;΄ǽ_C���A3ӷ�du�ָLa���ߦ$$S׈��mUҿ �I�1$R��n{���ܥKJĤo��o��4�"0�1.?z�)�S���m�Ƭ���7���:TbS��$ҭ��+�0-��k��k$\��p�6ۄ��.L&|k4�N(6�Ժ��ӟ9푟Uoj!���e���prn�IG���2#6uIF�_F��y� 5�,+B}C�^R��a�[O�u�2QV���(lN&�Bz�P�]��M=ZuVX[��ۤv�"h\�kJH���	^Ҩ��͙b:��4V7����ڀ�qw��t�>���B�-k�D`�a`�p��aX�}��EB�}r���a$�J=�|g<A�
���΅�5�c��"��\"A?��&�HN2���pHiyF�X>W�CT!����E�.0��oLJ�m�WW0E�IHA�?�T�ǅ��cYt��W9(�9�������8�WT��ESO�B/��a��h�l�κ��)y���}�ؑ����k/[C������y@�����;Q�l��SO*��7?�t�9N�S��1
n�G��CT�C��9n���;O���~��ߟ�|��T�qH%GĻ�E{�
8�k{}1�|�B�\�T��#ɛ���yO/��� GF*U�cU2��0Z��z�en�n�@����jg{���o��+�-�6�����e�2�X]�&�m�ŷd�m��� ?�0ơ�þ��~J�p����Hag��^k�� -��������IL��S�k��E}@i8�a��2��
#GVr���*:��Y��DE������ȡ{��ϥ��"��Z5"�P�^�u�^�XӀ[��P� ���mA�.cW)�1cAtƟN0|�d�25j�Rvn�y�L-z>@����4��K��:�MXu/$٭��5�i��V��G�6-ڊ�WCmvL���
N����TA�z�����F�cqf��K,(У�Oת��O���T��u+�@X����ϝna �C�<�P9Np�>!\�X��h��B�*;��E��Y�����\J{�j������ħ��`M=�a��:�ߛ� �*PDوN�V�]��t�pCMGk�E���N��"ͷ-q�ct��hzI�*�uDkε�J��ٹ�x�zhO��"��?�������;�aՍ�P���ֹ���O�����K�ly���{�r D.X��G�����/˯�Ǫ��S������c;���pqn�> �&Kcf��3<]*���Q�K��{Q>��"ů�I���z�?[F�j����]�<���,�$*c+U����@4�q�1��0?���N�d0?��8(/����4ڜ����9HA�L�W~�oa{�cPR<N��=���;��L��Nq�6�L^!�bd겗	��̞t3��\�3�k��5hg?w�#v4ݍRR z&�����D����M+io �/`�Զ2��~d���D�'X�� 5�i�ǥ9��R�@��o҂2�r��zI�M�jB�ar�^��|�>+mT��#g���]ɔ�0�����!H��0�dR�J�o�L�c����V�۶���=�Qř��$6+�JQ����7�#a:mԏ�o�+��a�*�N&�'�T���gA)��dhg ��E���דB[��X|�7��i6���Ӓ#�A�K}��۬	^�z
Z�wwMa����
����:A��\-�(蜇��s�͹.�g������T)��6��+�(
�`�>�`��t����v��0cF>���������_=�-뗉񄴊ʊ0�A��S�����@��T@��'�-��f��uaNh���r���N�'ws��+~��T�W�a%�yj���3�]�f���tM��Lǩ��&�h��\�� W�֯D� �aB@�Z����h�6&�|���b �	2ŹH��c!��X��xH�{�.i ��Á\X6u�B���9%_��9OxQ��[�1[:e�I�����@ %�jp �?���|p����t�x�7�b>��X9p�(�}��DT��r��=8j�Q+4s�_���b@95�D��^�_�t��A�;�Bb`�ڠ���n��}4��������2/�\�>Hd������I�sn�ڽ#��D�Ds��E�/fXa@�$�]�g�8G�e ���a��u4Z�K���uG|��8u\7��zgs'd�� \ͅdu�����JA�������>R)I���'OT@��]㻓7-��I�j0ƍU��3��Y?k<i��2<(�%G9F�s��7�nh<:���ZMI�E��,Q(�F[���>28q*�|H��\q6h$�2����I�pEm���`�*{��*%ʪ��#�����}��]'�KNV hڟߖ�n�;3��Op���1��Mm#ǜjLrrǻ�Ǥw���N�\W��- ��F#f+3�}�7��lA�i2>3�V�V���/���l��$���$I�m�<=��{��e�Ǉ^�i ]�4�P��W�w��.;0c[V�Dt�΀�{� 5���ؔ �1��u5{�LMl�E>�y����d�7��̑��p��:�<�暱�N���Clc�O�<�}4���K[��O�gS;��d��#�;{æ�2�;������O�LP1ɳ�Y�����1���Z�Nt��$Z����Kw��~��a�g�G�R%]�m�*��P���D$$rY��;&F~��e��2+���-��ɘ=F��sϛ�O���NxK�>q��>��h!o̒��Su�V��#�!�4���Pו0���I�2�)a�y�9*�W�j�K3�*îiA'�֦{�i�1S�J,��\�{+3*s���C$��+�ٖ�Z������fUf��~��K��������A���/^��F_�u��a��u�\ �٬y�Čm�J�dD[g�?�,�C�<����������d^����KC��6�?���E/x���?�u�[敁�Ͼ��������֨ڠ�����1諚K������5�c@�ۉ$9�jT���zH\��>b^�n��X�$p"$�R��
٧Rh�o-��y$~���#�1��0×�h�9�H�@Мp�I���-��\#K���T,�k��%�1��	(�G��:�s�tl/�P1}'��p"ܡ"�|�0?�j&����s����{�q~�ݘ���ӯC�ԍ���R�/��<.�*�-�
W���j�����0�ކ{�t "N����#�1{�����9V�����;v,�}�}? �5�1ߣ&�j4���mL�-=K�^�aI���ƺ&���OQ_��{s�F�3��Eܿ�)� *��X
Wd.|0r#Χ!�m�Uٲ������n��~���x�ywV��k���,cl�S���i��h��]1���;ĠN�3v˚���T�Nb���q�)px����`Wb��L(Fw���*J��As���q��jy�oy(s����hCI��B��ZU�\�of�^լѣ{=$�+�	l�-�$�2�1N��ڔ�z
U�6�[i�݅���|&�l���"�G�����AT�[��t���&a�� n��C��D��0/�H�V�� s�`�'���/r>�%~;�b���62j˫�o��-����*�4�@Up��I2;+A��,�'7�&�;�=nV @�w�ɗ�:<��%���������Q�a�"�t�&����yAF��]�	#%g�]����ji�0�b��y�y��k:�N)�]����;������Z����2�����:b,��`v�����>�[����ÊW�!�A�_U6Xױ�<�����	2�ă��T�#���S���0�=5�y;������/�ދ.�~2h݂���{ ���3�)����,�z��������� GaQ�U	F&�|DH��ݍڈ��\�$���_�QK_���ڮ�d��p�@�hn:b�[*%���z��=:�]�'���2���92I!�Bѹ�ř�<߷ҌA���V���Sc� ��~o��]�Q��d�jئ�&Z���A�H���2�uK)����C�/Xf�ڄq����MӃ�t	�bK{�<vn�qvsp��]q=�����6_&�s�T&͛Y?нe�Y�ϑ464w�~-���DB�(������=`�/�AI����P61�f�M8������ �4D�l��S�W�F�"������{J�	Ec���^�� L�� �6MD�������|K��-��$���_d�c��F��*��`�Iڟ\d՞�d��h�5Y帻~�������5Q���!�0fCc���N�э?Äω7�aL�9?�RC�(��I!k��`��)�N�A��?/�F����0d���^��6Bm��S\�G1w�d蚟����łE�I�ȤM1�CG��v�� �
�Z�1KE��ࡒ��[�z��ܚ&8\���^�R{(��I�s�n�Q� ��yL�>�������x�i���A��*�|��� �u<?[�U�p����yơ��W��HE�S�����|^��#��g���
wْB�,ؖ0��{W�s��:��%�����t��b�Ss*��E���;��8 R�G5���ʔ���>:Q��5�U�/����1O,/X#�,�/���peR�}�5^�u֝S�Usn�v�ҍ�fg� �E '����E���$B=��L�7O5����]+}��g���������4�3�NVFv��(���K�¹�"�yf e�zAk�Ԙ�g	�����U����h%�c��6�(�&���g�ϟ'��V����;���s�\�7),Wl�w�u�Z�	`=Q����h�I���k�����=�~�2f�T8�bqL�����<�������o�J�~���£Zs���!Qj��!u*3U�'��Ãx�DI����K]F+A��$�6W��T ���Q
3y�3���|����v>���F��yf���;Ou�y��bC(�j!d�84#ICo��G���F�e@?E�Y[Ƚ�������~"G5��h��x��9���ߝ D�|)N�o>�T��P�	���^�F�h$p�)�$v�]n��@ycB�!j{`u;��H�)�A1�3��C�f��T9�|��[1Pt�7%�Y�v� ԝ�(>	������;C�ը��l�E�S�4�?m��ؖjB��� �|����7���l�Q�6���G�4ᡥBf���9�H`F���� E�Q-J$h3�-s՝�"7���0���+�R�=��W�dڸv���5��J���Z�L��.:�'�pp,�v�׭������L�dYw�R�. ��G�{�-�S���K��}�C��}ӆ�ЗT�p ��D՟.(����(�+j=��s���EFh���
,J���U�Z�b��޺�0����"%w�s$c�p$�Q7���tyIȫ�U�͡ҷ2�Fsowg�!Y�A�����W��`y@�o�ˣ�H��]@��	�J��V7�D����w��C��j�468����5�a��S0��e[1虯��=I�89ٙԄ��&���遨�jc2e�*oM��(f� A
�x�� ��vDG�}��QF��Z�:����c�02q|�Nk����z�����mڢ��o)s�B��>?�^k��0R�x�>`��@V�78��ĀR�_|&	�%����K�����=d-�����Lf�rP��Q˶.�����G�Z�Xp:P��[�����P�5o�6��t��̤�#?���+�èe{�2�SYׄ���-T��3�N��n�L����|�>�:����P��'kZ�8�P�Z�wyl�)��ȉh-*h2t��,[8d��ʓ�tc�ŬT£�1�w�S-ũ��z=��.�s�ʾ�%����^�4�oQ��>��|6;����k4<��\�|a:�02�]�bb�7�\wJ,�o�u��l��Ǥ�)4Qoôm�z!��?����Q��a_�����|5�溼1�
�6���[ �D=/�$�{��jr���\�b�Z�,�P{x"�x���8�/I{Kc�m�=�?Hk��z/W�=�]ڋ�f�R�d�K%7��}�N�� �ޘq�W*��qS��\~D#h��"���rGJ��e�򵚲\��S�.9�ۓܩ#�<� 4���i�D��ݝ�pSj�66��ؠRZ﭅U��ܗ�z���+v���C��u�@�fK���u�.'�~��4��ED�Za���	+����2,ճȱԺ�<�|� VQ64�=�����4�&���ilʶ����G�ƢKB��(�8_��$#�����ՍD���-g����"Y;��t�� �nֳ���{�Y���������	c{��p�N�|�(L�|t���$�+}�Qv��Ȋ����ʼ�l�,;>��~|�t#R�x�`ˉs��!�;:E������ʜSr����O��Y`vtTI�4E|y�_�/���w����6r�?1��I1��VR���|؄#�[��"l�/�
��oF�����r" �G������{}'�`Nˋ�{v���^��LKB���)�T���E������|V�T1�����[x����Fo�<Ə|(h�/J����f�e�H�v,��Rt6AĖ�6�1*�E��{�u"F@@c����~�Y1)�C���7�@�C;�,�Z9Rģ����� !�/B��LPf���X��P����O��F��"�ܢ	TI�����w�8�5(ѦW��;�aw�%m�i�]<���89 �)���S֯�f���65�J�ݗܶ�*i#��;7�M*���ax��}t�)�Be�L0T	�]	��:av�*`�pY�ްx�»�Kڂj���*%�`���Q<#�ܨc�D�&�7��8������_M\��
.>TQw���[��i`/�"lK�O���w��3�dʦZNa\�^�^�~�-��&���?^���t-Ɨ�!��yÿ�"����,�S���T�O6Շ�0�2X}�(X<1���GY?�H��p��0�O��OW���K��>&�Fq2�ܔ)!���{>�����)8ʜ
F�@"_�<{3���:���psW� �{��75=�e���#�&)�i�A��L��"��\�n��>�en^��O.��)�"��`��Gd��30;7%�F�)Վ��-˙�Ҩ�Z���Td9�W�^����������#���ն�������C�He�rƠƇp�9tUƋ!���4��V.\��`GB�)ƞ��t�2����z��'���1�،W�0������İ��1.�^�뾾��F: x��
��{�sۓ��`�Sn��bn�[��׊7ۥ��3̧1k�Q|�����Kdp{[7�J�gO;�R�S��L����_ӄ=��������R����%�M��e����u�a��xFo��d�%uq�G���	��t�M�����$Y��%����G��5$^�ڛ�k�)�3R����U�*T1�����l���L� ��@�
kr9��օ��;��m"�o'QuN+&�R;Nc����%�q?�i�/����a�ZO�s�������$}s�l�<�%��:�`�g��̍W�j�Cۂ�8˶g}�JiY����������� �D�4 ݍxY��&=�������
i׾� �ɇ��_���m�ō���έ"�����J��8K�-$>x�����FQ^θm�fZ�ł�E�l��'� �'[٣����B�������� ���y��4[��v���]J����F�f]�&t�a?*�:��̺�a��n��Mv1���k�m��2d�
�=٭�{��"
fvZ�c���Gr�bh컫�<r�����!�R\0T �MŮ���[������%��
���r~�S窺���,Wܿ�m�q�҄��8�&f5�}�-Xpd�;�na�0�~�Q3���v��݋C����4Cvq�|��Z�O8Ud���D�Q�>�%3�U22��w�+�,�5i�h7�H��[��,�.#�}f2ړs�Pu9�!�*�5��GHm���%~ۗ�uD�:�,6�(�%=�=�I0���XO7p����;�0��fq`�ƣpH�tY�,��2H���ǃv&Y������PK"kI�p�T�4J����Q�˞��]�40�}
ӿ�؃L���s0���S� �������VxP�����{�H��E^��e@��J�{ ]~9�XY�x���-�d���ڲ*�qf�ĳ��+(V�:�,x���\�s=K��Z�	ذ��p��z��fi�)>%p�5���ę�jU���<m�6�݁��V%z-�n�5|��7�O45;����S�
�� Suss��DTv9I{��p��?A�!x���/�Ey�4��G�i9�N~�r��
���#���xib�"�z���v��Wᴬ$�Azq_2zФ�wԍKN����t���ʨQ�uu��r��+�����Q|�dI|�^����+�5�_Ż(��VLj�,��؍��І���i^�	��{݉d���Q*������8l��^�
13I�1�1�aC�7�^mM��\\P*���=��b�$����wNAӡ�P�-�xȓK�碔�.���S��v��D�g�WH�L�͒S��i���Vyy�:ߧ�h�͉��� �vf��@�v����[�;�J�FXJ�P��凗�U�QJr���H,[\�%�nf�lc�Ԕ5�y�24$��'�$�:'Xߛ,�7��]"�-�����d��"�C�pe 5�U��\C���S��M�=�#���� �Ʃ�	b���Kc��h�a�*)���ɶ<���Z8�s�!�_�[5��I3Ъ�D�賟'PN��7��1h�E�Ҵ�i�E��4�u�� �6:��$\��QŕM��O.,<H����t@�ߣmҧ��[��5�o�e������(١�����[<��j������y�+S5s�X�3�TJ̝���A�&tL�L��������t�hge��R�U�i�kT��yuY̲t��q;�ܟ����z��K�sC���?rp�qE�ԥ���l��s�zsd�\�Bx<��0�C^�W��U%�T���� �w�RP+��H�[�ǨqO��́�M� �-�PQ�ms��
���$E�J}� �.�V`����Շ�C!��R��}���������k���8��㮭�W��l��+=�;�~���P+F�FW�ۣ@��"���e�`5�Stz�d�T9��Y���_�7?8�[�eoz�%QQR����䰎Ox�xF� %��NzI�(�l�[A��Y=����ϲ��;+*�̺������-��	3d�ֈn?�1��i5���O�߷��vIt�98�/,6��)\��@-2�('$#�Ǳ�?�Q���cgܙ\���7m6��O�T�6�z�5�hz=�V��<�<��������X梙AS����}XG������^�ue#�&�d��Y�+�m��T(�!$�>֣G�~�I�W�8�5mL��!=����$��(v���;Z�\s�ꢒ�(��N�{�!"�x;�ۯ>`ߘx�!�#muG��u�*H�N����TB�0$��6=
i���Wc�E7��KC�_����`Z�Ls�CPY�e����}ՙz����*+8;R��ڃ(���@�����{R3�f��d�l!6��\��g˂�k�9�k�����/D�aF����q��M�B���h R����S2�����$p���!��W��{�
��� �t4Fb�Ė��[F��ǅu�<��\G���I�LÓ��u�UC?Iq�t��P���YD�Q� �����H*~X?���(��}v<m?�	����^66�oV�����Vvb�,0�W��w hbg��<���g�g��C����ؾ����;�"z�6����ݎ��K�OӫiyL�q�)���r]o�	�s�QK�r�Vk��4�u׬24��_U�ǐ���3�i�B�B�	*m���ZNfI�x ��,�Z�v�p�=-�V
��]�a�_+���Ȥ֒�8�:��8��Mw�֞M�f  ��^c�5��H}���l+���(u
R�
S^2"R�\���K'c�l��f�WZykf"�ݰ�t�~����B��o�%<�u�x1�'�]����$Q������%��f�$׽�9����[[��ve������'�f
�K�/��j�R��1����Hk�3����FV�d<kd�B��m:�#���i{?h@c#�SX�����[��������"V��1�C�Ԧú8�K�g��j��Ai;!<�b��C���^�	�����φ�$so�bvϟ����c����x��*��{�5�k�eU����0=X4T)��D��j̏��k��6V\J�\+X���f� �ʳ����u$�h쩌AB����w����v�����d:���y /�@C{V.��:�T����8�����ϳ��Ofё��xgt���J9; ^�ß��H����_���n��	�S��;�`	z��sD�\��OP�S�D�@d�WMȺ8�Z[ёW���}<;�Ti}�.�P��*��/������[~t�v��4-�v���D������<�z�H#t�����ڱ�i*P��H��̃��q��~��~��5ʳ �"��HX>��e���������������4a�V��h�A�wѹ�K{+-q��\��}���2_�t��O*��V��9:��ౌ*�'�,�t]K@[�O<�v�薹�yv=���=�3��4�t�I�Z'�/��ӕ�Xa����.Tn�/�����[Q䎮:9�׍�{Ġ(�}���z=�=�����Ew~&R��"پ8~ز���\sU�c�piAB��L!�
*S*�Ư�z���CcZ����첞�g?⸾�����2�)g�D��fr3���3��P�!R�����Xs0��渵��)P'�U�p���D�����$��Je`u%��J�ܶ���5�����h�FW-�'�,��z��x���W���"�36�)6H�
h�h��*ۘ�x=.U��t��\,ˏ�ل.a�\���zҋ�R�8[O�^���8	$����b뱢���"��p�QR�����'���.���(���A	��Ѕ���ܐZ�>c#��N�����G�%�O�--9�C<F��φ�ܴ��d���ށ6t����QdU�*�Z�T��	x����}Λ	�Faj��]���+��$�Js�]�Ԇb7Mߟ�6�~Y�����[U R>O�8c���n]I���	�xq�����;;�S���Q��%~���
��b[����Ԭl�i��?H��/�/<+��0����͎[�����Y^��I�2ݍ���7;�	2���B��P��9��3��`\��i�8�9f�bInc��
�M��H�����g���V@�μ�y`����0.���d��eKNtGd��~�`QQ�[��a�*C"SK��N�cPy�mmI�ώ4q3u�Z��HH�+��t(D��M$0N+>�ЊLi�������H�sW�E�~����%4d��*铗�H4;������RX�j�����%{��\KU��5��������볭�ħk������[��2m󐣴.d6^���4l���S�}�='�U� �45�1�;�Epl�6��)�=c0�����ۃI�X��{z_ /�HN�	�-�f(�~����%���g��s�L���"���n�v���v����r�7��d���}����q�"�L�- ���8n8E�$<@I$<�c�A(��N���S�>m�0ު���\���Wn���N�~�Dӂ�sČ�`�aͽ�J t��s���8���!:� on���v��z�%z���Ҧ���k���T�C�"���>�����Z���S����}�D����,X������������	�9W�v�KyF=��������<"��8n�C��~k&�sR�^Ñ��Z��Kp��%����c;k�0��N�:RA�e�U�/Q	s������&�n��Ñ��0����Y⿮�[�W4�7����1��r.������`�i���}� �^����++�LΖ���F�'C�j�V*���m�O�)�ʯ�QA�}���E��G��R�S���p7�t��K�7�]q\�p�����?�k�a|�-�
q�l�D2��.[�+�
��Dt(=Z OUL=��� ��6|:��\��ҢEU^;Y�H�mQ�i6�Qp�]	��5�ac`�95�⌥�s�H�l���#���'�k�v
�Q�;>B�����U,�Z�q�h�����6����?3��yi���e�� �p7��Q�z.XH����ݖSWңuH��*>-X^ʨLvMo�N�����p2#�?s^l��]L�Hބ��	�ٝ��se	�-9�M��
����r_C��z��7V&�`r���v�Rڏ�6�@tR��M��#Oȇ�5m�8cn\���zD�J�,��9u@�r������u|,�J2û�!���U�I�]|��̓b�h�H�y%��]�y����&K��>r�DԪ���uV���O�����}��aAa�׎���8�>R}"+!hzu���=,΋�_rRG!C)�Y��E�ʤ�R�nK:5��1��U�J�MG�Z$rA�=�7��.��Z%q�O�g\	�v�X�X�%��dR^a&���O�ҍ]Fk���������^]{����w���ik`=�&�o8w���Fz��'�e���u�~�m��n������'��Q���l�鷋�)�-��߿�&�Q�\�s1��G�R�X�������I��t����䳤�X��}=�/�G6��Ž���(d�Hf�g�wYT��!�h��o-Z�@u�3u��$L����aaW���yj�5b@���wr#�i���R�+�T�T@)Z������)������&�lH�~W��.�J��g���L�%�n�&V�l�BY��&��:RP�ʊI�X��%�t�#X���7�@ƫ�h��f�Ԛ����I�<�Jo�B�X��Q�B5�	S�JT+��sA�� �u-�Z�R��\N8�E�m���U(՛��l�5��.�#9��i#��oD�{X⥜bċ\���;�C�б�+H;o��������O(����ܙ�E
*S I&P�w�7r�;Qj��t2[l_y2q�Ц����ъע�
S� ��W�=�5 �\�n`ک�Vi�(�H_x:T#es�T�)�'_��%#%M�5�It<:}����ib�Df����L=��]O�
m�}Okm �>=��ɻ�}LMʺ d>m���ji��}%$nH/3��_T���3|c��YwSDM���{]�)��/b4����R0;,�z�Ғ���i�L��E��kFg:�T2qw�^�^��Ob�E7��
X-E��Pgu�EA���b\��i�,��ʂ����ԅ�9��OnZ�4
�H�~ԯ����%�8�l)�'��?#h�G~&�6P�-īƆ����<KrƔ��O�pT �6�3%��8|[����dBqs}��Q�)�g�ğ�9H�z{�x+��9WФ��4���8�ohLg���N�r�.�:�E	7^(�o�B���zSD�is�[�tnΩ�d�Ʀ{F I�o#o7Tr�T�FU�	Q�;��aMӑ�9ˀ�$�9�"�_	m��$�1Q�Rc��%K���e���,�fG���T`xY�K���[!�+�6_��x��m�Q%;;H�ά*)�������)���J�Z��P���Q�[��b�RQ:+����YJi��!t>,������A�:�h��O��|T~��l�*��sL��M1)��Z�<�Va��*�-9�)����؎+p�RPm9I��7�X����ĥ��S{/nw%ÍC���I c;������럋�͆Q����E��2��:�@Y��TԲ8/�9j%q�Jy�E[�F^	���"���Z�B������2���2�'ˉ�,_$d��kq��l<�y,��eݗ��'�G�5�P���Մ��@��_.� f%���E��◂��Lé�d�I���s��
n���5�%
�&��:d���L&ܯ.�l�fU��G���j!�\�w��/v�F��r1��ӗZL�����~|,Я�4�N����,�����e:{Oc���Ϡ\#X�U׶2��W�L��MG%���a���zo1��"��N2���֜���˩�k�)����vi����o�z���o~U��x!72�v�I�e����XG+i'bw�X]O�����b-�����#0�k��@wfϽ%?�+�
�	-���c�����uD5*R92��l�3�mJ\l-h҃(8d���ā_�� �d���g��[��;�m:8~��k�> ��p�0�̘eB ~�T�Gj"��Bd��jNcN����R����Z3R�a�S���lS1���M@7�h�\A�	t�6���k��Û�^׉;?��U1+��w�!;r����8S������9�B�$ЏzUJ�����L�G�<�@|	���\n;v-qk3f�όL���\��C����-�Ș����@�M[�}�e4g��#s" �NKjV�yx_�UpSj��$�zx�@��P�-��c1j:�pK�?�n���ﮉvyt0�'�%��`"t 	 ��eFR�7E��z���1N[��v҉��9#
WY�鰿�w,@ OdR_B�*���	� �\}�����G;�F�>K�*ަ�_-���N2��x�Q�y���kc����YA�':%*���R����z{�]u�+��|_?ɤ$U�lYanlZ�`�k?=��A��S���	t���F��N`�@Z{���K�=Mt��HoW�>6"g#��N�T���j�jJ/�����CϏ�uG%S����Y�A�)W���/k�e<Qf[�
�D��L�����W�In�1�b�6�@g,��w�y���\)�R��S�I%?D�B�i4�;��T�������%xL��T�����ڀ�c��;�c嫟<��]X�Oq��k�չ�p����&�I��� /9LU���.����.�t� ��d���y����$g뺇�ܳ�a9yX�Պ\��sb����q&a=�� �z��b����\x��ܹ ����<#r�����8����|�|k����	���_)0��ا�Sc�)��[T�Э�0���㕇��P<Q	�7�ę�"�*=��D�E�����n��N��:|�J�w��Jք��ي ����*�_b��!�N(��|��'��$�=o��E Uŋ���[��v6�c=��P����q�҅9��;�)���kA�Y�R�`R�z_0\�XkS����0�km3�!-�q��10��<�E\Zu�5�s3�+�B�W	&cꝗ���ք#�Xo�g�/���wLD���.����c��I�ncf@�#� ���K�w��++[���*�*L2�>�m��d�z3b]S(A�rYƀΉ���>�B��!��m��t���`����c�_Ù�m��5��҇�"ul��,j�ء0����/%�!��e�[��ԭ1��K֕=o�3*����,1vu��̵B�#�II�^��멫���mh���c2*Y{�sZ�~�I��f+�[����x3�Ϸl�~iVO��|@j�j�����_W�,9-����`�IA��W�9��bD��L/��?<r眶֛��D^�3K�Djq�؂�}3���]�n�[j��"�a���|�����72Fn�J]8BA�ƭPߺ����80'z���� 	���TM�R����I� �j���3f;�YaO�׎9���yl�c��q��2�2���VR�(]�!O��xu�]a=�v�n%q�Z�=�C�\�0~`Uv�Y�$��%2���sE�"Q
�4����ɫ2�a�a��EX���������k� o���@b�s���o�ǰ�z[$�U�(������dY�:�KQ4�)΂T�+d�OYj�i�'a�tw"��k��*fH�\F���o����K�a�|2s7M��-t�M�R���F�����^4��s����ҭ�fp��o�F+�E6���)�w%
����ۡ�������C�P������W.l̫��g',���y�����e�@� �e�S�x[���1�~:��\	��e�����D��� n�P,�dh��P.Dy�D�F3�/����R�w�.O��#��}E�Ҡ��D���Գ/��Q�l�E���i��T��ݍ:}XS[�����R5<"$�!�<��M����g/��o�a!yz%�y]��ŋZ�:pp��?�r:�����yz5�Jd�^Ē��k �Hp�YqA-��2��g ���6�F�j�ܗ��u�o6������g�7 [ny��R�)¡�V�s90I��Xi��@�Y�@��d��7mI
�(Gz�Vz�!��}�y�7���G���z{�����4t=�ܽ8p-�|[�j6���H�՜��o>"T_�//v�[�-k��o��*B߶Z6
pX��x�l�do�!��voL�7:}:V�b�ASD�#�F�1��c$����Z�{<�7:m��7^Oפ��1�Ju�]K4���b$��d�NcX@4��AY���2�_���z��+����e�Z��l��B� z��y�ϛ��ǌ��q�<J���(((�~-�ϩp��۞��K� 9�����C�MaW�ȑaX��lՉ��aG��~���`���w��U�i��E*��%?u�-�4��E��n��{��58�R���E	]CK'��̺�V=G���f�l}>�G�+���dM��K��7��[�𪑡��t�$K[죹1����[�y�,�:�ǜ�����B���	zx!���h�� s3�����	~����˺j�3�wU�)�sr�H�*�!�\aM�
�8��r��l���+͗�'��;��ņ��GW�httJ�~���6p�VI�z�׿�O�ril�=�o�[�"�l)��!�M�4�R�Z�����F�gD�}xkc;L,P�E"$y�h�C�{F�Ô�0�����Q�UBk��G����m��J���t[	�S�Pd�\��Gܿ��`��h�q�ؙ���c�� +�5�_�hz.Wg�Q��:��O�ht�WK��d��)��F$C��h���v�����#�"��Ru��}%̇;��:-�X��!ӗ�\HX&aL������RB��K���ys#���H\��1_m%���n#�(�D3��"a!7m���,A�`��gF�&�"p���s��o���  B�D,�
�Mӣ���qY�2o|��m�� �(�$�d�?�ݙD�N���lU��x+��,΢$`V>�^��N/��m5֌���P�|1��9�'=;	�?Dfj�f�[�� ���x%6��Sr����
�X#�Kb5���=Ʋڡ�B;��Z�M��#�x_��1�k�=#kN\�A��'Jq*u�!M�!����Mt�/<ة`�֕�y���6~�f�f�X��) ��[���3�3	v?���Y/���d��=䳨zF�f�U��z}�t��s�:}ӧ���>�>�@���S�2v%WiGH�m��}2�:�=)�R�I��A��g��
4�^�t��ěi�H!��T�Y�s���\�6�����k��+��U�o	Gr��Ιi>,�8��*��5�a��ĝ�k�ɟ��_{���)��͗����?P������.}{DO62͝,=�N�M��*Q1YK=�3��}?={���Y
�K�����Ȇ���<���Ґ�&�B;����@Q@eM��]���`dɅ8Ҳ�������B=����`�Ʌ�:ҹ��K4{J��a nz�W�Ĝ8��x׌�2�p\�Y�K�ES�T����� ��ׯ�+�@�b��W:��-YI�@�b/�]�GW��8
�3��,��[��t�߹�Dg�(����oDb^Y�l������I �NC�(��$�|��+��iXΪ��0�����g��q��ri�`���V�S��`]��4`�.���p6���p�M����&࢒����VU���{��?ua�����J!���|����4� ���~9،��}�l9 ��#��E��ܽ!QJV�&,�HZ�����9�Xn�:udbb��d�_�G��]� 8�Ӹ0bs�Oܶv�;�p���u�$�}��7aǈ"9u�af�G�\��9@Z����V5�8%l�+���N��A����;�z��+�CZ�q���5E���:Q�ᢶݭ.�81��r��>W����^gm�]�uC��C���%u�)"��궋�3��iW�FT8u�>����~�1��-?_|!d�@
�	Y�o���y�ع�,�����	��=]�o֨u�2/��,�g_6�B�*�a[�N�:���~]m�`�C`]
��Au?@$�+4��>Ĵ�u����0����T�K[�b'qSS���7I�5�2Eu-�hvw&�9�� KIշ����A��W2b���� ��c��"oZl˔I ��=CP� �s�g	�R��H:� �lF���n�-b#v*f*��J@W�%d���͖�#.���j�.�a5h���(��Z>,U�U��m���-�m��z�'hW]j7x�9��C�8E�*�
��:�C�@ڱ���hţI���LbB����w���(T�|�;��=�~��s╥\�e�i�c��23H��Ύ*�	�K1�'���j�6��C��rU��4K�#}��v����¿�ga�s\�r7����s��n�^�I M�� ����j��/Oe%��t�_�d�5�QHѨHr��h|y�,��B(6�w��[��5�bV˃��9����	�췅�}�-a̝���<����v��be;륁�dxM��p��jYn@і-=E��3�#b�h8*�.y{bĔY���6�x��~���-��#N�l����ɂ�N{�VWm��!Ǟ�Y�$��~�?�@!@e7�`���T��ᾘk3p�)f�{�$숖�"�J/�(HS>ԸE%��B�d�dr���w��ӾAdb�D�D5�f^PS(�x��9�F�gݯ����1��C�]e�ŪT�Q���0&i���>p�C�q>γ��Ԉ@e���?0��i�<ZY[�W��rk��rUw�������.�_/�ow ��w k�Q�?�!�U�:�t�^��␴����¹������Ou&9rXMg�cD���y<i8�yp�+Un��r�+�ي-�m-���n+u���iY�h?���=4 ��iӅ$W�<�l�Qi{����'!�؄����چw��w3�~/F�X�Ger΅��f��%՘i҉OӽǨv�}>�EA+�^���8��J��D�@��b�������U�Bm}pe-I��j>�'�!#G(�$�uF$V�ֺ�:�';G˂�|l�j��VJ��,�B���:ئ����Is<Xb}>ֆ(�������v�:�N��sS{�dK,�������㷆����
�S�P�!�eh�:hsk.K��"?է�@�b�8E�	ߟܚ_��1j
�h>`ɤ+7�vi�@L�Y�/�p.x�R����*�o��'K7v�����뼉jL*��,@���* �z�V��2&�6�i���w15����D�efw̞�B��7�~���sI��Դ7����!+�\�ࡄ�A1��k7��Ź��W��Qh��a��j*?)%0���:2�sA*��	xy�d��fzu/�������HTQ�5rB8�=@��Nx}��~���K����,��٤�B�����q��sQ�/ԑgC�F����jf0$ָ>���K�E=*5u�ĸ��
�U%%E���X�U��$H����)�~n5E��X�$�9�K�*����&�T��◮@��I�R�CN�6�#�A9��������/�u"�~*Sm���&!!�	V�k�m0�S�\l"]=�����+V��ݠ>�=4�@��qf���h�p�� ��0�5�R��5eiWzZ�^<KÆQI�(��q�Y�~�^���P�~���ܵ����Q��M\YM����t�|��ꘔ8_���onܨ�x[gFjKe����U�o�=����wxm��ce̟{v�*����R�h��p^D�Om��t߷?�NCO��)~��$d�i��/oi��6�="��;�:����3ڐM����phN�2��
�]g���L��bPw�'5*R1�H��EM6�o���� =��+�����)_Z��׹-}�X��:�(�|�\ߤĦ7�I�D����-�[��r	$��'�(�]��$�&�w�i<���ta"��:Ba/�Ds1�wd'�
Mg� �a}�A�Rw���S�S�̃a!V�\�Y9�8�1ڤP�����&ȭ��0m���OO��<�<te�����ѿ���=��)>��٪�ڱ�h�%�w3d�kA_T@�D��|2���f�g�%J�k��uq����`��=�ٯU�'q�z�qқX�jGk.��œ^�@!D��i����6<�r�����V�u�.�i9^���=A-&�bSַ��B��\�㜐{�Yg���0��ݫ� ���2�FL�S�1�$'L��������!mPq�g�ުz��"0�xz�hB2��DQ�dk���5M{K�x�%���G]�c�fG������A�(�A���d�Jz@��+��E��V���uc��r8\�T�
]�}��*������e���� x@��;X����9�a�*i�V��H�� �C�;�SP�b�"{�-�@0�wޙ��IM�����:��T���(���`*������Z*:ǭ���*��7���p��^�u`��l˒E2�Hj�_����i����rچ�@?|W�l����J &!@ ��Sˍ�#�2�/}�����C\"Mu���{����&|� �X3�#�����%��`�GBd�j�ʈcK��:�.,ĖJƪ�N�Ť�l����`?�\�p���~^��FҋA�Y���U*��8�a�.�B�%���he��i(&Ӳ�ɳ
̡�c�� W���D�T��Tm��Z58�3���x.�gH��]�����j����Uj���;9�ƍX�\��/O@&�%��@.���NAYY�`n|Y>��|����i�!�a��� rF ����9�A��GM���d�H�$�T��O�5�A�:sL@�0�nѶ+T`�j?NKb?�*^���I;5�������G{T	.n���_h��qlY�'�;��Rv�v��X�����u����FW�
ɪB��/rB���@�d�[�M%`�=�%ԯ��Vw؍u�e��S=\��x��K4ɖ������#������[�rF�y%�'�~�
h�����`UL_]����E���r0�>�^4n�������Ee�3�{���Y�x��Z���\�띅�&��09��{U�{f<�F�1]�*_�������6͏i7]���nX&�M���J�x�(��>1��×��X��D���|����T��O����gU`����O�\S�-���"��Iwdei�R]Q���jW=����}&Y�j�r����9��/�į8���3�Acژ��V `jz}�V{΅�b%����1��R8m��ƞ���
]36u٢3D%-S�=aXcsuE ,8��� �i�)��+��֡�����0�a�彝�hh�
�=�����p���aH2{��,~e|�8tO"6�,e5�i�x
3�؈5�v����L�t�V]"˶��v�x�B�	.0��
��:�<Hu'9 c2��v��y���b+o�T���QO���q�M1��*Op�K4���v��Zn�?Y먙�0�@���EJ�J������ݛ�ǡ�N!��w�<�;+)�|��dЋ4�b���)$>$�? D���v��|��7�I�)h`�̳K��d�|s�ا<�V�.������o�E��mx沌�rO`��6����x���G������5]\6�_guF4<�[�h��g���Mq��3KG~-ʼP��D��Q��x�J[O+Ҫt!�����o/����\&���1{2j����u �:z-�s�@���p_�*8a���6�E0_�L����I#9h!�G��x���tgoE:"
���tN�OB�!�+����2�GR�ɠk��DR�.�[7�5}L�N+Vm_��s�՚D��1gs���V�t=m'	��ʴ�z�T��/�(�h4HJ����H���TCO �7~�]+}�޿��!��&��P!����J18�j��-�5�5@
��`�+b�I_E.���X��:��m�0c�m�H�ϯ��	vq(����x�\� ����e	9(�'��닜�پ�����;�F���6����Zm�	������̼z��Lg&>#������uv���n}��#����o���{F�N��nw��m��;8na������Y�;��X��V�-�||lX��v�g<x!ĒѠ�l�f��7�m�Ƈm�_�2P\��`��[+���\ǁ���dOፅ��aȒ4�9�]��|���
�y���qW�+����B&W�K��gU�����/^�;�}H(���b�(~�����R�[ň�y��Y��d6���	INC��;�c�����q�JܶhR�k��"hM!�P����ehտ�V��:�x0�"�/��M���Wq�6��Ȗ?��^�
N?*{�0�W���g�?y��d��πVʖj;N��+�v\�Z����d��pB^��"��p�qǘ��s�޿�����y�fp�`d7��/2����NkeEl�R�~[�M{u��W�a���U�E���X:yz����o3�&�AK��(aje)"��h�y��O��0��m8iq]��V��[�a@3=o6��k{�e@Vg5���"4�l	��WL�m��ʄc�� (|[(l�K�p'V��Dkܨ�j6g�R]�X	�n��8y�'\��W�j��#BS	b����H�g��7���q�r6�9�QpE�1}�h-��c��X.4Ћ.VcK��k` � 6��Q:+�6�|�	�=(� CM�{7A��޸ؑ����W+gʯ�U�s���LP���m'@�e���M�ԟh��s�l�t]�6��:n����<�A�(�����}�������\�kq��&�g�G�`n�@��b��iYn�/�,|��2#��>��Ga]�#%�����/N�C��]|NG�=l����P.����Sv[�`穫�d�w��`��/�8bm/ˌ�s<�b���;�:�Uc��.9��y4�W�L[�h��\���.l��UkU�&Q��8��8U�H���ۊ@�K������ »A��y���M��~ �+�+�M%pC������iɾ�$��>�TR#�7UY�Y�:U�B��X��(a����z���/r�-@�K����Af�}V�����c~s~���g����	�nj˧���2pAW��BZ|�'�ig�g�Q�4����5h���YT����q(��щ �kQw`���(��>S����M��������B�μԵ�}������(9��W��ӓy�R:�H��#�;K(-�J_�n�L�]T`�!��yT��*{�����b�)t��f��n�[`v��
��!S�Բ�[�C��Z����VY="#v0������kM �zE��to����pa�����*� [���5"id�+ �M�.�$ qY�Rh������Ş��� !�ѬVa��ύū&En�#Gµ㮌�=����L�Q�Θ��>'�-?��e�o�r�.+��Pv=�%je����8�܃se
�/u;vU���S���X��}{!v.7=��A�?N��U�Ήr|d�c�ÿ��� q�S_h?��=��dA���%��_�ghT�LV[���lOkj�x�������>�gS�Ll>�9ݡ��J&xO/�T[MK��zύi�}-�F6�c��_� ��:�bT/�x��[ybB�wsE�HH ��
�;@NY�X�SM��7�'���*q��s _�r5"�,��6�?y��FB����u������u�~�>n5Z���Nc%��u�4�֫b\u�4��&��6�c�g�
��?s͊�U.3N��rnob|%~:� ��������!���b&Ó���t���c#�"��������ڽ���Q�LA� �p���p���> �#�E�oyc��&���˩�q�
Ku;U/8��vZ�d��ςUϚ5�XFH#9�Ort�</�������`%��J7�we����W��b4zp8:����u�R��P�(�y�0$E3(0�OA�%��}�J�c�	�[Jgg"'��&�8��3ρ���#�\��&��&lم��_y����@J�vL>�+�ox�)g�Sa�Z���uwe<�ۃ�F�D�Ǝ'�J�����Y�p�PL�Oܙ��Q~��ɬG�]�:%!�Nx_z�*�3'`��(VL�v���ru_'��cAxW�e��$�7}Z[��i��sH6|0��[sǏ�?��^i��G�%'j���*`��Т�ofa�j3>�hBZ�<�\�J]}Ϗl��=p?�hV�b�\9h��l�Ec<���� �:;�8<�]Aw�%�8������׮`�.�
z�
X���~3��,}�Ըߐ��)���K�id,��%E��E�^��N�������S��BC�FeWe��>���5/���A���?��\�k� 5��Pl��u)y��K�up�%��4j��/V�������9���#]E�J�����v��Q�dM)G��<� ��yd��-�F0�.#j&ϑwY>�C��m�񿷵�t��LNH�T���#r�Ta'Ӥ*���L���z��@���5+��B����E��{;[dh?�J)��<�9�	�VA�l�4z�2�Fq-���J%wjG��x�B�h�dU5��a�I7Ͽf���f��?e�W|�Tr�+�)��d�)YF�_-+�򶜘��FW���:���p��E}��76Svto��������o�����8����1�R����ӑ�X��IlR�^N��i`�P��[t=S�l%0���[V��ލ��>f��QX��ҀzD�����f$;	c��1#�,TW�� R7vFl�s	~���W�*z跌���>qd�Bs5�#�w���IZF<�� �p�Цy	H>��)�S	D /�:x�����>�CyX������=���NCi��iM���Lo��˟��F1�LW�<Q��H��}q�^�o��Yx�}W*���j{	yO��|0$�����t����+	��$M�1���I�:��1 �I�۱�x��ϕ�d�ï�f1��te���WH��(�P+�_��+U9�.Ym�� �� �}����%��6�|� ���#�����K�O��Ek3@r�7��/�$k��v&�f��� ���E���,�A���c�ii��yu���x��g;���B�`�#����
����M�dk�V��kϡ�	ŧ0�����q��>�����=[ɂeL��&q���Y�P���ŝ�vTKh������/�d�d�(\�9��f5��S���9H�`�^}��tx��O�ʯj�H�L0��+�.E����g7T�&�l@}_�'��C��w�_|�Rp�=����ۧ2I*>��D�n<ĕqj���9l��A���(������L�B�D�{�Z�5�~dGSi�1��}|�p䮆<W��+}�������}��	�S�Z��'�H�4�|�� ȬF����*�����)�Q����~�]`e�\�)$�>������[�>�R��L8���� >�l��M���c�UBR8�1�Z�.*D/~��Ux j7�Z�ꍗ[N*x,��)= \r�bVT��)�%0�� -�ݧ�|���k*�.V�M�9]�U�V�uBP��C��C����@О�2� �F#5\���$�5����B0�F�.��ö���_JA�"]�y�!�R\�]zmb���ǐ�΋ɱ��~��F"7]��/8��;�>aP��Nҟ��ȇ�<l�����Z�]q�,�P�>\ Y�N����攞/+�$VS�BA.�5]MTo�.�s	>"a3¤
� ��d��No�?�_Bl=1�T����.}p�S�'X��3��DRl�+�k#Y�T!Gs��������p¶v���vk^-T;yzY}�HM��SR��~���������y)K�E��uMyi���#�QC#I�X!���b�ձ�6�J�U�*!���H���9��	q��C:&������e�8]T3n���=S�i-$Uy"oI�s�۬'����G�飑�B�!=l=�8"#��,�8@"r��,�Gmr�<�3�{������ֲ�ܟ�e����wm�rA�g�r��+aCe�!��?P��ۺ8�{�5`x<2��X�w�n��4�4�!�<ӏc9�������w����gysr?e������]W��.Ŧ#��T�		o-�M}8��|1����Q�ӨT��z�j=S��3��>3g�����?"�5�#g8�#�.��qX�~�N�hG�3,b��DR��`r1�������ɃE̷�m仇�l� @�*=A[{�e8~Q����1�K��§�o�X�@A����ƚ�ƽ�`�f�����IOG,�c-��i�u���WP43�9r�������X���[9��˩&��E���% ��ǍeS��,Z(B+�l�Aq�B�6@�����c�Ô�B��PJXN��l������"w�|��ΗB�5Oc��1��=���g7R��{��a���X�,���
f2�=s���К���z�?�j������~�<{PDQ�'�b�F�
���%i�5@�!@���_	3"j�'����q@r)[�4�_��8�k^x{Sz4�JX���Ժy����R�w��JM�b� 6�1|!�X�!��SH�g������{�
e�d�8m��K;��F~�[��]Y�)[����R��	�(���ыT�IQ�,�N(�偭�D��pj��F�1f�n��&�$��lѤ��uL�*���ɮ2)�,��������x'J�(Q�z,q� ��� �T�fUW�}��~t䵃�b��7V�����%bqzX# 
�NB��m)j3�C87_��H��5�xe�xL^�aR��وL�F�����F2����}~��"y,�i���_��~B���@Ua�d����YJ�����1����B� B��%�hr�@���'�����v���%�b��-����Y�gwZ�M�g�7����ҨH����B����j�n�tD�6��$`(��D�g$䲃R	t]l|F!������#.�~}G�Uױ%��ͫ�1��+�Mi� �o�,�:n��3����/��z�9���3��7x�O1y?\j&L���XC����6p�5s���W]i\�{��LCn���Ә%�s�勹�� l�3�AԊ��
Wvjx�JJ�U�_�� �%î9�g,;�G�	�n����j�ɮ<�b#�c�:Q.�ۛ)f�BEy�0����hq�_T��6lG!l�j�{�� @�?����G����+� _�3T��ͯb�u	�Zm쑲�|t���r�Yւl�B1	P�$��߀,!ڣ�É=?;RK�Y,��VɶP~���f�1���F�Ga0wO,��8�iM�����ߢ��a?���+���ǆ:�FC�������,���.Yu/G�[ۚ �P��B�k�ʛ����h� H��b#��Ɗ��c�ډ�`\c���Ě�>�_�Jk��7�9�P�3�g:��U��;NYn��v0�^T�/_tw�2�uv�%C ���k{��ر�����ay��lpP����]��E_Z�l,NA�g��F����`b��L1d�Wa�_�,:zA���O	Ý흰bn	C�#�?J��-Kj}Cj���J�D�|��®�.���}bXoe:�2z�%��>��tpQ.����׍�n����b�>���ҿ9R{u�03:�܅:��B|��{���G3\;�<�>��{��j�����k��~P������9��e�|7[�c����ĜW��[L6+Ԯ	��a��g�h�VP��O�����T_mv����z!C<57@
M�"%@�ý+�5��l����(J�"�j#B�lw�_���1�|��L��ܧ٧�t����L-�旽un�dV{
!/����6ݥ�rIuA� �7T�X�R�㦩�^Woe��Cb��jߢ�P�T'�A�TasDz�X򽗼��7��g6���1X �����2��]7mSU����4%�c·�{+�Yo��ܔT������|�(ia���1r�J�1"{ܴ��Ǌp��K�Z���ܟͤ��F�<[K�+b��@a�)P�[�����!�e�AtMKb"��
��#��N:����ke	�'-��o2Uvt�_�����\ê�-�	O��Y���Aۼ-�9�'�'���\�����"���T��Η]^Z�@����W�/q�^j���Xe^*{�eW�Tɹ5�կң�����0-���y1z6�c6nz��E��0���1G�\	[]�]�۾�]U�_�ؗ ,t��E&z!�a@cx�j��~"�p6�6�В�C���撴`H�oԳ���J�jű1`��Y�8�XL�� �aFL� F�_������j��ɓ�A�˫G�����wZ���!��J�F�PWbզ��"e����<�[�p�!�}o0��bےS0k���1z�:Mf:x�\O{��:��y����������[ѕ�?8W���ｉ�r�L�����'֥H�T��Qa�^�V���8<�wT]t��xmy 0���r ��B t���-O8��|��9�R�<�|u[�/��/#���[��YM��T��2���YVbU�ƍZ�ү�0J�~��
O�� �[`�a����R \���#. �zn���_b�U ֢wy?]m�}1#��>k�{�&�U<�'1����$}��k��= �]����L3����H�/JwA,f�PPO��|U��^g���>ϫ`t�T�m�pEt:V�����Ҭ?B�J�N��pW�\ʐ�c#&_r��=��Βc���3�/�^�M:#u0�l;���屬߳��ض2i˕7u����$8u� �F��A�5ph��֔�QЦ2�1�x�?HS�v��w�K���2����W�GFb��-^��5�x�x�d0�^�%i�L�e�y��w!{�[T�gB��U��͆.TEё�b#	co�Q^�c�����q' ��p%�pR{�l� o���+f�#F�=�h�����r��ay'���gI��ڐ0����BY�l�p��f��5^q8?o8�2̥�S������JK*�P�w��0|-2�x
8']y�	��vf����-�y|��OS�{r+j�,W+��om��ze)����j��앆w��=�}7+�^�ڡ�D�z�R.��I�%�_��iq�)��r�b��:X���rh�&9(��L�oL��ꊍn�u�Q1��D�O�e���bFr.P�5���&��l�����M|��5W���յbt��sG�{�^��e���i���Kw����kVQ��v������}�|X6ҡ��R��pk82�j<�[�
0��V�b�`43�-�k�ZL���w�i��p���2���)�����a��|bE��QFq�N�)E��<�PЕ�s�g�_��C��ێ��c�W�$$�g(�R(zJ��cS��uGP=XOr�.O8>ZN����Z�3mk�T}�ی�nq#��D����߮s�����-��Kp��ecsĠk�4ɫ�'�m���MȽ���B�%Ų2�z�&s�t�&�zP�/�rQ���#}VT�b{� ��%�l��o�>,�Lr̴��mSԣ%OX���_�VQ�2�U���/��V#��!��_b��U�.$nc�a̘іkξ�B�Q�g
�LޙG\,9�k�F�vP�y�L_�z�@c��D�T��s��������±W�Co��%�B:Y�#|��kZQ�	�T���eYx�ʇ��8"Ў��M��0ȋ�yN�3G�L��+�d�"n��2~�Zm�9&�ψ�%"���
x�8�����������_�g�L'Jj�!���y��[;�èUE�%�Π�k���1�Xaڑ3�����.��h�����1iiP��:�>k��\9�z������r�R|��� �P+BZxZ�#���s��^�,ԟFP��Q�Pj��{%z�h��p��f�|k�x��k�ߎ^ߑ������ݩZȭD	Ɋ�7�f�������GKG�t��ځ�Y�=@e8��#���B����0��c
�z���@�4�F�/�jZY���Z�2�������b���#۵�J�+mF�F��f��fi�����ҲT�ŷeGm&0G�v�<�4�P���9������4�0���DK�;���V/�b�G'Q���z�&�*�@��6M����B��B���|l����4t�<{bo���'n��
&�7�?o��6�wѳ���q�0�*�c>�B¦&���I�t�t�S�8�������5ou'��C&FG:˘>G�����ڪGCl�i-��W����E.:���-y.�]HH�.�`zhċ)���"�����Ւ'��xΘ&�@3��=x�!���^i���*����g��x�ٓ=a���
ݢ��ES�?R�+6Ꙗ1k�
ʊ#�3��+��$e�8_$�HR��Q�)H
��"�����n������ְ��:;g/�6N�wyq�Y��8���c���Xp���/#Ĺ�+�����鼕�w}LL���4a��J]ËZ��d�<ϤU�kI�'��w�9����g	{e�t`6d��"����jy�����E�Y:g���x�\{1Tc0��m�	����� bk��)x�U����y� �\��U��?�J>Fo5#d�6�.�M�lw���W��L�/z�K��E�����"S����C���Y�7�Y 
�p۔�'D��3�&�oa�č�5�O
8�)oz+�q±� h@�˗=b0���$2I�۔�o+
m}����c,O_6	�V�sP=P�?���7N3�$��Oj��jygc�$��!�j��:���En8�����E���޷c�m�64��yy1'8���ӝDln��#"���(#�
�,�RXv�����+���R��K*�uC��R�+��~�1�7[ �|i��,lQ�g��V�� �¹�@5S���>k ��ۯ�K	��ȯ���'�U2�R��A���֍r����T��	A���؊�1E�:M�̥��|�ŠU�'<^�'��d�Y�5�E��J�82���.����h�6h�����������[�Ey�����8�ڸq�u�n����<bw�0�k!`���_ '��mtW�y��U���0B�⃢�v��3O]`cOjrl�<�1ΐ�y��G�)���ڃ.0<*�\B���Qci�����!O�}��uS��P=5R�ǓғLk��{"��*��x�=�,���T�<#Le\h����ꨱq|�¹l{��W�͉{������ɓuU,t4'M�	b�����)�VW���sf[l����w��愓��R�Q�%^׽�no(
e�<�W WUq���T�N�1����(��j%T���Kc���⓹�nQ���*	gy4�u�^�?M��@���Іi��[�b4?xzMӺ����6��@Y�K?���D}��A}{�H�@��щ#be!Y�A>\)�}�V�g��gh��y�fC{�8j�X- ���b���ĂY�����_e������{ş99���������u��-���ˮ+�g�X���O6�gv�y���2f�}X�Eu�BM����5�R�����񦈼c�ݸU�Ok�zDlG�s�E�2�9A���4mkP$7��UǗC���Ü�҅n�'�T������a� �S��}m�gّ�K"�J	ݹ����N����aY��������Xb����<.�b�)z;�g<od�;�&/U!�s�A�Bߟ��$��G��Q�Y�%b1�1���CE���m&����}�r�8{����P��DRm�;b�<�I솛&��
K-f�*`�5$�r�s���v�uT���BԾ5�#uW7a��~��%�s4ʥd�9�[�@}?��㮿T-T'A�W�q�4���";;�ZL��,+ِ%
^Ro��'*�~�}E�k�~�;��0ݜë�����4H����F^�b*R���P�#��	�\,��\��V�4��׻�}N�F�?y�<���c5��Oұer�Ҭ6��:P����]��@�
��jʎ��{��]���K�tB|߼��]w�ig���6p1,>���d�T=�5��V\ ��b ���,L0`��sg��蓦f�����0^��>�Y&{SԨ���L 3 _�;�k�~�'�R��5��͸�}���Pܼ8��s�LN�!wp A���T'�
��#G��K5�p�Y#g1{*�z���<������!n[t�in�0q�c�䞼���u�j�f�WY:���:�]�ڿ����H���>` ��
*�I�BO�zI� ���$�Ç�H��Y�t�[;=��(�Ĳ�6��+)�X��(+.�q��9�^�M�D��M��~-_��JؘË]��)�x�������Ȏ�5�*W�1�I�qf��p���4V�0zM����P��S%��'�;1=pR���e��ㅆېu\���(]ȇ����#�y@�rV�~�a]�]���9[V|����G�"D3��:���Upk"���/�v�*��m�B�-"--�Ќݾ�ɢ���4�yʱ�����Q#�C/3gR�����Hw�;U��\��(�I��U�κ7���>��x�>ﺹ;p��n<rE�eC�_u����4ث�oW��a����IL�y�+��9�x�e6B�PK��jf<Q6,�6�7�룕�{�"�;a���J���;��t��F�^��2��f?�u��6=�v����a�R�!�짉ds�YT �J��-� ��m�o��҈I�Vt37�,�ֆ�.�3hJ�Mñgq����ˇ�[�Rө�$���Y���K�Ӗv�UƂ"��Z�yϲ�������=���p�o|D&M=Ï��6�/����i����V�T�u�#O���t��4�M�9����
F�$�dA�ޅ�Ylb(�l�{p�	�@��}�5 ��B�j�d�M�x	D��P��!�c���� ,E?f��d_`w�.�8�����Q})����_'��!8x�UƙB;�mߕ�? Rf�����C�u�E��!]��WA8P]�j��ol"˦w�S���K��K	�~�����KWL�����-W]�q�؇�����O,fj���q�=�*rD<��ol�ޛ�&��H�p�2��-M�)�Ar�e�K�6:���A�CGD��1v�A��� �`���%ru�u}Y?eh<��	k6q!	X%S�U��!����#�]`�RB}�1�
���7� �뚧��p� �؝�x�ͤ��j�w�I��@��L!I�n�=��F|��v�)��Ė<�tɜ��9��#;�ctܐʧ���i��S�z�+�j����R�)�Jj���3�-0`������_a[a����'Z;��z��GK�qJ�VC(u�d�Y�M���a�4��qc����:������+~sr��(v0=�-�I��]L2|��^�7s.��s)�r�Y��r���҃��ɖI��m?��^Ӡ,���,m*�/���k�n5ɟ	�:*4�}��쟃�9�ɭ��@���-��X�?F��u�H�>����V�:��G���fq{�
|�]�,k�ч�/�x'�Goo��j8��1�Rׁ��}	U1�;��� �CS��U^<�/5�����Ml����p�=�"�:�3�e=��H�8�7����Nտ5������n����q�_#����+#V�֕��l�iY�&S������~��=��TOZr�%7Vbd�ݒi0������H��9�� /�?���+B�X��k++Cɋty2Wr����?�4) ��\ͪ�gP�Q�ڜ�Ili���Oj`ۑL�K����a�r9��&vb<׻���7��{�����Ң̾�J�@ʞ)�1�E7K ������s�v7����3�����G�T%C�r��z3I�?7�P�����_���|�'NWzd~���M�l�ǎ�'4т8{N�-�؋��qk.jj�����h<=��?�6������@�Ďєd�
��i�S����o���T���:f�	�-fs����ke)Dr���s�/I4ݘ��L�(ן]��h��O�~�ѽ*J"�YN\yGM�_0�d��ͥ�l��F]("K�_iP
R��םe��s���S�,2��ԛW���7��	�k��4n��دi��c���J� �"鑅E�E�GcC�����Mi���9}V!�2�8�m\�n�o��*֣.u��F�Sh�3
32zdd5�]��ЗL���6��=�^�LJ�,*	հ`M�O�׃���Æ��#!�����o��]��f#|kx�(���q�&*x�%��ˆ�]}�U�xw��Kߕ��b��.�76�a��JR���� ��{���B*�6���	��n�s+���l��Q��-�����庙^���S�y�)�ZQuSt�ب�	����[^�H �+��&U�A��o��\�|7��ͬ�q K�� �)�?��O��m�*5�u5ơ�!^�����%���oC{�SV;��M��3��� ���X�i�<恏˘C~n�5��Gֳ����`�A��j���W��(5�0�S���d�+!]�4��#�+LY���h�g�H}����(��'P�dG�������{<;������:U�9��(���Kd77�1r�;1Q�|��hWg,"��d��WKIŔA�y��E�u�"M����4;�L�!�#H`ն:��Ir����Y�5��C�O��IΛ����ɫ�f�c�\�);-�,�;'�*' ��)5�i6h�D]Q���T�F�����3�o�������.�WBQ�L}�����'~���c������J��!�M
N������R�����ւ��\�m
1n��&B���ӈ�T��L��P�N���@o��l�5]�����}�[ץ97�/�
o��?�
�(��˔w�]�7��a���";�\N�L���>P��6"{�1if�"}�F�e�;�6�8J�j(��}(��"�hPH������҃�M�af�U�a��=�,uX�7����a|��E�����Rj!�H���N���X-H���"�_P8y����G�8�%+�1�У�e���B�cm#�]/��<=����&7�_�q�/�) ���^�b���Հ�1��ƶ	��,����*f>`�Q�\�iIDCA!�hY���yC�,�Wn��fr��N2�6���8@��뇔8�vB�?��˝�-�q�>WHe���`硄g�'���/��J����Z|��m�(e�����Tt|)�4c�>O*�T���רk�)�����*�-���T�#���m�@\�O|�!2��i��jQ ���P�*,��ظc=��T�C��=jY�?]:�'�u�W�g�ϻ�a��.d��nЈ�[o�<��Ϛ7��^�(�u�;]T�# �����w�_y�T>BB�a'{�HKDy������Z�����m�m��ƈ�����(#���z��qj�}��a1�e����{�)geG�l�i��Q�;��%���fL>��6J�X,¤[dV��de��2Z�Ĝ�E�mu�������=���H>�9(\g̇<zlT �J��BB�vˎ��e��?��RS����&2�F�lh��@�Xxri�؍s p��k���c6�o�}���	��p����l+�_����1�����
-�)�cs�JUOv�#dF���+�֚����X�@��� ��)�9�0���7^�i���T�֪7������K(l�+�
���^�;�M�m�VOX�tm#J�Y�Ty��Í��y	PU��"�����M�|�?_3�Ɖ�GeB�}K���&�|h0L\p�˚��"Դ�l+4�$^*�čT=:u'�	PM]mAF�\�%��&��IۭTB�A���7E��fO_�m���'j����Q��f�a]{�.��nਧ-��cs}!?���/eW�F��Ybk��j~�G��Tئ_0} 4��<xGk���wx�r�
KD@�x��Cğ�
����l��Լ���	>�&i�Y̺���1G�A]�H��7�4@[wE�W�}h�N�R&��j��t��Q�<�%Z���4M�8ꦡU+���C�4|YKQ��_�0Sjj�.[��WϦr�V_�;�{�O���݇�����\���!� $���Ou���L�ew}���(��²,0�T�0ET��D�ǆU#���.�֛��m�v�ŖNiμ*ս����J��c�k�����$h�ė};�D��z���H���������isGrnj�.L�䧋�(=(-O�t*>�?*�(�C�kSt�1���*��^NЪ�m~Vp�>�L�/L�)�������l���>�]�*I��j�uS��#���=dvs��+$W�_�%�T�Y��� U��t|��w��xo�
��V�;�
��ZNi�=H�_됌5�m(��	�6w%��xp�B��l�r�Ѡ@�dHn��_n�6T�k�S<}�q� �P�A�0PU-��C��#��ߗ�j��^�'�AJs�1��%�Yvӏ�������3�P_7�A�[ u#������ԋAϽ�H?J4��ȴ{��)�D����,@5s�ɔ�]�o������,����9C-t4T��S���Qt��WO\��w��w2��欍��*ߠц��&�{��"����ڜ���l������A�����q��q���0���U	���ռ��'؅�C�0��$��
�fCX�]��~t;�&��ZP�U4��>`�f�փt��L�?�ˌ�`oAc��Z��=n���<`�A��FJB����`�w2�!����V��!Uq�\R_ԄY׆�s�O��2g(��
���'��!nK�g�Z�;g��}��4WI3~�W��g�hI+�<C�3��R�>̢�I�d�$����c*5Ə���K$�@�ܻUv�Ҷ�U�����P�<���Q~j�J�B�MW���m�3z �E9��`U��^�{��캿M�)2�Y�b'ü�_�"뫱.Y<�
,"�s)����2�̙���������Խ__[Cܘ�ػQ�X��ċ�n��G�s��jA�?U�5(�/�L��h��t�;ro�M����=rN^@�/C�c�8�[qغ����� �h�jJ�j�j�]	�}pߔ�q��p��2�`}F�"<0~�����OT������vŞ�p�<���Uz-V��_����nJ�7Y[�ye;͂��|�C���sJI2*d?��4kȡ��P#���DL�.��X���҅�I�1��)��!aR���V�4L�i[,���yn!��՟��RSB�UR3���_��!8�WY�D������֝B?��3�2�I;���v���f��4�N�:X{�E�	{�@^j_E
�F˸�����g���ݾ��U�Mc�����1uP�E34��T����S��[Tڶ��	-���նސh�oޟ��LZ=~�*SA���n��r�����/�|6�O����Y�tK��.7�br�JtS�pg�毇wC�j ���"���ۼ��1��Cu �D������4j2�o�H��[��h@YYDU�7%�s-nt���������m-��k���=(7���8^�7K�d���W�Ti�E��n/�s9���-�O�oM���Ŧd�k`S�>��=d�"<�:����g�(RE����ڣ��67�I �̼R�7u���i�� ����9�r�K+�^)9`��g.�m����6��Ƹ�Uշq�ax��N=b�ʤ�l�R������7�3�m���j�Nl��:bg8�N�	 ��0;��p���Sj���������ˊ0�'ϨCT��{�b�P���{L����i�c�9�̈́tL�1�D�!^w_�ls.s�f� �.T�d���P�@�+#ʪ�a���cG8���S]��<����!]�phn6�O�K�"͝!���^K������;��xJ��>ZK�-�q!Lx���$vaX��VS� �i��� ~-Xgzm�/� ������<�̻���?R��d����oA@~�
��(rM1���E�+?���tg�I�-��7��xg���T���T�᤬������b�j)<'D^�ΐ:�y����Ւ��������B���x-%��$G�yDrP0p�J��Ӻ@���P�	��TKi���4w�	��� #�L��n����GxȚ-�/���I�!�-�}��T^��*nv�����)�s0���0�j[�v���Nz������F�c:��k��(`x��ŷ�%����l\[�vmPٱ�"��/D�T@�W���8�"c�:��m˴@��ɞri	a�P⃯��C���{j�fF�����1&���L�Ք7Ex�\l��W��Yx�����|��a�.�����9UR�����i=1@���V�Zc�&3�9r��.�>~2Cu-]�t����o���[��I��D=�y�����$Y�F��H��)囕�6^ɶk27$�GB�Ɇ�C�*�V�:�>�u���X )Uq��'��F���g�������FG�!��C��V�&�܌;��:���Z�L�$�]k�"�������	=���ƭgq�ei�A��m�C�y��%�ݟM����u~�ڂ$�{��,�6��&�r�W�w�I�q��*V�-B�iYʩ�e�Ĺ�A����G��ˁ]��*o\;�
2���W+B8ӎ���-vd���C��X"$�e2�����ꧧ�T�*C�o0*����X+�~�ի6p]�l&�r5�7%+�P����:Gԋ!������ɷ��#�ƿ'�^dRܰs�Aeǚ?M��o��%ʕ40���r?��5w�/�#���C�� _Wi��m�璑�F@���7��3u�N�p����`~�$�CZ��J�х��3|={p�fp11�ғ��S64�q�_��*��<�8�l�����O:�Kԧ�.m1&�KU圫����=*�5��C��/�s�S8N[�J|A�O�V0��wr���[�H}��Z0m];�������K"K���|;:ı�A�TV����Jc�я-�Q���f�m����z��Q��yg��Etz>����O|?��B8���Y�(��U	g�p��Ű�.�`OP=��閲�,Ut��ڇAijR�U�D�w?�|��Q��L�6�Q8�ћ����KJAc(�RJ��M��s#����b4�M �M3D�ч�|ji�e��P:�2����X�׭�GJ6�����n��4�A��ҶJ��yO�-/A�ֲ��U*�o:�]e(ic��:�g���\O����$��b�J�jԌK?s��̼�g�A��M�S��R�+�-���a���c�n�xXY�U�r.Y�Mm��ƅ%��<�������f�N��!x)�^����ɼ��5�51� j��jV�u"Q@�.fy%�Ρ��a��+g�E58��8A�/^[5r��7� �K���z�f�ܖ�G����b�ݥK)�D�i���,?a=	�5��1J��4�E�r��.���P�4:����Jf�`����GG��Gʾ�������1s�fL�*$�\�^%Gĺ�y���50����l�"�N�A<s+8W�$`�o��y�VԄ����L��&��C߀����O�x��F����F��M���o��2=G��7�_E͑d$ŏ�H�m{�Gn��~˾�V��%�r��rk|l=VB�F���I�=ո��VoX:�9�|&�6�3�3�9u^)�H�5��w�Ps��I��8T�	�A�q����!���"7UU� �o��QH���ǣis��K!8���Rw���	4X�铌��9�������"�q"����m�9���>�\���I%��3����I��i&�B��r8V�fpQ7�Bb�Y`��ǯ�ۦټ�9Kl\�(�	bآ���,��*�Ō�J���ϙ�_�q���{<�K������6� v1r?�����Ӱ��e���
�j�����yS����&m�{;<�������V.�>��:��ϛ�M��::1��{����!��� dSh���k��&��(Ɖ�
�]:!��墜�VU�)�v\`��3�2�mZO��� ):��VG:-���5d�yN{���Q{��k��B_}������\D2y&��FzaL�L��|E�L5ј�hC��������5��_aj+��w?�rU��� �V<iU�.{��( hWD�h6����%�&f-G'�r ԰nVy�Yl���}���r��������	�C!��Rw�	!���H���G�k�	I���I�Tؠ�`��������N�����3ޥ����l�s�, ZX7N�FV�p^�I�<[E�w�HB��]C!�o�^����<����:!-�K�N�-{���u�~=y���U5`�����2E�3����!��p细�f�⻂��#���v�{YZ;�!E�IkF�n<����h����y��=:�iN�NUE�VV�O@]Ry�,2O�Wޡv�mո�%1ԭ�" ��B���y�2���yu��ueJ����??�m8����fsȄM�j�v�}��N��۳G�&?��i� �R�H�W+nX��av�xqfX:�a�����ȗ%�߹����td�Ϊr�wOQ7�Â �#�p}�	��=g�IM7�ט4Ѝ|T^v���P<3$/�f�k5^X�"��w�Z��Lں�?��U?@�
D�4s���)�)��m��=ӛ_ �t��Yvl���/TX���.�D-;���=}R�gGw�YQ�E,�0�C�E�`n��OC��eII ���j:2|��}�U&�i�zJ�y��c)�i��>���=V�D�R4�'�
��4�
��H`)gָ��(N��ҧ�(�X6��)�K�`�vڜ,�s(ge��'��;���=���r�C���T)����0�HL�k������d��9b��,/�.��ng[���8b���5.�DL�{���Ǐ��̗;�l��3��$V̚4'-��(V�Dġ����[�2$�n��U�p'��$��!����6��m�v=3@�5G3�k�i��I�9�~s��P5}���lv�
���s�q���c� � .I63@^���:} T���%i2[��˘	yX��\��l}�L���]�T��ȱ��"a����h����V�9�M� �BkRJ��.�̀/mEs��#�n�*��7{�̱vIP3��/ ˕1۾v}1��F]U%�m.2<��&��h���\V���5��8�؊���>
X�q|a<�;߮�W��X�k�|h��Y�r�dߙ�9y��K�WT��~� ��۠�Uğ_+�h ����WfmB�?��O�@��b?��t�LCEj��k^ȶ0�(�~x����h���Ov���~cm��R���wߩ��Q��~^x����fшe���"R���J�OZ%au�c>��'i4(�?R�
[W�Po@�Wt�*fS�Gce�es���`މ
-�l�q����U�ˠ�tt�n�$��TՀ �BD$0���z����C��%{�X� ܞc�����?@�z*:�w>w����`�+R��F5لQ�o�����W���<U.H������B6�Gϯ'Ek�x��>g)�["%�0��b�0�k�jA�1�?�P�_N�Fl�W!�/Uh��<���v�,t�4�œE{��ٛ������h�V�i��¾	��H�� Akn�E;���������\y�=����*mU�%0w��|�ERq��U���[�f��}}�����V1��J�X�9��g�Z)h�ShYo��3و+���3O�oU��aT��P�>c,�Ց�'�Þ���fyjG�<�htp���-����D�:q#��q9(V���B�t<��H4��xU:9�ɔ�JhR����vK�Ɂa��N,�^���4}��7?�Cf|Uہ<����b��Cw�K �>z8Qh����|yԩ-�V���(q�Ɖ9��X<%�keD�G6Y�(��e]F���q$֔Bߡt�!�8ʙ�>��+�QyR(� 20o;�p`_���i�Jzr�+9�F��de��
�؏[���������{e��K���'
��-� �%^��G��_��?��cz�k�^%Ш�5G�<�����:=F�������{��R��ɻ$t|]��P����:^PR+�V�X>�,�ŌAJ�1hU��	y(%`e�nU��v@�Ҧ(�ܼ��CflH=6]����/�$�QO�����V!R�������[&�{�Jh�Ƥ�LE�Phw��������7��qyGn��
��'�k	qְ���v�@�`i�?"��6Pu<Q2ȴ(�͝ws�3��`�<��"�p��9`��:����C��Xت4`�I�M(�Hвe.�l�۪����o����z����S�rz��a�f����1;��𜱨�c��dԖ�r�U���[œ�K�=��k��9��%p�E݀hr�%S�Ѵ���^�0~a�`CX�ԃV�/Ren��I%3�7�e����<7(j��3~p.��$T$�5�X�������@��	oa1-�o��?�y2�v�(�^�%�ַ���`��~z����PJ��E��9|���7�m��BF�/��َ����3`?9�ͽ�ȨQ΂��XS�� ������"�[�i��O�$M�"L�5�� %�Q���W9�ݻ~v�wr� f���8ۑ�Ҁ�;x����L��r��n��u(�K�B���������|�>Z�(����O����)T�+f���:6q'�����AϾ~d4�X70O�^���WR/-w5�^Tn������k\M��,PI��w����y������˪.hp4Vd}(N ���:e�v�'mQO,~�b�����?@����34����qĤ�Zy|�<U6�09�DmF1���B;N�5	 �A뙍&�A '�hs9aT���B ��]�����n?)��v�c'��@��}����8L���]Oi��Ŷ�]�4Eh�Ɲ6e�#PF���̷]u������?��|E�6�X>j��?�
�{)�8+��4���-�kղ���\a�/}����&����.�CU$D;��S38H]w�8{{����6vU���ع?�TsTȽZ��䂗U�&/�I�0�Z@���+ F?�h���%j6��Ta�L�ʽb�d4�[K~���d��7nw�W1nW����)��16
�K��qi�k���5�v�e������:�q��#���Uu �RC@)�P�3��c�h�:�XA�8���2�I�7Xb�?�Ҳ�5Jg�����T�-Ȥ�<m�B�9�ǽ>���-���g����|����iG8$���z���y���b�L1ӎJT�|���:����(9l�p��"�	���Y�����H'���ZuYϫ�@K<���
P/�
>�Urh��?NKb/# �v(���x�L��c8z����n�G=\����C��E�0�Ix/V�i���c�����)o�&��z�48i9�bE5��z�b��,��' ��n���dR���V3�ԏU�u�V�_��A�e���PA` �ʒEoC���(l|�x���#��\����}��B2܊C]n	'A�����É���s�3�e�����L�i�� �:P��V�uڅ�� �����hc0{)[t e.�iJ����:�˾���V�
(%�#K/��qek�0������ �'�/#OaSe�.M��W���A�[N������F}�����JɊ,D�5�
��p���^%��W�C�ݛ���	p�N-�)
�X;ʦbSu����K��i��J�v{�o�7ͬ�v��EL��?��_���PJ%̋��j�xf��%j�#�Y$�񻮛��Z�V�Lkh��:��j��>r�(�/k���R�Dg���.괠�? �}�?�S������u��7$���4��B�p�DZ�{���.v�$b�8�%W�t2lR��X�F0��TT�8L��wT�	�L'��Y~vi�e����#�<2[�+�����`��z��G��yMD���0�l	9u��I������|'��fʢ�H��\�X��\*�a�_�󪝧T�'+�R.#��:p^�{jCl��{�"8z�z1{�
�w���,s1����8"jXK¹��9����%2�)�4Z2[A�74���e�[����Y��tJe�\��.�t���_�j���41ѹ`m崉��2��ߐ7��s
}sm����˥iГ�c{��wW��/��]� ���z���˵��`R��_|����>j�a��7����8+��n)�>���4CWL��;��l�Ve����YC(��3��WI�j�L�ٹXECS�C�5r�%OG���%&&�>:��$����޵���&����sҁmi� �����Vyf�����h��=��#b,����4ޘKk ��ǣ��1�9T������Ǵ����)�����,�������F.!�����}G;�Q�v����d=x��?�Ā�n,:5�",Կ
���j����8S5�8ݔ�w��/Y�pVy�'|���E����2h:kZ_ODlA�pCTV"2v4$�*�����k6��yE��i���ҭ�"y��Gb�J�wݜ��sK+:�*�a�����8fL��Dac���o�g�����{��~f��1c��ӯ�����3Ry���AE�uk�+��ӢMN�p�LOs��=0A�@`��SƁ,�D;���ViSE%t�(Bt�,Y��p���Л2�pC��<��X%�`��P��4�V�f፽�YVA~�����%"u����.]�����/���u�����[9�Uq=�GJTޓ�VB"7|������y��S��nX�z��?��G��a��!_kĎ��&��ᤰ�t6u���ЮO>bv�V�Y²�P��o�w�3{
0�����mb��S��
vl�g}����?E����p\K��>�����m���Zݝ�e�pmN2Q7��fp�8��16�`^��;rM�y�w�$��>I����_�7���nH���ץ�o�^�3�@S���Iht�[���i��~/R�Ɉ+�l�i3�ԝ����	�j�3�Bd��4�@����v��7���gqi1#��A�E�r���pd�%,�
�}���NJC[_>���{�"�U�iplg�J�U m�֩�-'�ˠO/��Ϟ��C���)�t��w�;ɏ��O.�pvSiHxa{���%�go���)���djB�3���|hm��`��?ڴ�9�`^���{�XE��W���v��yI s�T�O�?������/"�ߵ�7�.9��Z^h;�4��̯�n�P�l�hٶrcȳi��3�#�������c�d��IR��8����0\!�W���K�V
�{\TBO &�<lPY�Y�!/3� ͼ��%�E�=jS�Q����ϥ�$�폍�1�"1��%n#����A��V��'�����17� K��@�)=)4���x�ԕ�|V��=.V���X�^����(È��{�9�ȋ��"W��,� %т��."+_6X�h�$���i��nq��5�<�����
1���գ���R��!�H�y� 2��ʎ`�2h������"?���c{�ؿ#;�����贒�'k�z����¾Y6������s1�>Fܩ��(RӘ{���"�0�+�""��GE�۰��T�r�|�sĐɸ��"-��m%�Ơ4�k�/�ɱ�~��'d��%ch<�1d
��:�o[���|�rj9ŀ .4$�9h�SsC�أX�%va��?M�pwyF!y2�wtGx 4]�p��,�$��Wv��� �'�ל{4��hL��tL����Z+�f��fa�6���Ї� �!��5�UƤ����^��#iSn�.u���d�]j�������Ў�J��P�GF:v����C�L��z�.�8S�hп(PRm�� �Fҹ� 4t|�H���b?gT���۾�=����4D��e=(Izo�ޙ������?T��o_-1���+�%j��G��+���x�SJ-�� ]������+�0�W^F�����c�?1F�&K�`������}�߾N�i,�;O�C[��M$�D�ưM�)� �<�m�X�DY�ޫt�<�06>Px4q�]���4rf�2DD;����TabU~����f�yT�E�I��#��#S�7KQ�[�@�mGR�)�sK-s�\��\Ii��؇��St�������w� H?Gg��W~��r���{>gN�U�i���8"ڨG� @���Z͸��2�*	X��-*�D
Q܆�﯊Y���������1��";L�|���3�@|���9;lbq�ϋ&�����.�=G� H_g|��@��08��b�3��^^z�O�S����8��B��i�0�5Q�>����������b��9��.��y��<�*HX�!%��>I�md���NiI�b�~�Yh"����Y����,Э�<�:��%x�&���h�ofC��(]���HK�SYL�B��iW�,�މ�~�p��� 2� �k�����d�G����3�\M�q�̗��U��^��,"��W��5�$j5�x+Ϋ�(�^]"�iIW��Ni�j��E�o��^!����3�\�=�u��
[L��z��v�c�I����ڠ�h#VZ���������ԇ��,ۮ�d{�t5A¢�魓�DNX��g�ӦE������YՅ���W�It���y�z��q��l���u�Ղ���Be�І�ЦK>��G�M� ��xغ�d�i�����	{»���Y:��aKd8��"-���g2f��. ͻ>��"����������Fn�jʹ�t-���\�mE�mؐ'3�50����OÓ$���|^�ګW�~�DGz�T��E��(�4�g�p���uk���m�ɩfb$;��y���d��s��B�a�X��&"�����ӃrM��#mK��B'N�h�i&+&��(�������3�ੰPyRj��k!�ӟC&�ņ��-��Fw��1*�T���O����[d�3�<�8^L~�2<~h�,�C�6=�6+�S-k�D�W����mB�z��7�N�vsV�`�ψސ���Mly�Y�yT=IlW��Qt�H�1�!$.<$�fZ޸꩛�b��
S7t%m^�%_\�|p�DN�A6�ou\��G����>�{�E���tYB_��S���r��@�����D���ǥp5W�5X��֓"�Sʔ������Z��_ߠT5�K��\�Q�����5`�|��U���-&����cԕ����u�Y���!�y$�<�����Л1�`oqv�vO�R>�:d`�c�K�M�9���5 �cz��=�W%���eZ�_���I�{c�&D���޽���+Hm��9���R�繿XeL�Y��.���c@:%��	�������!t[�Z�����і8���2���Ȁ�W,Q@Bhr��><�5�S�U[�x%�y^Bڔ:����]y	���!UA�wA�f��eU̱H/x+Q ��} L����S|���Է�/��j�l� �c��Hւb�X��EQB�V�T.<�Y�9����cì^HѩF�=�ȰL��ϱE]5�W�+R���٨�p�ʳ2l�
�U�UcbPzf+�ճ��Q��+����>�A��Cpa���q�J
�q( 4��VL.� ����F̯����Ч�(��-x���6gR]O�L����, �T��� mÚYp��v,$�}ʸ�J�0a�䘞�|E��8V���eǀ��s�K�oE�U/:?��r�d��z#���lP����վ�Ї���P�o�?�$O%4
�t�Fn\�,%�Sz�w�N�
��N�M��~�ya���%�w�'s#jpzaD�iazC�z��_���D7�Jy��ɶ1�Ë{��j�&q�W�b�-�v�V� ��m�
۵��HbZ6��@�sh��ű�l�L�{[Svh# �i��g��!G��#�6t���x�������=s3�>��@&�d�!�B(|˃.Ѝ��%-�i)��!%`8��'��K�*�)Į��A����]����d�{7D�=�^+�5�4��Þ�d	�j�d����.�*/+�%k�6?E`\��(wGBqJUU:fָ�̓�=c6;r$�J���r�Ԭ�����˨�R/n��P�(�����\	;�v;�j��o �����g1z��aÐ���"'��`�:;���s-�g=x��p�5�:�X᧹'z��{��4�_G)���Z�ur�ݠ�gC�"Z66T��>��D5�˱�7 ���'�۪�b|���L�e��[����j����~ڒ݈)����������E�5��SF��@ ;��)~�˫莕��{�{+C��Lo�GA����c����0�Q�A�ԥ)l�2�����湥+�<�w�^�m��<���>��c����ǻ�W�An��b�y��x��J�Qu,�X���� XW��b��������%p�p�KQ��N
�D�CW�Bm�x�e8�^<���BJ�ӑ��+tJ�;��a�s
ӯh�����s�<ݾ��=��E��X���a�Q�%^9�v�Fy�����pZ�&]c��{*cl��w�'ſ�t�����@x���Q�K�mvTv����KM�7���g4��&�FUf����+_�$�����l�M%v��$��V�iv� ��M�H5���b������50�cNIlW�S,�����_�hDIS�7�̺RS9#���N'����B�KAw1��$;!!P�.�T0�����_��P�-]�Uz�J������k89o�xw��
�]Ҝ�<(#z3��ّ���t� �%�gU�x�KK��5Wv7��<u�2�_{I|�ؚ��m
ӿ�^�Q�<��ݸj���_���� -�1d�s�P �S��ѐ���[��:�plx��2�D�%9R3l����͟��H9����8��bqhz���s}�wfsH�]�ę/�҇P�""�X*S1@���7	Ei���T�1�S}�q�D��^D�^�J)���g�����F5LTE<>� }j�K���)�@cō��!Z�H9�TW� &N��UM������,b��12�1/WL�%8ƬŁ$t��Zf��¤$B�C�v�}��
�@��tj��/K:Y�m�"�q���o3�g�L}�J�4\�T5��ZHP؆�H@~g�ɻ�Ao�[�}
3T��	f'�kq�m�d+/&]���}����e`qqq�!"���S�&�γ���3����d�߈+�)N��|�e%�@#|E��Y�m����ꝙ	Be���#:]��e˙�k���B��=9����¹�'�q%�y��w�� �$y�W�6����v*��l�D��Y��b�7�T��p��wn���D*}�uβ����!�5��6�b��F7-�RsQ��Ǟ��y�i��J����)��߬�|d�;��W�'�,��C������L�k��&���UvMn��{��̽M'`F����*z�D�@~�%B|Q�"O���
�N�잃����|VM]�3���J�U09w�������v�<��T��vXi{;�	>9���a���k�Ѵ�eOh=-�����2OU�Ā��T:PJ�D!�?��|^}h��	��
v�.K%U����E�3y�x&<���Q��$�e��İI8����?!`�6.{76���-Wn.ǽ�x��S+���S���H/�T���ӑ�e����w%!��B������
��vL {'����D���P����Φ���i��s#V�r�b����@d�G�5(������c-��l����N]�_\����C��>�:�^b:~2m�U��������ު��2��pǮsc�lĈ3#�8�z��h>al��k�t$϶���?ys�����Z�`.6�'��c�N(�8�4TG_����~�~~�0��Ճ�z���A�`#�w �fg�6ri��td�\�<X>1�&��^��#��4���-h�I��y��؇h��[�o*�/9� 8�
��^=���J�foz\P�	XjD�7��=Q��P��tg˃Q:t�Q��
���u����$A�\�G��T
���nR;�>�� LwZ�tl��{�m�ĬFdT�P<����|�b�o�|A��>��ҦR=���H*<�r#�Bx��Z�}E^ϔ�\�/-�} ~1�^����rnuBӲ~�G:�����F�@��#Z6)!b�訑(���VSIz�E8���*��G��Z_*߯���u������ˏ_\,��+�2/�;��3p�.��6H5�di���:�<��
S��mʵ�z�l#��ٞ#!yu��p��|qT]t~�ߘ��Da�0Kkr���� U=��L��e�K�r��a���bC��mcS������k����:	&�d����dp�"?c]E��ptb����Tr����=�¢�7s�uXp)�Ys�BѨ9~�i ����8F]<�q�t�t+mNT������zM��ε ?���l�d_��UgG44�8�@�hn'�|fU��n�>ȫ�&�Ƙ��j�>G��{|���e&�Nt���g��r�AK�T�!k����H�H�oW�YTiƞ�=
���;'ZW{�A�jKI��h�`Tkfaz�1��瓢U�-C2��
f�lm��A&E���w��䚚K8���wg/2r(�'X��BہmNR@jY5��?�Ȓ�w��d=wF�uU���D���s~�Ǹ��^
Q��OL~sOH���$�2K�p^ܴ�;a��t���,k��Ni���!��s��>���z'���%M��Ae���8E��[�����TM�S���Pe%�%�_ou���+$��}ԉ�d�[��QE����E� ��~1i��"��~�4�t�v⯟y��� 9E�Aݙې����Q륾�v:)��0�)BrM�����8�IP����xօ��~H��?��UOQ�%�'x"��w�|���Ut��6�O���ࣽ����x��{w��0�`�������g�K3������1��d�f�G�g��*���s��m��)C����c�7p����@����ހ!$��}5���z��A�����E�lwvM��`K����xi_�S���z����F��K�ĭ0�r�t���fJ�o�ʜ�e�g��?F�N��5��z����
��L��m�?N�L�]C�V�����]�>�x��o�d@5���-u��%���4�����曇����v>^2T6(P�,hx�t��նM�:bz��'�����j�*�:��w�޲x)w�K.'q��`�5�i�#��z�Rf=Gi�l���b��{:��A�����t�$c�w0V ,��,�s�J�6	�.*���!f��T9ŊDa��w����k�����|�@]لa�Cʉ��"��r��ʠ�S �}���ejeu��6a�g��������ui���ݑѮEUj�\��F`~�C"��q���M'��$�Y��w�8�T�*�����X�n����^���2`m9�t���s8���S��ݡ�B��|ڀ��H.�2��-���
��9���7�H^�� Kok�=a�f��z[֝���Sk&�n�*NU3)���1I�;���&��{�;���M+�'����&�r��Н���}%��l�~�� v����=ן���������^ �c�~-���xzvf�뱟׼e)	2F���̖��ܒ�hw�4,��}H�Ⱦ�u�0�WY?*���-𭂩�1��в|�wi��w{�}!��wQ`��w�<Q��+��Z��������=A��93��
�s9���ayW7�e�����E��*���I\`�[K~es�K��OЅ!E�e�����,]8���g�Y,XJUքT8��V	�	�Yb����Ҏ� <;�g�Ks�j��3���)��7��
��ԄU5�����:,� x��Ix��������t��A��������k���p�xO�e|��[j-C��E�vS���(�X�af�홸�U~�b��~�rLV�{�uq�2ܕ��&����S��NVp�)���������{
���;J�[_D��v5��0\���N�K�6{!�M@=M����t�X5���6 �+~ t�(tgs��0A3k�v�[��#=�Q�\�őj�[���m&��D���!�ᄉ�������V�m�Bv�yt�� 2�߹'8YW�dd��kfV�WV��_��Z�o�H;�|��2�p�p��A�T�*�����x��4�wF��mIͭ�i�+��r�O�	и���:Ͱ�yg�K#��v�~@�h�)�%�\��]bخ�"[`~�}��[5/����(�¤����/Cؽ��]4���yRb�{;�yz����T��)9X�a��_m�A���9.�G�Rz�	�;�å�.9���07��-��yR� �R?үT}6�F��S (���4tb�9�;���6iRNi��E�T�1˙9<G�����$�9S�?y��S<�=����>� (��#R�`�
(� }mn@ЂA�S�ܱ%�*J�ܙy�>�0I���Eg�,��|2�.|Za�w����$�g�.�Ie���c�x�*�/���y�W7�O����ꡢB�#c6�S��:�3��*��6i��4P	��ɖ͠(�7��Fcg��2qfx$�|�Ļ�������˖��[U,\N�6PS�R8�HJכ u�g�D����n��Vs~/V���v0�A?D
y�v$
�UM�R.��5��5[�|��m�4�C�E:*r���9�Ht�H�>��DT�����i�L�?�aMtLK$�)wn���%��w��m�Mn��47� G���Sc�f��}�0�ȑ B�'��.$`>@ Rۄ9dG��x�y�������xy��Iz_V�߂И�X��=�:Z��|�ײk�*��bu�t٥�m������c��>]�G����"\�'��F��`�7>�Ծ�8�cN�����зt�ӟO�h7�����j#e��_�w�����i���3��6��.兲�i�����<� 4v� I�O���ȏl	BQ�O4��X�!I��Cι���&y�9����*&T�l�D^)��鱛q$���m?��Q���T������ɕ��5v�׎�{Nƥ�wK��I	�=erY��(��z�[��$��񆗠�w��gd"�Z���n�6�S�!���ap���"�?XطI�j�զ!z��HaN���(�I#c��tӟ;������9�WZ�34����[�Կ
�O�+َa�,��
�c�0\��"�'[#1^@k��r�@�^�1��W��������
ဧٯZ���I���#6iWtߴ?\��I*?<q�k�[A
xaAy����F�+�h��,�.��������z�\Ќ,�&�ҟD���i�Q���*x�V�����Ee2�O��+X�$uj/��D=�&J���.{6b�]���x��������θx�������� 	A*�+_��J��"Q`�t����j���U%�����m���O�q��v�#/e�	��2qw��A����ه����@��L	ժH��-�
)�#�*r �:y7�դbb�n/�2�����u��PÖn�S���' �����(Ը�o��K��+��_f����H�na��;TC�F'i�a|��f�TF4yR���w�
+�_RKL~y̺�60��xy�!�ɤ�����U��aK�u�xw�(�ܖA���Y����w�U7��͜+␅�2�r�]�l `q�� ��X�-k�L��B	R�`����Pq��"z,��%�[ ��6�6��Z���������c!�;�ϝ+[ը ̼\�\)8�7�Q�K�!�R�BHwsDi�SԦw�j�$rQ��7��*�	"�%&�V����:�6ԙ�_�?"����g�yu�-$����g�:%S�g3��z��!/��e�J�ǝ����wL-��Bn�ҍ|vl�@�itE8cޒ�:����q�#�����Ϡ|�	��-K�0��Ӷ˲>|�*��o3������F ��:�į�q���+oA]�%[>2�A���O�!��s�&�L�����p��0�A~ش�A������&�ܲk�إ�)�f��|��}I�̱��*
X���/�7�n͵���mz�	�_ ��S��%B,�`j�]$������j�od�,��͈��@"~�g9(���������7�m/^V�4��V�?���i�P�����?im\)�'$}�q	H�z]u��f+���4��[��c�%"ԏ��J 缺�S�jv��5�/����M�h��-Y�\1���e�\]����7z���U���e�=�il�ha������y~����
�`���F U�l�S&b�ؘ^z����;���@D�"@j����Ej'@�E�yX����@f^���K���aDV�����y�F�=U� �oϤ���{�xe!�Q7������=L%��^Ƕ���5��u�b��g��dGZ;�WK�l�
�ڲ7s���s]�(�5����-�x��]�ע���N^�j�q�(
`Z��)�N��Fе�����X�������0R�D��:�3����l���+'ʫMV�ŧ�K�T=^ߞ7���*���0&i�)z$�Yv�XSm*1W�1�� |Iq�T��!4��nK����0Hx����C��Y��/S.��=��w3��v4t³�޸z�%������N{���UV�r��q��4h��ⲇzi��Hި#�Rx��E�xl3f�*
�Q�{t��'M�V���C@�з6�����u���v������;K���4�y�xA{Ib�!
]��x_;�����gKB���\U!�տ`4���e/�����C'f������ڣ���#%%���S�n;���q+Y���Ӂ#��|������V;HIpyMl>�������b;O���F�j�Βŷ[�fptB��T��Al����La�:��1MLӶ�-�w�	���\��Q��ͣքw��[�8�Q3��p{�@"�X=V�p'Ic��x�Wú��[)L���*�Kv�X���/��۠M?����������֌�p�ܩYݦɳM`ϻ=��~��t����������1�]�s��8kgR{��~h�T��p���׸�4p.w��������x_��k72�=��̸�Y.��=������g���Zȗ�m������QRGo��_�!"�&����$w;Fx��=�L	%�p�RJ$MM�74��>~��~'�Q��Å!�����h�]P�57��"���VhOk+�q!'`V»n�tǃLu����x�w$����A�j��䋇���fq�q�J���.E���b@4,A�M�9AJ�*/\��yr�#�r����צ����5H� �F�(|P�`�h�,li�:HAwZA�'��(E�D��=�/�J��CŁř`�*D<*p�v�mj�gD>..*y�.�hO�!��߅Y��'��m�Z ��v��5�|W��]3�2��t۰�8K�W�|2��"�Ǚ�sB�a�BvJ�ٔekq����|X�-��6{�f{j�KJ�S��}T�32��x�ډoT!qQ��H����<ãL��i�'!��ŖC-����@�u}��i1N���Ks!�4��;&��ˇ��rR,�/fg��L��|�5���՗���Wn�mժ>�U:u���aò��X��#cQ��yvb�`��E��_q�<��w
�?���j���b«���<q�&�
{��ߏ�,3'��%Uc|���ɨ��<��p�-m�d��Qh^k��ԸX�'�֘A�+��� 4��۞ ,0�L��C�L˴2)�ks�O'/�|'=}[�*��T|i��l��_BDzί��L������2	@���.`ˀb�t��ʋl�Z�$fp�$%��a��A���|Aw�SWD�x�r9՗'�\�̋��`=~��*z�MrY���P�7�) ���Z9Y���hS�����U���Yɍ��\X���(�iT�)��vvݺz��Y�O�.$�Ї�td����W���0,��)���;�}��Ӹ_���ߩ���DL��}��{�+���ӹK��`A$�˖\�GhA�A�B��m��s�Ԍd؟�(%@�SAMz��S'�&*
���9�l����HK1A�Q�$z��*L[f�u���Wt�֠x��k�?�?������G'Xu*�*Qq:�0c��si,�LE(X��en'��j�sA�x%gV� p	��"cɺ�=�uz�)jr$J����^�d�-#+�G�:ƃ.z�Z�GcqE�L]ES;�<weY.'o��=r�}��h�-'B(:��WK�9F"� ����h��ܱ��59��S�(i/#������T���(�(��#����W5���H"=�+��2���1ȇ��}���z?z���Q���_$ ����?ɊM�U|��T�h4B�u�����s��ܐ;h��,���nf�+'J�ĥ����17�l�b�G��\�m��3B�5$��%��(<ҧ�5r�jB!���o;�������;�%
�43�n��:==���O�T����r�Fa�$�Vc�iAF���`I�J�#�?�}��5	�ÎIY��Ȧg[jbc;�pQ��B�����;*�݇6�=O٨���ݞ:�E@s3|�(΅tH���ț�Ԭ����R{���g~��J��	��4��Iͧ_�,4Dɯ����I��t�Ƿ�in�>l#M/���wទ�n��˪��0�o���8T���P������_��\�2���*U�StC�_�8I��W���Є@�ԝl���
HN25�]F�����q-������{z�=���cՉ��"
��f2I<�%|"��{LAQ�����,�qp� ���\Z�mY�����b�"���!?��4@���WAc��r1 l��	��o[�gf�D��R����ݖRk�c��%6%��L"�G�)i��* �4�X�E�{�\XE֨��?��F8�eص5t�
J�6�n1�Q���1� �Q�$��IYt3�$޿�F��#)V\�S�{6���7�Q�e(��n5� ����>���
 �Ɏ�ƧP��i��=�4����E��+ Pޣ�=����3�=ߢ���C_+�	�,u�W�	��d� �[��$F5��o=�1�o��J8I��!���@uiivqj���͔V"�5���M>-��&8�S����[�̪xKY�A5`#sqל"��s�����x�܎%��k�g�]��Ճʻ���>|���n̰~̱�7��S�#��G[*h\�7g`6	[#��U���=����c&�{xl���h+S���C8�£�3�=_�Bv�w�NLnI����e	A<����/�9=@�+�Z�{^���BVf๞�Zz���1Ǭ,�S��{�9PfZw�5S���5'h~��?�o>ʯ�R]�~���8�L�;�ʮDF�>�\���o����9n/�:��S�DshQW�"��h��-�Yo���Oa\8\��������k�2,3K9)�-��X�;���G��|z��.��eY��}�6p�w�������p'���M��y�/��<tS����!'��k�l�jթ҇v��x}	�S>�o�����c�w:��P��BX�	e�	���S����K �Y_�[!��{���[��ԋ(�����yԩ�W��C� }���ioc|֣0f�I�RK�A1EEy1p���_�fvo��<�'�wq�Gx���������ׄ�Q���+A~٤D���Ok:��=��؃���^�N7F1�����|C�ݙa���oL�<�R3���RL9@{���I�[���Ftru����O^̍���򨖍�Wo7�J�aau��AӸaQ;�I�a�Mj Q�w�&eJ~u���-��3[[�I>Ybo�x�$��}6������Ǿ����u
��ߋ����Y��t�}(ד���q�*�A�+�%�խ:Sm͙a�n�S�Y�_�������Xi6u0-� �'�"�LC�����O�L�&�Q�����T��&���/�(�|17l��J����)�0���;)�w��xj��<� J�':��¡\m�8)'�n��|��䦈=_�f�J��R�e���� �c	���ـAkP�$'��[%\�t�I�S���8�	(�?ɮ���&�
�ة�pbe[?oE���@ )P�*��GzM��k��4hX�B����'�#�#�}т��_ h�PF�n)
��\��&
��"�T-*�4G�O�nY���K{�	�JԄ�G�� ���z�}�zvλ5�C��@�p��P�4��ԧ�2a�=��́�&J���D�k�����"c�t<�c�fG1OӺ܆W�za/Ra_�X�p`���o��V�RR�PT�n;f��?����Coۇ>�E�vT�n]1�h��H����[� �_���t0c��_k,l�@�.�<`�����(nF��D�L�g��9�)�7{F��']G�;Z�LD�~�)����jq- #Q��M�!>��U�p�oo_�.E�5d<W��8�-����!P�v��g�m�!��	^�
�p"�;��C ����`��� q�W?�	�=e��*�����Z�R��m3 �v(D��8����RF�U��U���A6"$	�C�[���6}X8��;���prj/ڗ����K�YM�U�3���R���19���}��������$��������Es�x�e-������.2:�~�w0��\Dfג�,Xom�J�E��qϩ��[���z�q��:��,t��E��8c���!�`�
`5:�L�QT�HJ�P�b�V��7�A�fG����2�J|������Å��m?�H׏3k{�M]��J��\�܎�zD��Z,��1Q��2e�r9���X�ce��Y��X(�zI^]O�S�u	_.���ެ���"���B�#���_���Џ�s���޽�$���-?&l"��PD�9P�����
:�����y�9��;�w �4�R1�؝��
	F��Ƞ������f����O[ѥfSwFz�_9�aҿ؂�>����a���*JaaPq�z~�-�:�0����躧W�B��V���a�Q��W|R�������=�����O��}uo W]ӀF��6��X~?��(��$xÏ��a�"�����3��&���؛���fH�xJ6��D�C6�}׏����t���	�ab y(�_�p�x"�j�o@��?���&�P�r���${i5<��ߑ�=�Vݳy��xps��uysS���<�
1Cp�s}�S���y�!X�5m��}��Գ���6���j7ԗ����8��N��@���nn��y�@/ŋ=��"�aGx�.rq��h�y��Ϸl��fP�����V�tr�����β�h�����^\Լ"@���(�9*g&�8%�T�,�M;����SȌ�ԟ���&d��NE�ZLz��K��q*1��,��>F�:=s�m���d9m��vM��'�҃5�f`8"g��s*������aO��Vo�� x��,F�w�W�f��gT�
����ͬ����}���ׂ�5��\�:><��)�r�RѷC-DT�6�~��˃��ƸG�.k/]�'
S�����}bxF��Ս����ISF.1�O�K��f��c'�x&�_�%��NJ�COf��SC:���؆X�~q�AK�)����1�^b�p����h�15��CV����<�_�U�����F�ׂw�����G��|>4�+1��=�D=p��-Z��"��a��gB"������39Q�%
��n7tW�C��d��a�xl�4]p*��G=��q� �6�^�F��Y@�8z/ۼ�O�{�rT�����rl3�W�va�v����5! Y9*zN��2�rܴ#�G���/���т��y�#%l��
/H�?Q�?�9�{R� 8�,�e+ށ<����O�0�~b�a<���O�%I ��UH8=�9G�[ē8������\¾d��ێk[���=�%!���B0?����g��Ӓ ��� ��I��O9�oTe�$^���,�CD$�=r��n@���P� n%Pw>���S�*"~���Lh�xO�D�Ag���2��F��9�υv��|�~���ɗ/�漭2Z�)���Rb?��m�[��:���0���"��o)�*���$M �p ��N�C�_Y�V�6\�$OHCδ��;��4�k9�轕b_����˩��5TJ��szR�պ������x�m�M�6h%�&�O�?tO(J��Z�}΀b�N�T�Eq�-7��{a��A�{��%H~���5��_�������D��><y�tNǺ���`Zw��GS�n�����A���r���r�a�a,ZH���r9�D���Ff����h%11�PhÏlR�
'&����t��������c��U�cF�W����ٍ�VQh�������!�
Pl��?Ν۵ֺx�����,�Y�xF�-�z��^�4z��\�6�hA���k�ۻcW1����0�,�Q���>��V�`h��� SR��t�
���Ǧe���������DP��0ڴ�}@ ��C�j��u�PY;^���E��f4���M��I樹`B9{f=,��>&`��8"��C^-��'c�! ����*��M)���@����U�X��@�A������,�U�T�<� �x�Å(w����`�\���#J.���^��5����j
/��2��g�Y����� FZn�g,j�v�.�`,�]A�߂���찅���[��|�8���]^r��٘�{�ܞ��!'�ǈ�
���=�4�{a�hmG"^��L��]w:2��)�����s�MR@I�H���c��3��0|�x�/)�S�SbQ�8ʩ���'v�$�Fn;�j��$/��&=��a�Z��J��-����$�Ț3�X��;iyה�T覌PD�2����m����%@:�f[��-�A��%��u�S�d�.`k�U��:u�_��d��^����	a�i��W��<dp�w����D���ԢQn��g��������B�f�����p����:R�5?��1#�ʳ�r %��S�����+�o��B�@q�q�s�a�%ii�l�|T,L.�+�KFg���7p��z@o�L%,h@tI7q��}Ξ-�5>�,��z�d�����j0��U�u�'�ZOJ��VS������~���膄,E��i��+�,3)D�$Qn��J�$[��ju<!=|$�n���	� �)fΈ`c�D<xw��1L�[,�Qy���� ݐ�
�ya>�=�PE�%MB禒�;
�)E�b����[�b�Z�Z�Wq>l�gϢ�mV���� �7��I	$X0�� F��!��#A�[v����.�g�!+*qL�_�t'�K��vT��7 ��M���͟[i���[���*xT��s6�*6�z�k��V�y��
�=3�1 ���~{@&�B�e�j8�Zlf���ɥ�� bE������XA�r��a~��~wT��[��'>CSH�v��?�zY\WW�_�,�D���s�1r�6�>b)���F��3;2d���9��!�N��c4b��U�fr�d�m���C$Uv��:�]GW������Շ�N4U�r^C.چ�wAm�?o�,16�P`G����2���N���䀹�Ίr*�c���M�@�#�U�B��p�^�X�1�>���^i���VӶj� �t/'�(_�?�&�� �H�Qa��'é����w\�	 ��Y�����~#�`'�wx�M�~A�y��"`�]ԟ�7jLG���1�CŃ��y��zy�O����G�u)"n��"ݒ{!��Ak��������l�m<�Ҫ�ڹ��?C7?����\���E��zB�)-�J/�F3Θ�'�G ��pCy�wacQF�0��>r��Z᩺-��Е��Zq��T��m�n�ai�5?��i���5��h���[�x7	��,���r4��y���9<%/�d$��7��*�f�f�#�^]�u����':U�?r�?<zZ�~��>i��#�d��W�oz@u9Z�{�|���`P�[�R��d�[ZӺY?q~�r�W:>�צ��2�8����� ����"�N�f����T����l��g�Bv��)��O���}P�t$�4�� fe�{��(F��_0{�B�D��{�spJ�G��H;į��xSP�\�9.�:ޜj��(���c]��2�N
��dQZ3E��vR�F���lOs�Z�F��uX���x�0C�
�")jd�A,����P�������:�n�YoOC]��G�䐞�2���30/������z�:�����茄���3���%<�ٞ�`���ۍV���k}�xǥ�� !w�;^�s�����j��r�{�|��5A���9�6*�3�9�`Nm���F���4�`O��jW}#��ĠlgY��},2�u�􊨫�ӧ��))�>w��v?G���,vg !=\)����Rǡ3v����&�%缎��5�+��ɳ��m:�,�����\ ��ic�[6����������$�n{��U��eX�z�+۞��t���?`T#Ψ�(��!��n1'�6u�g�-[����!���_T���w��xm�E�P�H��:�w����H-N�d��������������1���y��b:MTH���w��<�º�!:�ZZ9�qn�;�gOi����}�^�TX�H���n�6�јTS\J�⃹9?=�!��G�8SRZ�~�3'��8��]o{�����?q���F~�6qE�Ҩ>V�3W|�(�1�6�e8L�y7ů1��W��;`��31X�ӵ)��ָ����x�c_)���,� Xqx:n���>:xs6)���;����d�n~�l	����;f��.����V~��^�p(q�������e{�Xq������Q1Bü?%�)t&��H�liN�,	�?�/d�#��\ 
�F��,���$�|�OH��l�+z�. �H�0K�ZF�o������Ő��,�b��d��qL�_4Ž�lo]#
h��5f���钭P.Ɇ�X���P�ᕘ�H-��oi��r�����qׇ>��XjZ �E�� �M�+��⥾��J���dZE⴮�<���C��,��\ț?�;n��!�*�RS�/w^���u������\�0��G/��߿X�wzE�Ӛ�3�VҜ��g2���(���ϗ��y( �Ӈg��1E��=RM��҂�`�q�� ���ݫ�u�n	i�fRdM��+R(�̻|��D0e�vf�KT5����[�=\�X46��s�ż:�gsTP �{]%��Ů���x����2�J�76&�-ԙw������C� Y���/@8gJ��w{��Y,)k9d�Y��ݮ���&�\� p�9�56��&�O��_��_+�k�����<ܛd$�^��m��g`d������[�J�$?�$Hf��[���-��I���!s��]S��3o"M�ɨ�ӂ4�M��y��l�����2wv���r�`\.)HP���!�Ѧj|���Z�)x^�W�}��#��sk���H��{ո:��6��s�@��H�9$��^�+_�`cK��j�E��g���:ߣ�ټ�#�:�֘?S�\��f�?S]��!�`SH�|���-Fy�OmX��7qJ�a����˴�x4�ޯ+#J�0�k��s�3�I�f��A-�|�	0����m��xO"ϴ;��˃)o�*{O�����fυ�L�Y��m:A<��J�3iS��W ʘ���ۙLD��1��K��ӳiO�?�PM:Y�JJ��$�Oٿs�KxHl�F�xD���uK��o��~�'�y�q����Kv�;S�/?�Rq��L���f<���-��STN��>d�½�	���m�v��r�2���'�cQ����5����{ȶ�Sy@���Yy�&��#[u��]�!>��gp���NV�t��as�Y֭�Xoβ��d�.�"%WW��t4F\K��Oh9�z1|��`���]��f��^����Z���g?_.�l�5�w_���z`3��i�G��&�X��������Dh̍ttăO���F���F�7=�F�2r����o	z��~I�@�H�u}KJ����*a�����]���g�q��T���UQ�D�4id�i��jN�S��c�D�w�w��_�,�qK��y��Hs�����z(�P5Jl�"Gj :��K�~�v�d��R�νZM��UW�X�����ZTa5�������C�o�Aԫ�^M*�C�ϵ�Eˣ�5����ь�"8�S�͟�A$~@r�]��
>*w�u�ok'�Z�γ�_0T�͓[h�����0n��ƶ�	[!R�	2��7�diB��K���ωC��z�!��'�V��R���v�ôU�v��L/=�q�s��ؒ�yʒ�^r��!��fS�K{
���xA�s�%8��"����ط�D������D�I�-�h_hMr3X�xy�晕���뚥c��v����vISb@xt�F~������qWN���=��͢���K� ��'o#XgT��j,:\S�BB1�Ff��ؘ��"�$MY	������R�K�;x|q��!�~���AO*i��\g������=n��6���s�R�/5�qE]@F��6#��6VކL�e���=6�pg�?����D���h���<�4V�L|���R���$?��x���&�\��~���q2%���+�[}]ݜL�ډ<��P�$t�l,e'��ƹ?��s�t��*k��!���hj jeԊC�L��tXKu�aUDz�0�ѿ�����l�-.{����i�E�+��L�,��u
��%k��3dߕ����I�_5��;1"rja���D[�j�zit�5�.�ʏ5�딢�bw��h%]��kE�0���x)^���(�
> fl{���EU���rP���v> .�3]`�'{j��=��A��2�}���AN��9r �e��$yE��#�?UrȘy��Rvg����@ޛ�{4'�$Ї=�����]�M'k������Y4��N�	#H!]L�8~��'>��	���p�7����w�W����p4O� 5���#�i$:3~>��~�:������� �W��fK{%���'�_�$F�M�W7f��
S���8����ZG�#���ĊR}x�<�K���z)���.���Cs��"5s~��x��� D�q�?1�U}2�@�y�h��/Ϟ��w
�ɿ�����#�\�3f���W�@I��B�׍?)&f7r$c;�}\p����j�H:��a2KՊ�b����y����rD���{I�F\Y��i��|�zƠ \�����<s�z��t$��)�$
��/-�����H���g��}��V�-��ԭ'�<�(�GQc'��3���c�aB�nۉY����~�X_
c���M���l�1���K��vFp����d;Q��%a�u�B݅�Q�cSx5Q5����q�<�?�z�v:�Ӫ�b<n9�"�U���Hj^�Ѵ�P9W�v�s*�F���z�`0�C�Z�zK����#_B�����S�R����<���`�,���[*ʦV�$6���?�����x�ӨTH�ٱݖ��)���Q1�*DX����Ѷ ��S{���&�&oAa+L͹��e7������kڵ�Dk�+�8�}��I���#��*f�h�'�˾bwEU�E9[���[�&'�*���m���Wv�l�/�m�+�����A�@-����^M\r	&l�P�'؄�VT��&��.3�-y��~J��iV��X�W]f�4i")࿞o�*K��=�sr�$Dg��xl�d������UfX�e�a`X�)���y���P4'@e�M�,X!�4�j�e�|��Xh����(�e��hF���h�y�U:�'h��#��Y+�N�i[���p�l��*2A�p���l��ɿ�ߒ�%���{�h�����T�%��\��2+p��W��m��Ke>�x0�.i�s21�8���U���b�8$���h@<X�%D�x.���5��"d�ص]��*�_&���= �7S��[`Xs[YÑzi>�&�X�i��rs������~���2��uO/TK�p��(Pk�t���7"�7]"�T�l�&kw�[�&7�B_�E�|~0���.W�HL',���|���55Iנ]e���AhY]0ꈊ���n�W�����MZ�1b~j뢆6��bmdS۰d3����X�_� Q��˽�0�[�X�{i-<�כ�&�0S ��;�ųK����c������	X-� %�����@3I�/�4Ar�`x�=�p$�^ӽN${׬O���Б7��
i)�s3�Q]ZZ��]}��ppZ�&�U�����.9�n~y"���KQsbʩ�ppQ�9w>����N�#DFml�'vl�٭���D��e1��S���@�⣎r"6�>#,x�,�j���BÓ��,`��ȵ�Ujs2M�h�=��K;��=5��5�r�5omȺDog���c�\"m@�bۏc�<�ޔ~hڌ;���R�;)�����c��"3(��}�9�=�S�[^�8�+���lKl��D��i�k_�D�0�;��K6�阎a<��Wg5�k�1i9o�a��M���3`�+�m`��iה���2>??F%��9��l+2�/���s�4dM����z-OW�Q>�N��R�1S�!3ȶ6��tj>�0�\hT�����Z���O�D38G��xz�Y��#�/6�������Mw=-�ܲ#�k�3Q��x��Q��p?.�?����@�0=K��>G{y<$�N�"Ű��PD�vBx�M��O�w>F����T� �����_����&���ϣՍ�'� (>��Y�WP,oYY�2^�m릒�Z�X=6��f5K~�*B7Uu�l�ͪ����O���#���@A��5����1�֪W8��í+�m��DR��278e���Y�H���>�p��ą_����_=�j�x��F��n%"rh��G�A(<c���8�C�	0��Z��
L6��j(�)}T.%�� {C�s��4FL6�0z2L��� °����}������@Cd�;�*�lb)��t	[��&.�U��JH��p<�DS��@���J`2�S����W<8�aEߍr�ŵ##ZikUX�e21Ċ`�zr�l���R��E�m%O�O���X�Aqj?��@ �n�?��|�{f_���ԓ�1�T@ZCyQ�b��!�/�K��Ѳ�m)�<;s�ʹ@$;կ%f�� @mKgu}>�d&��L����ɣx�&T�a�^�pCͷ��J��u���I[��l�E�H���nｃ�ˑ�T����"�rgV8��۳1H�82��bT��@��|��}�R�����|';*f�cd���b�:����$������w�"��e�Ph>�G�2��ɒ?"���R@��#��W8���h�hq=�ª��l����\��U��q�ag�ހ���nu*�L��g���_A���a�,�3Q�+Q7��n�eD�K����R��*���6K���C���̱~~�Т��&j>׋!4奤l���]i�Qq�^�6����n?\���	����W��:D�:w<��1��ʢ�r��
��i�L}EI�>{6hbV>�]c7LVBb�������-W̓�0}Ǳ'ۊ�~>*��Q7��?�2!��\�?����oa0nŸ��ZyO����d1{;�S����3,\�RBz�l���92�V/1+x�c7�t�>���@ ��d%w��쓡�+�G�/��Ě��LY��uB�8r������[g��f��3XŌ`�Y(��/�{S�*'|w�n'���(C���vd�&�2�Ѫ�^�!�[R�;oJ9\͈����3X&c��T��^�m=2�����Ζ��k�h��b��*���83ZL� ��ˁ��SǄ+0�����u�cߑ���Zf$�݂��O���c2<b{�a���H@<n���\.��r�~�|d8\ؠY �/.w��� U���J�|��j�C�W���d
~�8�
yt��L�Rr���R��]�46GZ(�8a8MC����Z(m)Y����]~!E#]V,�#��3݈�ĬNq�A�߮^�K0����u~� �n�x�dەj�Q3N�p7���$���NJq��6
��y�v��w3�����^CeYe�'!�9.Z����TF|;ror4[��z��N�wQ�ǀA��"�u.�E�7׿qTW2
=�%O�/o���ܻ|�*]��bI��,����};���`W|k)�]��0h��,�=3�h�����Y���-��n��h�:Y�{�-�L1��O�xp(�y�Q�Ǯ�������yS�V����N�A��?�e�d�_D�3i��T��T�=@�NF#��S�\�O�y`d	��gE�*T��)�.Y!���Y|�Rg{�u1�q���-|Y��^*�)t��ޅn�Fx��o3&�s��A� ce�1����`�K�]P���v�Y����v�jˑ�؋�o#���Y+���{����iU=Sb�L]Q���Ú��DP[��Y�i���Vڸ�o'Q����F�0h��V�VZ.��'��#5g4�V�|�oa�,�	n@�Y+��5w�,e��'1_]:��J��bF����AW
��ٷ�Ƴ=(5��)#� ��y%�}��'��$Q��@K�O4ʕu�5�[��eq:��߸FR�-��^�I�JH��X�z`��F@~^IGE?�=�hw�� ��!��Z�������@�C�x�������9�Ay���_8Ĳ^Je�8P]�Y�c�.��h�{n7ǂU⍰|n�_3���}�E�z�S�O2׺[8�|�y�p��c�O�h���}D>�0�GxF��.�z��l7i��&��]3���w�^��u�{���r�Tʩ:���;X��Z϶�;����9�{�]h����xLZ��=��'ku�1*��]*��YUZ߲zɏ�
��p�s�@�La? ;�b��������g8�Ub�0E-�R�����_�zk���{�$��`���~�oh!�WL��-s߷��k���~L�³�@��d�lW�Q�Э�+aKqT��4V
�����9�J�ޅ>48t��@�+_��غ�M�u����3�-����e#��qǑr���("�����yH�G�@����GY���Pg:�{����~#�y�5�443���1}}U@�c�n��[��WMO('/��+�T��M��C�d�q���:c�ׄP01�~Q��%M�zK7�BOEJ��qu	�����qT�\�tc2}q0!�[�n��k��i�ۊv���JJ��V�/��?3��ر�wd̓e�_u���^qB�o� �$jV����7�x�xs�ҋG���w�D�t���ҟ�Q����|��1~w�S�)��а;����l!�Ь�]��i{��[&},KGY?R�2���3����k$P��4��)䥓pjp�v���v]��F���y)��5B��E˿Quo�S�`c�!-��B��ѯ����ms�>�S�\�L�$A~|g6�jMH'v_l��'�T�^����/Q_q�w�f{a&�6��I��ld�Mԗ�J,Y�>Q�d��ni�"��L�6����	]�o&fT=�Ep"����{?|/!$M͚��/5�����)�4 ()��I^���b!�K�>6��B
�0tE� ?�Y�y�D���Ԛ#x�����ݏ��b��^���x�������l��U"�~����m8��mË�l�\�3,�*/J�b��xDpR�b-+]����l� "F=���*ѓ��h��؍i]�Ǔ��MB�'Tz��=3�����ls��PpڵS���#[���8��X��K�ѯ{�b���ʰ���s���I��)��,�6�������A4�+�m$ፊJ����������r���4�)LcuCҚ5l3Y����|`�;wJ'&�L�uk9Zjٗ�g���EҞW䯐��_����tmB�J��;��zf�b-�R�um���i��f�) 64�[�8��W��K�nu^�$J����;�S<F�/�S���������D��d�L�/3�d���n����&��v��Ȗ˂"�ËsH]���rb��8��~Y`ϔ����Md����^��8���ԭ_��Rp�Dj�ͱ�>�e	Z]{���K���H�U���Э�O�j���~��5W�T���EqG��f���葽pP�$��i��O?�f#�}|�[�����6e� �x�����ۧ,,��KέQL��%8��Ʌ��fAR@
գv�8J1Ntk#��(��s�蚊wV ���]��]`�Z���։�� �Q�̀��9�\L��S���Iu��rx\Z�'ΡT E_���枙qh�[r{��cXa�ż?t����3����$����Q� ��R�	�ۯ��$�>蝱�DQf}�j�M�X/�-S��wW�_M��ۤ7�A��46OH����,�� *��(v��x�8�X������E\��{<�����.+�ۦ�P�8�u��G0�|��;��@Ђ쮉���>�/1����J�!-5dy�8�\�5�
o���T�=�c��R%o?Is�>@8�z��>F眲b��b�X'|_	}�l���RR~^d�Z���}v� #1���}���j#��T�	+č�`�^ؑ���-��A�\qS��_��IH�����u/v����O�Q� 8E��gw¤�O�-��~F��������c�H|qds�]8�����J�K�6?�š?���E ������W��dzOo��m��e�D�;���2.���,D��t��1���~�}�il�L<>�^��kȑp�=p��u��/���~n���:&/��{�>�Z�p�3-���?�ú@���f�A��8y�q�@����H'��@��a%)͝��/2�ܪ�3��ؓ�P�[���N�P���Yi�c3!��Wn�7����2�B3U��>�<��*���9��kq��Gi%xBԟ8�� ���χR����*�nv���	�c_#�$(�-����+�5��8�BPǡ�H6�O�I��F���6�͝���Pa�9�����_xbYY��2��j���F*�>ի2*T���_4����v�:T�'$D�u�����74pӌ��@�*j����B���H�d�T�%��\ϐ��8���h��.�v�p+�Cp8�L�FˬXz�c���`��_� f��h�gܐM�Nn���;�"x@���~���\�~E�t�m�����d<ad���u�'bj���(��BH�A��?#�N�z�Ɍ�ݖ�d�g�`��,_%�:��t�ҷ[�cJ
��� Cy^�KZ^o!ĺ�q��36���;7Y/�-�Ni�*�fE��A&��Rb�e���1=}��|�Q����U�.�<�Á���(M��V��N-�`S¶��aU<Ҧ��/�O̲	�Ye+�r�[:4.a�=�AU��2ū��z�<� �D7��*ކ�j�&�0#��߿��t��Ts���<ހ�H=B|�a~R+1� �f��%��G���.�@a�D>n�w��gi�� !�h<��w�ǘh��A|��aI�G��p�v���4�1�A*���\�UJS���t{C�jY�ҁ�aǒ( -���rSbmҀY�gAWJb���b�����p���S���Iߤ܅6l�|s���	]CV���-�#^l]T�N���N15�	mםb��hY�F�2�Àձ�
�<�k8��*{���������G����n\�a����a�pp���:���h��L���D�����G�y�"u8)�*��u�N��t��FK�����l��T��]��W�
�F�_��q�_�߶.��l��	�e���y�ȂG�w�/u:��Q��1�yɰ�Q�!���a���V��mK@R�0�7/KA� �ay?5%<�Zd���ف
�U���r뷷��%A�w@����ۑ��]Kވ�M<��"L���*jxN����vk����ل�e$-7�	��]��9ۗ�� ��q�y��T�ry]K����E�@��KT�.�||R��Ҏ r�J,��"�6�ߩ��� Bx���B����>���C�5��Kc��k��o��U*ݽĻ�Z9$Ǒ�}Mh����d��B��;�~MpBZ��my��9;H*6�ƃǠ���� �K���N�ӄ.�����/�c^����a��PL�u���b|j�d��+J,�"�.*5|}��Q��{�n�l$�`���M�V�I ��GH�}dߐ���+?����p��"_pޙ����:��hI��C���d�f�t�9*u�Cu���Ul����+�S�)��ilV�:��pD[e�b��<�T�1���ĺ�q$�-���3=�FFg�j�B�H��mɡ���.~��4ߴ�X #W%\�o�����?B�~	N�������Ok,�2v�KVƭ����%���G%")�k�1M��0�Je�G�u���B'df`������0^}�����fI��Q�qS���`�K�}h��⧗T���
l�ý�? �����
��=�=���ch\��ۃ켞��c�9�D�D��H���C�R�/�:� Fy���<��	���鬝=�ى|�{���{P���
�M��'��.ḕ$		8>�p��'�d�f��C��]ѳ�X�S@f��4�㪷J��A�<*8Bxe�� 	�6�V@/eI�?g��FaZG�:�_lg�LV�"���S�n`��e/ʌb�[�����Ͻ#�P�OS320*Dy�:�#7/��{f�����b�U��j"�~��|bN�\l"�@��A�✊�l��y�C�Gv�M[��p�96;��,�8߲ƾn�7m�˖��!kl_V�-Z��Eg�m�Aő�:ocl����u�����o�����1����NJ�t^i�!#2nǀU��J�o���0�[�e��
�	�����ݤ�$ILV��A�w<u�?�`��(���Q�\A8У���c��l��C�Rr��n7�Ģ���ef�� �F�{�� ���|�n���M��:��2�"i�w��+vgJ�b ?��d18��<��z�b"��_��-�6G�ٰ��Uj�k���w��#-����ė�E/���hj������������{xb��݋\X�k5 �Za��!���Q�uTI۲��h��(��
��O�j�z�G"z:7��͜��, ��1�1@]ۨ�,���露�l؇�B��˜D���+rxmc���p���*�A��UnÅ��9����m�=�Zdn3�󲈎��c��N�[��C����s! N5���NطO.k���]��Lu=ּ���]I�Z&}O�~zqS�r
��}���a^�Ҿ)[�C�.c���WjJ��bf��]�4��B��Ե7I��n���9��j��<N! �-�a��1 ��F�0���>,}����H�K��[� ��8�<v��j\ZK8�I�w..�U3��l��p5X����Z��)tE�����W@�]s$z�������kR|����2�{͝Wʒ�Z��Ɩ�L}�n(��)��'*�E㪶F�(ؠ/.�j��C��a]�����[x����/���Nԑƚ[�s��,;	L��績д��zތƁ�������B�#s�y�1M�@?�_���%�茎XW�C:F�X?!�	:��K4�X> 5�B|Uw  �S��kU��G���HX*|�@p�[�Qq�>u�]%��BV���z'��}��ɤ��\&��U\\`�V
9�E5� C�[�(���b?�ƋQ��:U�l$�y�򳥗�\A��ȤBs������g@#G�8�N�u��%W0�?VL86[ɱcɱS ~�������O���68�ï�X�0CW3S'�*�C"*��~bB	��u6����V3���~��婬�T�d���`Ir��s!6���l����ڄ�P���ٞ�8ıZ0�c��GҎ���n=�Kx� �����zZ�;=�{J����3'���ob�1����TeIs�!LE�[�X��q^������q���Q��l�m��ٸ����Y����/\)�x�T���8(�~/6�-g!,���ٌ��"F��r0>��|��a�#l�p�B�/!�R��]u^���F�q���Y=��J^�A�;���ޏ<�ы杘��� Wn	��K�y��i�'���=�~K�ӽ�۲��e9�.�!"RC�L$;[ّ�ײ/O�G����!I�튔���NǛ�ҽr1Bg����:T(*;��|;n �  n
�7��{�f���>�d�p���G������߭7�#�z�����:|о(���c�K"#V$Ka�����h���wM��t�
n����qTp��ɥi�_���+�Q0:7��#�+8ArVq9縈J���h����CKf�� ��"R���/�C.�l���N�FW/8 S����D+�Ɛ���Fȩ#�p���Q,���ni�!܉�@2g���������>�lLzH*_A����T>����m^�֋�ċ��K ����
ջ��d{_�_�8��:���N S���JѶ��d���>Qr�����0�?t������U=Z�B%�1<Pri;.�yG^����iW �?�-lJ��Ct�9��������'��p��{"����_�h	:�$�.ud	R�_4���۞��+��JA��T�ž�j��d���_�!�D��5��jE�G�¶�T۽�k�xi��v&�b�g���T���=���	���d�0ƌle��Τ��z$�5�g��n覻�e�=,�]\)޹^98ɻ�50�]�8���&�����Ş��׼�5��b�%�Ԗi�5�fB��.V�/��`l��e,����xh<�K�T�c��{�wg��h��'$E�:6�$���5�2dIc�{��|hoom˝� �A��V��@��P/���O�����^\�C:���j�!fY'��"�=x���LGn&�G ��:ɗ�?�����NS�[ P|t�ɔ���ծ	NV�u�ȹtP�@��ʟ�b��n�MY �T8�)%/�q��� ĚB�������	�N�_����cP�`��cM�s>�.��������O-_;�����9�y���e�هӉ�C7ʸ>8Xj{��(?����t���|u�Z�"��:1��_$�`
���<�z\�A /�)Pn�73#�T<�x��tw��6��F�n�LL_Z�¨��m��щ�݈����b�4��  �	;�Xؖw�LԵ�N!�9}�� /�-|��N�t<?���xE_��Z�Թ-Rg���hF�l$�Yzҟ������l�?��[�$�Y�3N��,�M���8Ztꁰ�3���;�r��"t)�q�
9P���9g���aٽG�2JB���a�ڛU�B̫��FXݍђ�X���h3h;�w�n$��BA�@���s^ RK�; z��8q�"�����q�V/sێ���(��,���<�F��ub��xQU+d@��Y0�ë="�k������a���κD�l���xe�y^�1+�2M`�v��z殅FJiO��6��]�p釃us�0���u�E�`���S2*J)���
���V3_=�Mq^8*R_�*җG�RH7�/�h�c�)���{5�2��!{����F�z�������������>���̫�{q(SŜ�0��0)����"P,���7����Ν��_r錼=j�#-��B�r��|1c[�꾳nɫ�R#פ���?K�8.�=M��*|մ�|'�����/4�'�O4FT��
�u�X��݆�b*��0
�A�9�q�QX�����J����v��0��ޚ��bf]����VǤ�q1��
��v�&�gJ�sI�$�e��Z\�0cy�̑2sQ|�jݖ�Q^$�1��-�O�A��Aq>
�G��03��V���k]Mz�e��Nj�����������r(B_��0n�b� %�ʵ_�5�����=	ǔ�<���ŭ�e��7�ת�x2�  xUj(�rU�F���n����U�o����U�Ť��@$��ys�JQ���T���2�)e�ԶG#�%]Oɾ��l^�BTZ�ko*�|sd����c�ƌ������^�k�V�����*2��V��.4I�('D��&և|+�'�Tv�Mh)�;%;?���0D�+8.*�} ��҉GG��1f�rSe��.W1<�~)�	�������L�|&��;z�1�.������1p�ɐ�������4qbH��q�r�x�}C�r��D�N�	ql�~��h�������Μ�
��a��m�z�!:��	02P;/�}��5�Qp�*ڻ��[%�[�K���9��kZrk֨��P��F���0$3�JV�S�Z��g������KǖkD[�<��Q%�5"�$p��j�{[�������I�m-~��\I*�LG�ۙG��Aw�Ϭ� b�8��[��|�A{�M8*Պ7��i�
��������)�k�?�Ґ{9K�׷5��%�`��$��1�8�aE���q�&7)�.`�"?��`&����	Gs�κ-bV�	p���p��Pz3����A�q�N|<ҍr�R���\Aݙ����b̡��C��sxG���EeE�z^��*�����u���sj���V�MP~�#^�l�� os��1�s��R�D���V�,�,8�'YK�'�owڼ��%��L��k^�W�З��uS4�y�t�U�[@Ϣ����S	�M�{Rú;���Q�w�v+ʯaV�Y~/?f�i��u�C8�x�F���=>Xm�q�Y�t����B"�͚����(k5����:|j9��; ��O�)�-6y�R�����ԙ��s�L{+/&ߚ��m�q45#�J���i1�v4���I��I���s�CKWi�J������%-��&r����`2%��� N�n�7Y�{�r���zmե6?~_�4�����j���/Z�^k�hD"�au���6���8 ]���h�2^[�!p���.��f�	�����S����8�ӵT���aAK����n`���	���'��Q���՟r�C�";��Fh%z�����#)���k���s���w�e�9XB����M�S�ޫ�ȧ:�b���:s�]�:wLEX�ځ�\{(4o����8O������׊�M��u]�q4��p���')�	'*o�8,��8���@n��?���#�5����Z-h�i� �y;[$p�נ�F��T��`�7������Jm�������E���1m��A��-�O�L��K����u����iNռ!�z��s��(\���L�d����`�yxpz��r���0?<��U)"���:�_�bow�h�ĕyخ}Lк����M���:��uh��ό|�e1Jb
���Y.�7/\�m���q�x;�?��`n?� v�;3t:���r�P���u\ēb�V�������ex��2:'�����-sg��8f{T,���_���E1*8�y�:s�Iή��+�#�����uS�'����L~��YQ� Ʊ�7͎Ƌ��3��c��j�|�~dQ�@:�,�|�����Q��b1�¤8�������?�����Nj$���@��u�wt��!x�%<��9/��W�Hbk�V�EG8���%����g*U�h�q^�7\w��9��U{BS���4�K+�Z���Ӓ����j�c}Hj~n������0K�o�~�S�^�~���إ�*�X�����tX%�w�,�����';U;�m�*���]׈ �3��G�׌Z��rp�������Z5�6yu$�������-ҁ*w,6��=
~�#��9'���B�����hƢ���H.���I��6��7�SV;�oQ]����$zYx�s$.+dA3h#����ڐ|�~'�TI]zZlS�Z^1� 7�2�Ͼ�E�ŋ��9Lz!ߖ&��^�L�JϾvj�i#��|���8�|�ل0�k�c��7���cN��'i��uy� q�XjIP.�-�Wx�ןb�@�m�S0��Y��423W��m�!W�n(\R�{�פs�����U����!�e}L�B���E_i�_�h�o�����XS���z{0鈙HU�y����@��ks������:�04��W��m��F����P[0z���B�5� GҮm5�w�څ����'�?�ߌ���7�*���C��}i�i����x6Ⱒ�
x�-�����nr�|��81���6ν�WÅ5�ҷS��F�
�ǭ�{�wP�윪f���T���=Y��ę��L7��+�����3!����R�$V����a<<�:n�:�eU��i��r��~4� �ԑF�XG|u���������ӏ;��2�H��"IF���ے��?�uw�K ���]�DY�?�Bb�̉j�;㘃r���v}�h@�s�ۘ�������Y/c	馝���}p��єC��!���Ʌ᭬g��ŏMQ�ԩ����hU�.(����m`d㒩gG�k�B�B�A?��A�po-9Ks��# �z���=#���x�L�����D�G�m������4+8�o[_Ѽd%YL�	������r�P���/󖚜�|�
�f�:��w�֡��4����aX�Q.�a��w\�zCzy����ԁS�B.����V�%��������x��%�W���>�Eb�T4���=;�O�f�wQ��[^�̈"�
��lqhJ%`Y�y�ĠQ�%��/{�A-	dn� �+��(��<D螪TV�.]�.��r(Z7;
ՠ[��J��4N���(i⥰�� ���[[N�<�5"-o)8PhU=����E�R�V�Q3cx0����W���֠���b�¾�xw;����R���� ^^�u6X)�5瘄�V��l�������L<Q%<��\cL�U(P[�g��ER�3�����-�7�#�S	W86i����V��61�_�y���"R��Հ�x$�36|��ɣi���FސG6�e}���ɇ�m���t��Z�DCn����	���!UB�A#���s��l��^,)�y��?L�1�~���j4��D�l�X6˛�Ď��2�с���ꤜ������{)��%�Ú�/X{[�>ưya#��5VzD�P1g_��T�CiP��Ԣ�����E�z@�@�d;?��)U�0��Y�J�X bK]]��툁���t���f��2�@��I���g��t��p�D�
�QA4n��L�]q��F���K���Ӛ{��}O���^��SU{A�W�ܸP�l�8y���G\��;aquo��Q��%P���nU��)?�ӥ��H_�S�Щ�Z�BH���
'�i�3����1s�;b>�P����١�xnbO8f�!��}d��&��n�:���b;1S������	+�/��cJ׼��>iE��=r�f��(��;CgH���K�c� |�����"�%h�4�t_'����q�!Շ�����(c�N���󆅠A#Ń姢��bW�B��N*�8\)E$D¼[O���bޮ�	N>��je�@y�5!��r��f4�. [��p|��Z�������*��w���|z?���!���<1��uDG'�y�`W�|	�횶������t�ԗ@�Eͥ-��=��M�~b6|�X2�4?ےw"��}�g?�@�*_V��˒��C>��9 	����T�<���������<J�:��`I`�C�Zx^$�E��L��Q�]v\�(^3��>��R��v��(�yE�Z�ZQ�V�h!�|�\x�G<�?D6K�wE9�]�A�]Y������J�;�ȠH���v����E͛��:�MC�V�m�9Ip��)���GX��HMXY����s�Ѓ���������V�Ͳ��E�g�!�kߝ��P~j�fI�a���%�Q���7�a�7:4p����/'�١���D9q�B��� 9�,k��9qr�f�e E�1����#r�LI)������&�mȸl[T+�G:��Ƹ"!�n�/��Ф����קG�w�?�*���<��F��!b��T�����A�1�=��_��0j!k��Y�<m�WݩN�Z-�Qe#���U*�(�~gA����#�q琻�J`a�z��VA��<f��%�,��I�d����j�v�f3��Ė�1NnӍ��jsR��B��O��r:FB��l>u��������x���"O!4�ǚ!�;����[[6\d
���[{���,V$���³��f�|��6�2<��?�������~�6n�5�	{7I¯d�\�d�Dr4�,����(����вT~:�.�_��`���O�H)Ī��'�?��M��T��p��E�佂!<��8Rh�qK\���X�df�����P�y�c�F�� u��a��#G�b)� �8���ݙF�(��f�R8~AB���m�[wĪɗXtN+�^��y��C�>����A[�cW�r���}�K��5�ӹOĩY�| �]	�O�} #V��֊���ur|ӱ���͚&�c���4ʾPS���@�S@H��.<@�i��a�d�@%���O�m�g����Z�+�l�g�&����3GBt,���xB�EA��Ѳ�n6�hIɄh�	7����+�+5��3��)0k5�iCK&�<���#�,ɹ&1�iY^�#���y����o2���J̊	J�ph.��@���n�VI�p�6_��?Rħ���_��(.|9	�<�5	i���RVy=C�Sh�u���,ɐ)�_����V��|�*f0?�XQ#1�4r�e˘SA�e��Nb�^��U2q��l��?֟S�?#ET�����C����&	�9O��2��?�E1�Y���rC�;
72 J1C�~��W�a��Fy�|����������_��ut��H/M��'绺4Y��E�c��D�WaYN�l��-w6�r���ddzsY}z�?��D�1�+�L��
4��#D�o��J��d5�|m��Y�q�	�Q�*��w���[/��/��?,w� �Ĵ���AuC�s�Yd�h�$(�4�)_�̇��jn}�;^�����0;�5�(l��R֠��XV<�/������������������	i�L���&���}�+�ťǇD+؂(�K��6=�!��l[�2�1%�\1�!��(?�ʘ�#u�`�'�^w��_u�M�ac�O< *���Q���g����"���l˜P7�l���d��7$�S],O�SW��]�t��f�h�&�k�ɔ���F��a�v�����T�������8Gy�Z�M�䕻�h|�^� FA��=�R��v�5��6�(��3$b���-01�x`=�l
�Eh!b4꩘���J�քO %����(���z�Ca��G��&��>�#�Gd)'ϙِ�(����0Y�M7ܠ �&�EeP�i�wbX�]�{uq)NP���?� �>�KN�_��_r%����T�m��
��&1p�2���$A3���+#`�vWfIA�:iG�Q��u���v���z�1��+��K9GH�槕R�q\�!�Z�㭛Mٳ���a��ƕ>�>�%
"�[��;����a�IQD�w�ie��~�W��+o��lTܼٲ��je���X�v��P񧆑tI�����2D�R�L�]�F�3t=%6��������	޼M�^3��������0��[�d:��*�Wkj�8����+�Y�r��@>�=<��+� �_sёKCZ�~��K�hRy��/	�m.M7�'k�qQ�G�;*z�<]��YFSm����-�I)�����W�H��@�r���fOW��9e�fN�">�"Q\3�P >ںD���)�d�K� Oߌ(.'p/)�q�=+t!<���x`lor�z�f�T�"xUU]�|�"I�B�-(P^گ1�� B�����T�����w��A��	�)�Y`��q̲N�V R�uRڝk�Kt���I��bX�����}H�s���z��F"��:������K6s�k�^�?����גԶ�.Më03�
��B�'_M��N,�ujYM0ɱ<j�'B�SN��0�(z4��=yt��Gؤ�#��aG�󞳗>έx+.��ȯ ��@�\l�{���:g��{�U,iOw'��W���/' -�Si�2�����}��ڼYA�|,߁(�c�
������-����d`:��!�����7<#�yG�o��>đ��/�N������gƚ�pr��<�:��<l��j�	xz=Z���������z. ��i�=�MA����U�\����<�G"��Qp;��fi?29��}���C�S1�!�)&�~�X��}��ieJ������^5���}�Z3 N�����x���Ʉ�����A�b9�?Ɓ�_�-t�q�q�?��с��/4�?�X���GV*}�Z��`�I��)6%���	eN�y�Nv=�L�����&5ۑ4�jA��o�ɶ��<(?�g��#��A�}��U���`&a�K<a��G��D�1� $6K�|�<_`�_��,�;���]�ҕ|C�Q:XZ�V�u����&�í[�鍕ݽ I~b�Sn����h�>�#�����&��R�Ŏ����}×c�Q9.�ZU�2@�����p*��`jeja���u�hl�(��l��:I��@�.4�&��f�dP}W6����)���\�&r����Hs�U �oLfI�d��T�ʥ	��*�c���5��w������s(^!p�g���h��H^q�]( ���q7��1+��O}�n9��X�Wp�'O�6��01v4{����s�.���H,"d�R;�n�����`�1Ћ���җ$%�=In�l{��I�3����%1�`ԛړ��πe���_v�{��z��Pq�.~!���&����ǐ�y|�pU�Ԙm��p�I���Y~z�9Q�t�H�ёe[�!�T%�	���DYo��ր�'Ȱ��Z��c�Ⱦ޶�TtP��R����Z�����x0�;�E�:@���8�Q{�MX��]�HK�8�ur�p@;gı{ b�F�B��<��5Y~|���z��_�n��=W�Ƥ�o�2��z�?�W)�w���25R-�l!.�_�CGNVh��	�F/o�7$N��l��هZ�J��Lr�Y�/N�����p���?x�}4�syu7������1?�Ÿɢ֏mp�~~�>0��D�����o���������B�-udT������*C���.VAd��/ၩ[ȓ1�b��������Մ�|^��h�$�A�dqM{��JIE#�:�%���F��^doB�<J�msG���K���*&;�M2�`���&�ay�r��^��B��$Fa2v��Gu[���"����gY!�x���'M	�z�B���F&�>�q-��PI93n��Q�A"��V�z�E�eN[�n�����! 5�~3���'�� �
�ě~ǃƖ�\���e 	%c��/7�����}�Xx���j����s���9N�hb�]��:�<r#'�H��zJ�1%�b�t�!E�SwQF@er(c���oɦl���%��X��~�gtp���uw���!K�F�l��wgk�E�^�́d��D��1T�C/`V�x��8�(0�u���x��W����Ej\C�z���BXwe�����S|2>rc����Ҏ����{���ĸ�c�͵�;�u�L�G�a)�,��ga	E���F�rv�x�0M�������HR��e�0�>)5�F���{�[(�a�^W,% ڃ��YR��wU>��ی\��Q:��г5���@���Իwv��V8�}�{g�|�&�6��|�+�[ �G�ww�(K��~4����ˌRV��3i���#w��E�L��<��-u�����]�ԃ >��<�(��x��騔��0�ځ	:�����i��ю y�`tf�Ұ�n��(�	r8�(S�q�M���	�$bX��x/	����q�UЧ*��[� ,`��c0bP1����F�9��TY}��ڿ_D&R:�"���$��-��V`�����CV�Z&�qܾm/�c��Wq�B(��V������j��$��2�{��	šSТL;!H	
�#�X1N]Ώ�������w�O�h�����zpNqm��ڐ���υQK�N�QY���^P�^��x��dǒt����^�Uv9g��<��C��߷pƙ�ybc�e�ؽ����r>'�[��B��h��/���¼j����L�=�VfN��ެr��(��w�d� ߖ���N������P+���|�<��.=丏���1K�;=����	�����Z4xZ��)C���w=r�6�SX�"�1*�[
��v�����v
<��Hg�s��|(f.mv��4z�0�����K<�M䷪�.��`ǝ	g e,���P!�;��g�h��hnX���[{�k�l.S�4�,��f�rȟoG�Y�"�&Yb��T�{�����N���t{�R7�p�|*̀.��g�r�'#Bivű��DiS�C|Ґgq=+�ﰩ{9S�x���1���U���C���E�K��Y�:��B�d7��΂��Y/kwݓ�@h�o��P�1� Z/���p�*~�Y%,��[�"�!�l�in>g���k�SQ�?���ʭǌ�9�[���i�����;{�ª>'_�F�D2��P�覆0�%�sO5d,ɷ�s�٢�bS�V�K@�|	R�^xP+�u��H�A� d�,�� (��;ԓP�����uP�ww�k|Pv��`U$˳>/���N�]�Y�+�P`���%���>�06�iC�S�񶺹}���Nq������3��N)��h*����_\��M{�F�:3E�&�����1��q ��Kݨ���.(Uq(��N�=X�����#��� Z��9�K(��ئ��5�zJ�d�9M��L�"���}js,��=i8gά����+��i&�.��g�_*x�,�|�N���9��h�X�
�	��"s�ؚx@�BR9ӥ�%�;*}>]ن
F�r����|��;�~��g�ۢ������k��ih�ր�O�>0f�ʑ҅D��hǄ9��Z f_��@G�Ȥ��d��L[C�pH��{ٳ���v/�}ŹPwB��^���FI�oF^��d]f���
��v����&܆�)5��P`"?��bP|t���-e�Ɛc� ��^NjE�H��m�"gk3�;}#;�i���N�g�}�f�8GܷJU���,���q�?��:�HҮJ��̥zD��=��F�`�^��C�=T���]�<A��p�X�5�MgR�Ӥ���y8G3�6Z����D�ȷ�gη�@�iG��ly4�\�.�>k\Ћ��]*���V�D�Z����R�m#\�Tn�}�^-c�$�bَi`�h䇭S\墉;5 "������+�x[>�
�C!�®�x��(H��B�фз/�G��9�5��e-�߶v��wR%a�5�yUY�:�Jqm=Y���`��Ǆws�e�+�~�(\�Py�Z���k1�����i����p��R�K���v���[��r�l�^<��V �������8Z������M�����Q��䬲ʹy�R�X0��eet��G���9��&L��Y��w�zn���F��ZRmKІD�B�6��|�6	[7�V���M/��F}G�N0����ɶk�׷b�T�S�j��X;D�ι>��������֪�g�q���iL;���Uo�B�b�P�7�>cɆN�v�-9�=-�S!�$�o���*�.������Mw��\���n���@_x��%{H;�)K�ZU�,��o�U� p[S��iE�"R<�j�c}�����6F��&�K�́/H6_m�C�=&��Q��T}��bi־j��E�Rb��T���x�d�u�[fk�o�.�Á)T����Gy�� ~w_�`�07����j��
���]I4�*�ڏ�@��5��`����"C��K�4t9Iݪ�(ڇ�����v���-�j�����vf��1s@tk���Pv�J�<(%��4G�����J�i`l������w������QX?<�5:��Z��e�
y��pz�Ġ|)m����Hҩ�.&��������ṴѠԪ�]��J��tU�8�_�U��k̈́���������I����gRYɒ�r��(ph�5{��2x�e5H�Ϯ:= {ɣ/A�+�;������n<Ɛ$XU����o˚�S�-�;v�Y�U.p���{0���&v�v�d�^�O��w�t�gܨ`��@A���d��9tߦ��S͜ĝ�!��u]�f=e�#���	�9
�&R�B0u�������p���r���oH�6O*|�x���ԗ��[cr����:Z�Ͱ�7�c*�m��<Cݣδ"�H՚:��9��jƺ��+�9x��N�!�؉B�K��d0�x����F����w����`1 ��}u�ab� ��3|�L�#��_-�ˍ��](�
�|G�PfN�M��Q�T8\�9�m�f�M44����>���*o������̒�����&�4�4^U4��@y�}�/m��r���YS����F^�N:��7ݍ�[���<oP.
�o~)T2�D_1^�ds�f�²�$��o�b�&f�jiJ:��S1��)��he�"�;��5��V��9��m�![����E��g����N0�[�)*g������pJlA"A�mHv-�Դ�Z2������v۱|�?��ڈ8����w8�9�\���l�B��JE8��C�1Uz���9�L"�B@.��wY�2u�����O�~ ,���T��щs2���-@�^aSui)g��	H0�����/���e�Q��ᱴ�O�@�P�r���w >}Fo�i�g7��5�_�42�]�u�����
N�:P
6j`*
���,�P� �#���<)~FU�ͯ�>ڨ�i�N�V��?�8��EF�y��omY���Q7>Z%C���5��C�p��RC�7��(um7��3w�����_
���3����X���/�4/����c�l�dh����@?T�
�^_��&�WH4����ˡ4��[��}7QQ��Ĺ�S��.ϥO9����#Eĉ��'�R喅w\�i�k�B��q���k���v����|K�6�7~�US=�`�'x��1�/)�3+����2��*w�0�fx{�.���� JN/zl�c�����h��]W$Q�o���'�5�&�G�>R�������Z�.O:Pk��}nد/�����0���M^�^�ٯ���°�zz�"?u��knk�m)��~�ׇ4�J`������y�[@��0檵�\��s��(���:g8�[�J�*z��1,6��@���Pݥ�h����B��p.l� oK��2ˏ��G�?u�k�ێ�]�Өl�|t��'`^�`����c��4��E�ҡb��Ef��?r��hŇJ����Dq��:0cc�lV�F�rCl�H嘰^�THX�;-{a���A�t�����v���n{�
��E��ո�S'�a�Z̻��̈́��B]+��k	� 9�?�'%@m☸U=s�c4��z� Qx�*Z1s`�E�l�����8qI8�
4���)G�L�K� �1��]�U����-�Tt���������=i��ש#1��+xsJ%�: �9!��RG����GP&n-9^�(QUэ����k����k�HX�0b��İ@;���[B�-m�~����-x����?��B�owo�2���}��sN��6G��軸sfQ�>�[�:D��]T��$�����+�˞F@�Nǡ!:a�!,F�ϱ���۽ɢƉY��*jM���OvA�T��	�|�f�I���Ddh�@�:�fNKDSϼ��ZA�H��+�k����b�Wؘ9��mfeX-����m[v�­:`2k����^I�\8�E���� M[���f�>^�k��&2a���������%�ۖc�\ �i3JA�(�[^���}xV���j�$��p���@̅��`W�=.�2�E�%��ﮣ2}���&�7���U\��:��Y<x.�7�L���^�~���f+)�uUM���;�R�"�5�L��1����נ9j��1���&V� -�q���yDG����$�~�-��(�,��v��󳏱�<�#��p�ǙE���%&�����v��N��h" I����,G��;�9%հC�s��d)K�"�r�ȀUhx1�B�����=�.�׻a�x���AdUB=# sP�����o��1i�{ԇh�^�5�A;I��Die!>��f%'�_��g�8�+��eOk�^+bb�����L��a{���0$^���
�Q"�@�7��nt��_h�#�������sq��i��Y�f*�����B6yIq kD���Y6�^��c��:�nz�REաz�iL��el��51��Uw\�*�T���q460��ɥ�/K��p���Wk'?�Qm�n�{�'���u�2���b���8�_~�,�L/��W�_�{�����z�A!	�~^O�p�<�K��T�E�~�-�%�o�����f����������Ŧv�b���b0D����D���N�\����0vŐP���=�1:�0��x���⁉���I�'|9{$��9�SA�h�`�HX`0�|��v���˧IԔ>�_��Q�W��Z_����N֓�5r���Ou�Ns��k��q8���N�r�Y�7Z�<ߖ�ښ8S�Q4��
Cl�X��|�� �6������t�0P��Ń��p�Z�a�K;���+%��Y-��}ɶ�W���Û� �`�Љy�7,|��V�-�Ţ��s�#"�d�g1��t�O�1����P=h���O]",��e�\�Sp���.<��̢��R^�dS�ja�c�6��I���!̪�w0��ޥ�)��a�DF�@�P/Y�V�.���\��s�?���������c	k������[�<���U��ʔ8��_J�;7NT�[-CZ6��;�[�~C�$�����ERy���7E��pv}��|$�����I2 )gi/��G�0�ߥU��'x7���P�pAA��>t�Br�!f�v؍^� ��M�A|UL�0�a�����X42�E��k�ڱ~Lo�LBw61ő�/�> |����b��
s�����?����?���!�7��yطi���.W��p��$���'��3X�R�n#����Ye���Ӷ�x�N��T�&����
dĄ��_��r�5F�D�#�e��_FO�q7�Ӎ=&X�Q^��e���!���s4W�Y���]
����}~ �Yc�?cV���j��0�KLg��rGSt���y�C�şB���d]F�r��->.�6\����D�"y���/$�]^9k��y�s��`+F�y0��K3��vZ��b�l����Iax ���c�&��*�A�@W3���jWŴ���������B`Ө�\u�.L^?�Bg7	F��T��e�e�����Jۂ��1�`��Ǥ!��8�4'�þ�c���~@KɽcD4�S���
;�54��BG��m��B��Ag���3�<t�~��i��@p������6ƙt�S�eS4�A�$,Q���<��v����ŧ���"��'� �}%���ʝ�@�W|�����ey5��&�&9Wo�����r%SwY`)�����s����B� �&�O����wY�|��U�H����Op����l�jDJ����H�@Ʃ�FQ��rZ*���B��W�t>�M�`?v�]Q;r�u4>�L5F��0�Mk�Ρ�,)��U����g��/��E��ZC�W}����w��tO-�2�����	�HBFT��Nأ%UCW;�<�l��PW§a{��_�h�k��a�B��+�C������\�p3�����Ĝ��両����\8���Ih�oД��N����� 0Pq��i��RvHsLÂ��ɵ�!��h{D�W�(���o�t3�2���b���?7��A��!�Q�U�SK]׃��L�/:��'��]�8T��_
�ڨ��	���n�'��sa�P��1�e���4i�����U��<7;��l��"���ѭsss�2L🖛��y 7��e�J�����R�jU��A@>���T�/�t��f3,K�ʈ=ǯ�<`쮵����Ɨ��}m���^si(as)�Zn�X�_�+�t��V��ߺ�$E���Չ�V(���,!/W)Ǽ����$e��"Y~��Jeg0��<�
��|*n�a�\M�1'���W:@�k	8rot[�3��ij'�ٮ@�#G"�K���d�"N6r�*����#�n�ebo��
c����qL��-uB��L���H���#!�!��픲w��c*"�����u�U�ܼ}'�ж�V�,�̓$�=Vz��Btf�v�a��W�B��{��O�N&9
��P��k�%Ϗ���vv8�gY��r�h�(Sz�M4oIQ|^(y����"(������_ŉ�\m�\�N�xd]qw�����"�Ӷ)�� ���3{��kΏ�����x��9���mJ�h9kK`cWmOx��l���!VK�[��a`�XW�p|^�_H�b�$�������c_)(pm�E^vj�[q��-(r�<�H�ڕ*�:���G<LAH�6|x��^K҈
�~�ܝ#9Ő%�_�e�a�N0	BX]���U�M��=W	=�e&}��<���A��U���7�ϰ�i6<���15lmy�";�MknV����O���0p�ҬתIN��^k����K�IV[����B!9�Z��S��HN�/Mq�K���c���
 �h@��V�����qW�v8��o��Ξ�7��
k���z��c�z����7�(i]C��$YdB����/�����:���n�ތ�q�����83�l��	˃�-�4�VcTi�Z�=c����?84�k�pP%�a �Y����ID�������������i�LS��o�����/�����e��E��w�hH��5g�޴uЋO�U�������'��ypkb+-�M��S���
�E15�W	R���y��g����	8��,x�L�m��D�� m<*��=VH�v����07�rY��$�"�M$�]@�k-��Q^*+Q��Zw��djٗ�3Rt����sY�B$���G
vSZ�=q�2i��ZgVJ�?��^^ɶ�J�PL�"5��§��.B��%��@����@�\on����Iu�������n2K��7�Ӿ;�b�}L�q��T6D��\���s\aޯV�AΧ��ó�l����>>�;�jF��^29�W-����&�����YK���\nf��N�i��"ꡆd KF?]0�֯T$��&Ғx�W�OAv^�Fxg����~��2! ]���˺}�C��2�D UjIh �q�V �fϿ�e���)��� ��Rz?�����v���[_8�p�0�߀WA���Y2kL��}��~�Wǫ���p+���r�4y.�^["�__UB_��9�5���r����N� µX5
&�(����a-�$��.�74|J�yrΜ���#���x�}
�S�C��/pp�૶�c/��Q8����'�)Z*��	��C�B̭���������"X� ;oD7�H����/�X�e�x���B!@�:�k�ӻ������<���W��r���	�a���*��6�Q�}T�)�'��o��z0
L����!��L����:����K@wH d���X�F�zP�J���u�JbE-�K�v��
��(ϰLcx�>q��7���w��������n1<p�1`���|��r����`N���v�$����W~��t�-H����aU.�{u����tR���J��S�������"
1����ZrCT����ܫ3Ѯ��4 �����(�Π:*��\�TV7����3-��@#'�H�N�2!��g�e���F�F�(�R+[1����m!gK�:��� ��J�}C�r=��|��XvGZ�8U�f\<$�Y�~�m���
$��-�ڤ���ʆ_�YӀ/�w�TܣC�`�s�K�$0��˽��%A!Q,]�t;���m\�Jv���14��@Z��F�/ eQ����z�gX{��Q6�]�)�7�q�Q
(2f�W�*�biRηB��t����ߏ����ޗ��7��ܶ����2Sk`(a7���`}]l`yq�:G_G3������fz=]r�Yr!⮬>�ʞ��©t(f�w-Q:lm�7	��_���B49��7�J�9�����A֧�[]=�ʞ���%I�ѿ^�wy�"%|gї͵>��$I�Q�&�B�X�#x�,S��7m��8ּ"�l*���8 ���3�����+rH�p���a�Ũ�Vr�7Do*�����%���Bu�Pèq!$*���Z%Ys����Q6c½����4qU��l���%h��bV:�]�0�Dr��{����RX_�!ü�j,����Ȏ���9A� �o?�s+�ő�P�9�[�JѼ�Ytٞ����$�K���W[�[ߕ��Rt'����F�7��N롺�5� [=٭5���&���s���j�LW����7Ʊ�O���|��0��"��J�\�|#Y�0Q?�%�Jqq�mo�#+Lm�&���^v�c�Č�ɬ}��<m���F\�G��e��>��eSēW�R�K�V!D��Z��nE��������,���| 
4����$�1���b�m�.��c1�)ּ�ͦ�����%A�]{h�9�þWz:8�����'u{�m�ֽR:Ptn<fXT2���V?��|fz<�u~h�
�D�d��d�D�DPE���y��[�-��ɹ���v-࿁&�~�m�2����s�4�Ҽ�ͦ�6؈9����>�Lxy�c��ڿ'� Lch-�ج)� ӵ_O�P,`bī�>�d�KS"^�o����Lr4��� �	�cyş@���ŀ����ؗ�����]BFBG�M�m��=�^���р~�sj�B>�����iZ�BQ��K=�y�r���}A�s�>��S(�^�a0�򏪃���[����4��X�!|����,Bݨ*ӹv��Τ�vW���S�(MP˝N'�]�F��e�f�0��I��XiH0�m���IW�'�M����_gS�Ą�_J%D[-��G`/]1y�(�o#@��:��X{ڿ5��pPҞQ��i��<�i��Yî�U1��ҟ+;�)�6��&��K�8�z��#-a<)�d#߫���t�UD"���c����zH�%j���~�����T���)�$�a�uL�[�������㏓�r�s�����z�?N����Y��=�f��e8nCJ�� ɲzt�D�ŗɑ�3��m}-2	�v�TW�(�A��{�v:�9 Ψ����"�b%�[?��3`>���4�,�)�)��-Ân��?F�f��=� d5�)U��Z-�)��4���ἦ��c2����bά�_�Kf��u����T��5@��r[lrz��3L��xN8�Mx؎h3â�S�:=��H�M���䞂�5�_�]M��q:?8a���\�$�h9H������p �T�'�)=&��YV�g��	�g�c���@�r��Ŋ�v�=x�<�������{W�����qbB���Ձ��5�o��]�|P ��q/�l���6�^��EjuofW������ѹ���paG����?ߎ����_�#GNjU{�5ğ���l���M��WQ��0z��'N�۷�����c��$iIk�t�F*I"<�����jLے�e(8ͪ��M1f�Z��2]�BR	(d�=���bX��@CH�}��j%4�B�L@S�=K�3sA[
���З���[&�X|O���{��]�v*+���c&�]Y����!;�3h1g����{�lj�����N�/���������<A��g��K�}��6�"�6QYH���u���I��n�"���eb�-ߗ���3q5<��R�Ζ���mp	�m����k&Z�w^w�8�-���<�p#��2�LEǹ�i�����j�2� +���.D�����H���\B�|+95:��ǆ#�)�k-�|W�p��}�.K��РN�oڭ���/ �@�ND��f����|�"���ʻ�/��u�CUIy��֎��uQֺN�*iÿMf�;.���,F�}�-���7��F޻P3N%R� r"�.�n/�Sr/�0�ɓB�G�}�⦭XGW6�f>|
X�~q��X��ꇊ�Ҫj��X*�����.�!ZIF�6e�M�����z� $��\���������/�&� I��|T��7�o=��� ��U�T<by�+��6��wtզ=&4xE���V�af�ފ�Ux�qn+��������2},�WENɉ����Pb�:�W80~S9-����ܶ���#(v͡g�m��1�iTR`��'蹕�����Z
qn�:����oIC����p?ϊ�U�࿪�:M���=G��'��YI6�h�:��Hv��|��)��o�P�+����;�m��c�̮��qs���˰�9��?��on�;����P9p@o�8i�΅bHl�FHu`
�QOj��_�WTT{�۴;�=�[�\s���^�d�񗗌`Y��&�C� *iC�nF����!@�v@��\�u�����/N�E����?�g���60�����}��u���D�m���ZX��V��q�՟��"̣4�`ͥ@�ߚ�d�<o��i$���N����'+���2 [f�R!���� 7Vr^�-Q�^���ES*D��>+��{���zӖxU������P�4s���P1�q�Ox@Կ�̮p�H��|)P�����c�&H�p��|���6��������x�6q���Ҥ�q��n���yW�����(mW���f��_��&�_��QH�8�m��°��D2���$����%Aw*������ף��UN�斞������)�.�8�C�S�Ľ3G��HH݃��A�B�s�>��֍O<׈?0|+_�݃�����^I8$�{���lA���p͹�}}�����a�0�Nr���AװYdKd�Q�qP�?�^��"1��M��)cQ�dU/P�+�cH^�R�@�i�'ЌX�P³D��Έ��>0ޱsR��DYa\D�t_s�4<607��0��-�g�����5�/�Fh�" �D#�~H�y7����(m
؇ß�N(#_���\goS�2�r����gǈ�CgUw�-Uv"̦�������Ζ�+�
���j�n�ë���TK��i�O���C��C���2v�7u�q�������0��Yq/^��+a��TQ�dT�?F�?s~pJ��t:ԓ8~��A)w s�����$���4���숷;,�?T;#��T@uh���OI�HJj�X���LlX�)�uh���c'#1�:�OF2�1AbY>_Zxltfq]&
�e���gH*ᵛ�T���R��m!%We�r�]0*���.^��Qi�Z�"e��:�Ř1`Y������s���	�D'�vАj:���q?��57|�?2�R\;
��\Qs&��~��{�a��#��J�����>�����	.Z������"��s�{��Z�`����hH�앚�}�/��9��R�������UT�h���3
��pd��U"A`�C6�%���{`�I���K��SJ5�~[UA)�ri�N��#L*��_Bd%��(�Ҵ��r ���c���h��K֣RM2QyAK+�/�O�#�b�/��J5��۟V7��������Y�i���`��l��O�B�$9�Ü��ȸ.\9�a�[��h��-�ϮQ-�?�tJ9Ĩ�).3Oq�O���`���=�qK��Z��gy��Rb��p�ǀxae�ء �`�~j��=����ۻC�n+���/�_5���;�U!��D9PR.��#�hx�Q�UPhn��x
�)W�, �L���& �:�ўI0��K��=�$|�*Hc�;ȿ�����A`�2�����.�ENo���ZW�D�����֗�)��4׹�%��C.�6Fd��ن�[l�(>.{d͡�k�,��Y�$W{�_ɹ!n6��蛟ð�$	t����j�_y1�eK@����C�9HDd-;�m$���l�sN�bǌ"��D"���c�����L���y�}����粽����b?�$��3��sG�W>�����������%���[�?�~*���A%��:$i"�eɊ1v������b�\�?�Bn2��`5�ڭ�4.&6 Qkʲ�x�UEx�eI��	G�s׻�,��6�l� a�+��Qǻr��4%�)����La#Fڠ��w���u��(#�Q���<1gv��48D[pޝ��VH�-A�	����KL�׸�K"�6G�ź����=q�
{-t�ul1)�-J]��h�p�=��kS|V��`��4�St	���k��;!��_���Bm�o��Nw�D5.�DH�g�����7�>�e�$������ɞ��B{�y��
�S���&�_S��s'��m�G�D_t�/t�F�S�1������@�Ӥ�cqB7GH.�9	�Cy��� b��.�]�����F]%*���η򻧑�Fo;�]ۙ���������-�<|�vBj�6e�~��t-^+ݬ�ݷ����39Y�j��_��N]�x҂�L�EVqp�Tj��\-�ښ�J$�5��v1V���|Lqj֕~v]�{�ΰ��JiX��yPr�I:<8����8�TI�|�c�L=��[�X�|.�Bޱ�T�\���M0"������Ɣb�1ʚ��P�?���mz�{��A_Z�S��{�G��`� �k��ֳy><�%�����t�/�(7�.l'��Y���.�+)�+(z�_��NM-�,x��n���w�Qd@�J�����h������:�0Y�{�EN0���@��]��cR	ZV�C�0��g�P�f8l�5���X:�7Yl���_�`k�����~�rb�8N0����1T����(9���|MKZ���ƈ*�'�kW�։��U��%���=a\����L ��~5���~`��xp�ǐ��	������y5t�U�ɵ�ژU��g#�6O��9�] �Gq�K��x<-
Z�B�/���b����C�V�d�ے����:G���w�MKL�X:���u�c3}�ri:&f)�rTQ���=D�.4w���F�6Sc�������d�n�y��>ﳦ$�������ټj �ޣwU�^�o/���'��R�����X�-��_�h�~��o�z�A;�%�՝��"�)��ǯ��3[k<�~��!4F3R����;X��v��Bg[$÷�OF�,G��4E��|�|x�]��L�q�x��E~���Yt��O�KU�qBR�p�ۅ���ͧ'A�I�ŋ%��p�:�1�VM�P>�xi-4��)X����8����{l�6�L�,y�G�_L�ٳ�O�?�] ck���_Y��Rr	��h�� �"W�)���������Du�Z�=�z��l�n����%5����>	��B��H��~�ы*��K���4����/i^�f�)�4�K;nz�V�:� 3_6_�m6y�T�?_��I��ß߬��Z8��;'�����-+��,�o���!�<{�r$%�?R�*a4�໪�Ǒ�@ۚ��tR�%��/#�au��H�V;�����rZX�\p��Y�$���Z.�]r��W�s=�?SIвS��T�3�?���_yD�I]oJ,v�H]H|�ڄ/��앀̼����iym�K�!6��<=�|ʸ��\�� �x-E��!m�;�����Z�GC��5j>��9���iU;s6�a�����e���팝�@�������Ճл�E����+����kJ�����»��A�:�
KZ�Д�*3�@I���II��$���3����קQy����5��*g��G�!����C��3��d3qEft�mE9a�{��3��?�$�p�]�R��~O�n���].���c�6�d"ͷ5����L9Q����)%Q|��x,4�i�����L�A˪Y$!��I#0��/�x�ֆJ��O,#H~�ah?г���	��:�2�[?c�ק}@H�\#6l��0����2�V���fVm��g7���,>Yk�e�?]�I��W?:NЖ�w�7�4�Td�h�z��n�]��?���6��P "�O�}1Anw-�"�ҍ	H���H�����n�xXH2�����i^B�w����Р���xO�`�����xq��
|�Ԟ'~�u���YA�H1�`�pS,����$�Q�� D~���n��K���Xf�1.8�2�e5�X�Q S��A���c�^��ٱk�	4����c��}���(���Pom.���xOL��{5�&��m
�h�����Г�&���!�O�T,��nBt4B�����|��0�{T���'����1��{o�ɮ�67aH��}���x�q]U�W���}Q�RA}f	-Q�vԳ�&j-��g~�oD|p_+�y�����V�b�m��9oml�ljzVP �1�{S�5׮­$Q�6G�Y��o��4�аɑ�.L��v�d`�OF(e[%�:Qu�|r'�A�_k��:���F��^��ٞI�jB�96,�d���&�RP�Dn��A�?�O�#p���@��yW�I�s �s]�oo�@JA!�ĴPOZ�3\�T/"����q��>�\�t��H���b�12Ni/1R��mD�8��˧�w��94�S���:>1�c�"��d���R��m?��3�'Zf,|N$����؏G��f<Z�0���/��	
W�����Lc��d�E��^�e
B��#~k������� ��-��e���ʙ0^������
6ܑ�m�M�#S�tR�������s6l'�·��1_"���笘m�����������SS7�1���\t5���9!��O�2�T���(#*��w��񟱜�-�Q�׌��U[ړ�|^B�7 "x+�uf����Vm�dO>,ܯW;�6�C��������Z�,A�I����wm'�X�2|j��v�d�Ե\yD���p����Pʍ�l�����CO�X-#|?��Tu���O��s��?�#�,�׳�#��F"M�%I����#����@TVÊ�S�@�o�y��u����{cGZ�R�K�37�&�2�!���C_R%��o����Q�w=�ӦN��{�E_�G'G�`��Z^��pt FIz��"�fn Fs�Ab�Z$�� $e����9�,�w��i�����tT_�l��.�y�v���1hZZ���������}� l�}�X3
�3�ɛ����-�1��`�0��upHU��v'���]� :'Z)=�@v�3���E���J�6k>]㡅�K/* ��Jy�^�*N	p8H��$wĘ�����`������e%��V���u♈X�A����eL�hAU��V`���W��(Gk�.��_y�x[X�����05кY��Wց���D�~6uۖ8En�&���J�������b��Ql.�wɘ�&veql�C��[�"��"�I�2�6$��t[��w��m�l�7Gj��\��f黧���k�/��\_�}.v���o3�9vc��Gnb:p��Z����0�2��`��q+	�g-��_A{2�;����׏��Pɟ�����%�C�|���}ݳ��>=_��؞Q�d����y�b�(�&�[F�@�Yb��`ZM�n�3��	G��M+_T���a��}v�V�ݓ&"�'��
R�(+~��S���G��Ф�\���/ڈ��D��KB��A.��J����h��_M��}�3 �G�������{q8Ar˥ӐoD\��;MP	�N��L�%��9��>�i'�ʤ��%���=@~�㿶.�?o>>aip��k!�:��4:�?U�J�ȶ�>�{^0P\�*Pj!4w]����=*��#����.Зs���Ѥ� �Z�/Q��$���Q+x�ʄCľ>ȵ�ny�ϻ�[�nyJk�������aJ�̥��ΈBbF�?禢�ZgJ>��Vr�y�Fj_D1.�	���&:aڧ����.�Q�P�Hm
Q%���2�x-1Qg�4��⣹�cO��)����,�:�h��)`�x>{�RE/���G<�k���gwU�9Tt*Z��m	
����Iˣ��=Y��'�Ov_H� \5*������c�	~ {T���U̵���>��W�3�
룘�C��v]iҬ����E4ؙh�;��E�ɶz�Y�k�c?�N,\���1n�6d�`q�N,��z�����ghT������#o���`������������s��h��+��$V�����Mb�J�}1o��#�q	��f�F�Ė�3���Kĉօ�p�Rb����t:�������J�n��"�p̞0������ �PҎ� 3���8��5|I�E���x ����1]j"=X�S��T�sF�;&�Ѯ��ul�?6��Y��q#� L�-۔T��(�����HG��WT��,�_�-�i$�.kp\@�J��r֗_�@��~|��֥��:���wN1o�kiBz]'s�/�3=j��M��MrL�P�U;Os��2���]����^p|3A�r� 1h��m�"���} ���ވ�ѕ��J��a����ȕp��d�ʿ�����~A�b|�AF
�T6fT\;��neh.�}��&�ښ��NȚ��k ��묌Ø-T��#j����r��PW��ý�_f��x����.?梾oDe�+������s�������:�k�L�O��z��1������'( �d�*�o`���z֓xx���	R���$]�X�@�D DI���=$��PI?�֙���'&�76���d��f��U��>�K��=�p(X�ux�?�u�X�2����8\!�@Ş-�ͣ�/~�7��(ЁS �z>�<�u �g��(զ]f�ع~��=V�R�k��q��t�ב��&y�i�Z�%�q�)�pC�I���E�v(��\P�C)��澦�$%�kB�vb�"D
.�:ү��5�B���)��:�Y��x�4:4B��'$	��F���}do&�Xj���r��ĆT����� f�#1˚K�5��/6�k|�ڔv�~)w}����TN.F�����3Yl�^b�Y���w�tQg�hx8��G����b�tK�@�Ww�#]lE<���;�-�8�O�#����@�2�������F&��t��N�|B@����7{�N:�h�,J���#�Ӛ���y��5R��=��k���u��&��f*E��҆���B+��|�v3�l&�E��!�Ğʅ�d�{K�S�[G3���}	�T��¨£��y2ž?�x���_����x4��MS)f<�9e��0��I��?�kh�gG   �4���d*��)+u��ל�\�8�c��κ�SGa}�K�����Dh�� �J�=��3�7�Y�J h����?�`��LAPJ�U".7��pD��^����Qp�Ҏ��3���E��-��=hd�����*9���x�sD���Gt��ͪ�N�2� *7�#�����Q���C
��|�8`�/�;yk�c�'B��A�}�����ߣ�zGt.��W�����#f���6ܒ넇9�5�H�]��7u?�U����m+�Y@�%.�`���j8h��ȡ������$؉I�	۹���T(gtM�n9w�U6�yx�(Hl���d�)B����lM�^�o�/0��g���P���������r�1L^9Sī��u���T�ϗ̫	dΰ'�C����,sn��i�ԣ4����o�|cU�c��}��ʡX���x���#��.9��?����� g��Jn�Z
�c`W>Wm�(���H��}�� B~�[o�we����|X�_U`d��O߹5I��dN�|��������$6&=�P8�� ï�4ͮK�`͖��7����t�e�Vת�X�.�����]Ӏ����C^>�׋E�'`L)�T�_>�+R��T�m�<�ԯ��40��=� [�*�G #��&,���iކ�����U��^���KiL��6�>0�1�hO��'�ڼ W�����<7��1��Z��I�|����Z>��7�͡��RIo�H���z{�/��h�� 
z2��YLx>J<�z���r�^�_I<��j�\ ��eQn+��E��=�	�5�h.�a�e�
;=��w2��p|�1�3nm�]n)��|�����&z΁Mr�sz5�������'���p:1����&������̺Bd����}\�յ7V�K��ƺ�4���?),��/��\�ߺ��������K������r�Z>�3�s�yd��Wx�ĸ!�d!u/�%J\^Gl ��ӱ^���������U0Eaڈfs>��a-2���o�y���c�w�Skұ���龢fj��L�n��[m
��[#%�ޙ���r�:M���孥��$O�%���`x1=Z��#YN��~�[�wA�}X�d[��i���������#�EyL� Y���=2���+��s�V���gC)Z�*��6�#�,��~�~Q`��v���dڱ�b��;]��z���e	T��k.�P!���n�ja��Pk�>��,��+�A�V�'Q��g��$�d�o]r�v�������p֖��	U.ݦY���^�hڣk�u/$�	+�0�ӎ/�{��M6���g���
Bx��Cm�7i�X��U�?��I���$�E�:ɮ�1�:`#?�G"�:��M�@��3Y�%e�yp"�S���O��^2P��Y2�mr���i���PWv�e[��i�M乚�q�T������D.P�0Uv�'M�Z�s�=�%�ت.�@ �ɀ�E�A4 2�~T�xQr�+�
ܮ�p�m��σ�>��4���|�[@x5���}�՚�.�T�]�+Cr���/ӱ��3�/�4 V�?�Ӆ_��VX�������5n���Z\�B�P���%|��u�L�db���4��q�Η3Ze��h�%���)\�,�ܹ¥tN��NlT��U臅�c���J�d6k���p��dr2�pe����C�4�3N�$�[=�Ԍl��)~������R�3�/����nZz�)����-jZ�4)I�c�|���gs�:�SH���~�p�U�����q��$cm���.�P�@���f�ڧ�^Ò�zb��h��Զ�� i�T�~ӵ��[o�&�V���ìfrI1����O|���L<�2���A\7a>�����&p�
o��!X���o�x�ݭ�A��I�FJ�"��z��l��(fM?����m܌�M�`��%����O
*�PDf������<�#uT �ԛT�޲0�1�	���\'|骍v�xKO���yR�4:�t3���}� �ŝy�	�\Y�4W2�l-��O>�I)ȴ�EI��784�+�Ȁ���ia��K#���,�R,�X����x$����a�`%P�?Xᠥz���@6o���r.��6^��ϯ�s��*�T�c�V�fAx��J�\Xd�YH塏�P���K�C���D���5�q��6pd@����C�n�ҼO�S);���n��^��(��f�.uj��#-A~�&�-ģ�|����bF�
�&m�lz�sG9E�.���Xlj���"�����]A%��[�+��G��KU�UYEڏ�C��G��V�/"��Q���q�~���U2	c&z�ä�KS�%�����9��Ȟ-���Bj w�\���#�[�6sYS���s���:q���f�sqrA�T���L�TUۡ!��5e��������W�7K=Tǒ�����5&4��t��:u�$�:F�D����|+-�m��֋����?�镡Uue�V�;=(č�`ɷ�5BQ�B<Rh��עޣ��ƅ�o}/G�!���y������]e��q��7O��3��8'���f5&�j2�ժ��j�[-���'�Q���RO����Q\��4�y�-��3���Ǧ誮g vw�I<��z�k�ݨ�����7C�\��Ѷ�UQ`�6��`R�������X;�xo�B">����O�&�G&��A�! gg�3~� �d.�N��I�����xY��@DT�cLdi���Q��FX��3j��> Ft�Z=����o*&�Bm7v�!TQ5�+�<�Xc��?c�a����F���dǞg+��5|ߙ��dc3��}�7�U�UPQ�ܿ��%昀�Y �eN!e)��]��y��W �Xe!#��.�<��� G?��^,���� �����:������wg�-	@|�2��|�F���:�� 4M}D?_)�F��b�v��"Q��Y�6k����FVQ�,�Bj5Er�����2n���F�̡�O{�tu�F�o����rdo��xWH���BB��U2�]a���_�a�Ci�V�9�q���՜ۘ0�p���؛��`3忲L�Z;M;�����P�#��t$ђ�� 㗧N8Ļ��S8��87S�3u�Sm�f�Y޴���B;MM�T�>��Q�	���bJ#�?�p�V:\�5r��������Ų�,�Ĥ뀏H����������xN�]�x(�+��[���o(��bq��RjiTᚄ�B�?��̱m*A��0טO���^�e�͜������$���s�@MF|,=�\���������Y����s`�Z����e;�u�'��?RJJ#��
��F��pS/�-�V�?v��_�m�Τ'�UI�����!ڶ��&3d��ێk�9�3�ﵡ@F���H�x�/벞�q$f��սf�������b��C'�k�R"c�o�@���=˛����]��U�r��	fY׌m�J�]:,�Q`�"�{ܫ�M��#��1T�qgw["��H� Рo�HQ��[g6�O��<A�Ҷ������-�g�c������9�������d�o��&8Rע�Z�3�'u7da�� k�H��a�Z��S�(9i����r��[������,������>�k'!תi~J dO����l)�ELhʚ~�Ȝ&uR��{�ȿ(#�D�Z���XA����ߎ�\0F���`�J�y�P�Y�`p���U]<�׳D�{h[�kEu��nqE�Co Q��;�qQ�-���i�|����Y�,}E�"���)zޅDL�w��F�t��[�[j@9�YS�'}i��J[[�_��*�9�U��>�1ÛU�z����I�El	��j�,�6�%g���=a�.�������@B.t�EZ�.>�:�I�!xF��ю���v����Z�ؔ�����1r�EH4[��
��I8CP���xc��>�[���t�RNi�΀N��g�`��'d/�9`�g���]�_�[�?��൤1Tg����،�z��S�����5�b�W�XC���E矝��/�������@|���t}RUأz`�3*y�q9��W3-�}k�	�۪�|�8i��&�G��?��s�Os[xi���Ԅ}�Z(�i�����%���=�7�禹354 ���8�FvqϹ5�T��G� �>��J�^�*;a��ȱ�-��C9L���1�KF�-Oзui]��i!�1Բlu=\B�׫>��A�Q���������3(ﾼ��H�&�$��w1�[�Uf�.��4`� ��G�]�z��0��Ab��ּ�����_j�*ɻQS���YkI^o�A��F�6�ǐ$ń g�{�m�Tq���{s�K�(A-�Ͼ����N��^�ls:��0����_��[��i�נ%z����f�x-���vBx��	��nDX4`�(��"�nwv��%���-�Y����k[�b�'C<�Q�S���K��h|HK���c�1+K���Z���O�D���*6W��ב��7.���!"�~ ܯ#a�Q���i�"���oBv�~o�U���B!͢}��F'U����j	���7�H�`�b��6�ӌrZ���l�u�JvFC`P���I���	F�WX/W�a�K�n�xm:D���l���}ɐ=`�ΐə�y�ȉ^'���u��*��Ӏ�ѩ�
���$� �� �)�
v��-�H���RL�~oS�E��z��ܨb�L�
y��"���()����
�����՝�L�����ڦ���0�V�r �"�+t91��
���`3zi�Al�S����fu�n����x�F��h�EPg,rj.��
�sWܜ>�8�<y�}E�F�q���f�]2H�ݓ�D1DN�Sy$Q���|�d��^��9���	v#�a��T�_����+!��hn���)�i���M5����Xo���3��n}�Ǧ�E0�d�'�p��-�KJz$�nΚ.�a'^@8B{����i�w���ۄjK2�I��y$#�!���_W��g��+���T�o�	Đ^Zr�TN�K후L�r��ɘ���B'�����i[:�&�~�^��;�;�����*YG�"��uL"6�t��m�l9
�o,y0d���A�A�F4�.1,m'.�H���:葁��?�o(׸`��?&�.6�����k��\�=_5��U�p�>xv���y�,X�XG����d{��j�ϰ����$C�ANTZ�q�g19�D�[/��=�ɴ�\���k{f�@�n_��A>�Ї��`�A+�B�����k����W������{�����ʪ��ʣ���٬*(rcd�a�X���U@�0�|�X�7Ìi:{u)\�y;{"2ҘJ:�v���;F`i��%q4S��U����z�h\������<��T9��c�\�����h(L	�t9�bU:�S[ti�?�O} �<eǍ��L�/�߳��!+{�| �*<Hy\���p���X�J����~�N� Y�
<�Z],��(w�B��I�t�S��C[+�4���
�޽���ޣ'��m@����2��A3��7PR����'��%r����X�ɗϫ̏M+�Ć䆉=��l��Y[S���R�4�.�* �?�d^���Ԯo��G��d~�<dh豹�
��~,��j�c�Qeb/��Y��eC�A78���%�V%�l����{�oWЂ��%�~����]�}Aן��9���o��f^�B>�FF��K�;�(�-�(�<��9u�R���N��&����ı�B����gbid?����/u'l r���#2�X��@(�\Y4��G���ȫN�Luߍ��&�y6@�i�K�fH���5r� � �FM�`a�>���+%8(��)���g6Zb�����q���(�ݸ��Yުq�ڥ�+�8����RT��Z�\_G�D�W�'�k�Ke��޽�</�l�:���S��ч��b�HC�P����㻓�2��*�<�C~vM�$��Y�*��<{��tC���y�*���Ŷ��gϤE���v������✯���d�J�r���(�;t��t	A�/�E#x_H�9^����I��Dk�U]�E�-ss��ORq�.���~�T���]%�"yr��<�iZ~:ʈ��\:^���c�x�@��zh<d`�=��z{���d�Z�V�|��@d2�7s8�;@�޲�� >��+��m��Y�E�^���9P��YM�4�����2p�02��ۨ�Qr�^<���F�3�l��"��*��F��t�B��[�9)^�
�k�:��L��W^�T��}T>\������}�-k�%�]�-q/�/��	�X`�����t��V��)�vC��~���>��@��v�/ě������{B��8dV�5){ׁ=gO�H�쟹�^`�c��ǲ7W��dͺ����	e�y��0�o��'��EsĽn�5v���N�	�HpST�`W�����*�?@ffj�Οp%Ɲ@~ۖ�y`�1ș��\�7�Y8I(��>��ۦ���6�b7�D;X�	'Ĺ�l���'��}����m�G��0��a�����nkJ�,�I��N��D�~�."g����sD1~�o��3�m�aK�6���9W��*���|��)�uE�3���_M*�$!�r��^m{ޜ@�dA������4T�i����5_Ŗ	�ﱘx���[a�6��>0*k��w�G�G�b[#�ʹ��,��
"2�Nʜ� 2+��� ��A/�a�,���ȦwTAEE��V<:@�..���e�OM�ʩ9��v����6����
�*EX	ۥ�l�y�G���U"�89[{�rh��Nt��Tt�8����I����cѢ#M5_S ieXm�;vY2�~\�
޳$�>�~;5��H���f��ҫ��"�/�j'����m����������@��p� �NH/2�Y�o�1��I7[���E0���{�ڿ+�ݨ���
A���ȓHݠ.Cx�R�^�3~�Ȥ���a�4�s��o�2�
.� (aw�O�.sm����'������ދ�����a��9�eY$�J^e���	N�KC�xan�/\�Y1&٧���F�9liFR��jG�!�A;���C���#��B�!]�BP���v8}�֟���Ԉ�a#j`�ͻX�
��?�d�#�je#�_23i���D���O���V�o5D	:p�ͦ��Vv�l"�8�^�'��]K$3��w���h�Ё�<�k,z�W|�u�p�8��L�I���1�b���p�7���O�av��.����������ؖ�j����
�PA)�_��V�I���5��;[[�;���w�wy���J��d�������Se�a����f�����3�R�A�ɳ?}M>Y��<����K�����-�>��m4�9tI��\�?"s��������4�S��x�䠖~��e:R����2��i����dݳTJ��F/�ީ�	���TG���j�O�jE�<�kS7Ց'�|����	��:�#hL7�����/��h\���u{Bz$F������vK)���yé�r����x���tU�Ov��(�ma����j���S��ӆ#����%�����L>s�܎��cd\�p�݊���E�����O��(�?@� 2ey:���cB��abԀ�cգc����`Ps�i�Y��b�D�����}s�C�n�ѝ�!*��4�V���$�#�u�s�%�>7Jg�.���R��U��o���VK�]�,כh����
��i
�d�f����掾�C��@�D����x���&8P���A
�U�kH�C#����O:EA�$�w�*;q�$�0�AT@���	A��V�k 4"P0���0XN��\�10k��mN��y�z�R#�a�l�/���E�$.v����)F�^R�*:��Jr�h�2V�jx\"3�gk�v2��n č��S��l`O�[Hd ce�_�/Yw`��^/���O2���%�H��h��&#�b�Φ��2ˮX 7ǈ�Z'xA�$�tDli�}8�#�<�'�ċ������S�&��[��:�"��|��u�(����9vo>G~��>C6��Y2ǿ���H����$ �2g��^�aB2�6_׶�d���)jg��b����؊"oIHD�]2����>�7L���dػ�]>�^ƛ.9�f��
z��Pf������G$2�N�R���s��#�4��s�H�53<�/^2�=`���&5��;i����3j�m���!��v�</
��G�� W�����B%�*���%n�g�xt4?چް�d���@&B�^�o�hЈP�^�6'9�H���u���t���f������\�y��c�˳b���=�`��X�N+6k��a��a��g���v�"���^��E�`�|��:�`��&Z�zt���h���ݎ,[��-�pp!��;a	J����{3���ʫ��T��/ѾְT��h�\����W`�7x��K�t#>���-�h��F�Vf@�A2�z���D`���u�Y��A\��\��I5�����|NW��Y��?J�_8Z���N��*9Q�d2M������MtŔ߆h�v�5x3w�Z��ΔU�-�p����wa��iiL���<O���s���ݟ4��|q��؛A,z��rG4��w���z(�^}�ZW1$���=�H�8F��OMQ�3�>��B�e���P��u��kX� �~�<�[�u�D�����f�U��x�qׇ�05ط��>"A���B,(8m<r���V��1]-!����͇���xo>?���d�X��Q!�Q������^j���Z[(iR�ޡ-H����b�C���5"�/m&��靄w��x#�DF�N��������+��PG����V�O���ْpk����5)3ʇ�K�ؿ�⯓:<S��t��u�֜J��-�����W����U�ӄ�#f�x^" ���e�j����d��M�؂�pm$i��e�4~��Ⱥ^E����"/U�
o�/�7��Vp�j��W��īY�>#�Mb����|`�{��ۍ��i_�v#b3D�J�$@�P�e��sR�mp�����;W
�q���tj�6�B>�dIT�c�҂x7=�9G�p|.��9�[C2K��u1����J��\8�S�wջ3rN�����<��&�Pjl�PR"ic�W57�0K�pxכ����P7�Z�p��Y�:	��$������Y��K�#$<�1��!I�����Q|f?4�uo��C/��:�N�\&�c�������n�dqE��w��3�X; �^����n���DRv]ғF39gw���	z@�(}#�4�+wj�	��I���O��U��0w��40��v�<���Z�[ԣ�\`wg��f��Ac�=w����������IaL���Z�P�j�]í  �b��+f��"����&@����=n�*L�j�<�w�P,���`���!�z�"-�l�HÖ�[���A��T�:/�f�[���o�(;���M�r�i74��j�#џ�L��@����n"����%� /_�Q�*�f(xeJ6�D�z�c;�N\�����������6��0C��ιw D��p�`�[�g�j
疈PG�@6��������q��,�>�H�{m���ت��G�M�^`�C��D�"��O��0P$t:p�t�`�ϭ�În�BTK}q��$aA����r�x'b�
8��֨ r$��Q���?�>E@|t��qT%X�ۙf��(��ԟV�9 �.�1�H%φ�1J��q7�d'*���t1��6�'&�!�;���䣘��Y��N��3X������+ۦh�tC>���tl��Ҙ��O��& u̪&�g<1���B�����} {6X6��-�'\`7��M,Z�O�Im�$�{�r]/N��6]���#������P��wowO N����N�;0���������QEQ�"g�u�uB��O���5�T��-��4�	���S|@'�;
C��G�Y�s����JBp��R0U{��� ����6��d�vv�N�%���A]l�#���<�џ��q����'�!�f�!�S��2�I�˶癈����-�h�l��)�v��@Y
$�L�L2W%�v�#u��	��m^�/�P�V�>G=G倧�ڋ�C���c:��.)��tv���g�����1{\�Q��c<��'>S6?n�Og?�s��Լ+��&yJ	��l�I�𺪝|;'�c�$�9�r�,�	S��c@ꈣ��=+�5�E��큌Y�3���|��
ל�gj�T���U{�-m`c*�\�\&�cQc�!�:,�]��L�U�ƻ�Q�tP��#>9{��!D"�[���IFBe�π7��3�9D&j!>yr&�K��(,�lR��� ���>Hl�b��'��\���]$=,�M�839�:�� fY��>���X��9���BP�\�:>��x.�Z��-��Jǋ�f<\s�<�+ů
���g�Q��cJ�~�'es��T\�פJ�����8u�Ua{=	3g<ƽ��e��N�(򘸃G�����\*�x�_C�'�#�y� �=��Ŀ�[h�y��B�	��#��.q[n~G7!�<�����ihp�W��%����$��W�ח�;8	��D��X�c�R	w6�L�k�5�˰M]�FC��,��7��Mַ�L{�Ш� e�d����v󬒺�(����3q+*��r�Zj�5f2��ȴ[�pC��S>y�`״V������%X+�1�yVf����ģ��������bH���"�,Ir�'y���N詂.�俖��8a��ӛ�D�ڂ(�n�3�T�J�p�-����>��#�nL��ׄ?M���(��U�g,WA}%{�2Y�3q����@:oT$w�� �.Hf�9�Mq�F�#���~���Τq�,ԣ>�$�N"7h���{LS�@G��QÀkF����g�8��	!��Mw*�`}����A����j�?�E�-��>���h�(��ȫZH�����dk=_-�W�%��fCk�?�CRu�W%�����΀F9EF�Aᵀ*��P4O�����ZwC�/ƍ�r�4��}A�r�<�o��r�����W�_;Pq����_�tz����yE�������k�6��h���yd���	_"�F�i��m�
�G�!"����ƨ�3���`�Z��O��������eP�zG���H��M�#�|I��
�]����hg�uǋ`إj��\�9�J�lz"���pwIy�=GJV��$W�����ǣc�č/�A�d�����D�v�x9��ޏ�H�V�6��2����.ඩl�C�)	�kA�������Y��������GI7J6}�FA���Bk�� �$OxE(�<���{�c��]��t�=�d3K�dGW#hǾ&Vˀ,O��ݲ�1��|�gL�S�J/� Qצ<�B64�Gͼ��R��u8�_����]��h�BݖǟI��c��$S#4�|P����:�P�)�]+
�P���J��g�OM/�}�Sߒ%G��j��>�(�/l���z�X!�&�N��qvuG1X�2m��������!�h�x�<�}Q\O�m_�Ɨ=X�E;7b��%��u����mJ��b�u�g��j�@~��rؠ�83���µ���s�g�[�UUX:�_ڦtΧb�0Qif�����Ϩ����s��$��O}�r}d`⇖sn�]#�LfH3|�i˩�A���QD5��rwY�/�:���2�ǐ.������g%j���G���	]��P�%��g�'��r:���(B�>T}ݜ����w�_�R��<�3�ҭ�72��J�����
K��}/�⦩^�_��
8�/�ϑ���~�ۭe��KE�T_�%~(a5[�
j���oxWKљ����c�W��~یF��`�φ���-	f�-L�%�����f�:��tl};r�4�F�ъF�,eP5a�XA!B֗��,�!��7�c���1�UT �Vn�ȩ�EOƕ��S*�`�_)�{����X�#���W��G��^Ǡ�	��
��ο�y���huR��������^v�3�,����mBa�G9��KP'�CY�0B��K�2���v �����&��ݗ���1��]�D�9φ�Lj��:��LF�mu����������ŧ[~A�9�j �%��ؽ����Y����	���]�3�q����%ncjH\��(��/�_?15	I�7yR����n]:�)h�y2�߂m�tO��#��'X�~AQ��i��f�����W���+���P��\�L�n\M��Sb��"�8�΍�����pz�&����Dnw�7�Xd���hʳ������:��7ż��o6�sN�="a�i�W�5���~��>}�	,�ŋ��<P߂88����;N�5"�d�2���\�^�p�]�cY��w>�Z�	��������泅y���/���%9�	���sI��`,�4bbs��d=ľT�c�ߛn4QZ��f�ȑL�����i�ot�̹�m+�kz��B���?4Z��e��4������@���}`~W���(:��I#���4�o�#]ܗ���MvK��A|R 蹄�e�n�R�?�.(��w8N��I9�L�����/��x��%�?>�4B��<Va1�&";V�n����3<3���D|�Ñ�4^7���&�5�a���c���+�C�N s�l��ў��������ߦJ��*y�&��b��oZO��3%����DU@0?�qL�����u��)s�M�"'WJ�rL>D�f�g�c��;&�X�o�i����4�C[N�s'���{Q�����G{!b�PC� �(Z����DF��1<�X��#�|U�1�V�Jdw2����0�ͬ[�M�����T~�ŪDԁ�1��M$r�����a;��8\��Gl��&�>��a�+�y�K�Z���i�J���O��p��=�{p"�\dUT�=�&��tYX�!���z�X�Z���%��n���$R�T�ѫ��y(���r��ˆ#�렾*խT���]�w�kt��)ަ��^h��d�3�|9R2S�Z1;������1G��p����E�2%,�q�.0�ڐβ�uw`�,���1�oj漲�.�\)���C���3���ƾ���Awy_6�^D�-!���	�!Ie�H~��> �B�K�2�!"��}�T�ٿ�&r�R$w/�/���낹�U~�$�����Qc�`��ƑSR��2���uQΚߴ�.{�ŗm�<4��=�}7���,Л'�-$��4''�������r��Ǘ����!�>>�/����)s���]�'��\#,����lw/U�S�-��',�է�&�tH+͜L��Ȁ��u<N���Қ�.�X�|jb�@KS��S�[�BA�oW8T`�P�f��u�ߌ� �����1�8^���ɠ��<c���d�B[$�H�g��s���y=�~1K�&""�H���@�r��VS�~�+��6۷o�:#�]��ɌD8���FV���<:��<!~�ăJ$H���i�%��I�D�Z{!NE�[F#��IF�σ�7�A��dt�Cb�b���f<O<�<�VH��ٻ}�����4�k)��E��E:E�7:k/���_�Es:�n��}b��8c|���~�ؤr3��{�Kc�ƘM��S�ZQ}�O���֞.�繋��H"������ ی�ȇ�{ep��,���1��F�ˈ9��ˇԊS�cw������J͎�$���)L�)h�I��-Y��F������������gi��R�-�P���v/��DgEӓy�mPGZ��?\�P��������}�ȂS��St	8t�Fn�j0#%�k��V"�=��Å��X>���*��:�|:�n~#�TV����I��I�C�7A�{��̊��-[�$z�c�c������y��a�<��XI�4�h�)X&�%�ï�'��c���
����J�cE�4��eN�LC�	��ڃx-���C��Gw��L�-�s9�<�H����r8ʻV1�
�ٮ� �?Щ���R��d� �TwDwҬ���(N�*!T:|�������Eg���޳JkË��ͽ�+k5B=�HFd������ա��0�N�T�����#��)����)o���Ƃu	W|8d=Mc"���DUÊ�e$&U�]qQ��%O��+?+v��H�������`w���=C��p*��}��NV���
DG(M�* <.b"#}��>C[������E^'�^1�Q�$X��ۀ
��'iv�%~<z�o�!Z�����;�U��[By�#��*�PF;��'a���6cS5h/As6���'�o��mus3.���%>g��#��Uמ�/��t�5��g����F�i����G��������g�
ufpݪ��w�/��D����8Y��-UT�\���؄kȰCn���
�e	����c^9h���J7��6q��([��P�-�I"��ڀ>�����{� �(��c"����V��pؽ��4�����t��.I\�F��%�fJ�
�׬�]~��.������U� %�o���M�C��,��z��'��j�Rk�~�a�	����e�T	����1�nZ�R(#�Ř��WZbEm��(H��n�t�<y��=��e�.����ƞ��1�X�=��sV�_�>�i�ؔ���2r�;�1_}&�gc��!�tM@��U*�=.X�&t:��� u���o��J5\�	H�5(��_��=�����
��QY:�oh=�{��˒g&J���ĭ����^��ۡdT�=�ѵ�>�'�������\���%��^J=U�e0�HQ�N�ퟦ�F9H g�D��P��R
穴����眼��t�w�c��.VmCΰ�kK�����e��Z��\$���(�.�6�����1��GN���4+��BԲ�#�Y������y2Z��Ӡ��������[\��7�R�tv��Zß3�y��T�ӡ����a���\r&lw�z�}|�7 �aZ����F��S���X�To7�t�"�7�=} �d`���n��c'0��J<Q�2��'v�T4ׂ�c*�#�=���� ��<���T���s����M9�ayA�l����6\w��������Xe�

mv�^����&�<����ضm�q���9�n��ҬI��	qJ	^���@%�:HHׅ�a��FI�uS&�p��|�Uͯ ���"t�țM�-����^Ll�$�fZ���nP������bڢO�vY���V�:���}�d����hqm�T[ϻ�����d�/��j�����_�Z'��P2z�w\](�~��V��-��'_R ���;�G�����KøA]SWG�:B��5�9Jˡl��Ҋ͓���b�'B�ښ��I7󘼡�z��~E�,I���~����C�n��t�Вo��B��۔����<�aQ�1H�y�%��Hd�Y��."nb�ɑ4o�P5�������)E���g�6��b��(�p���c��i�f�v�rE�lB�%P�U�X)��3�@V0��3��a�
S��~p�uUGP�Fb]���Bjk^J��ׯ$�NJkD��'�Ȕ�p��W�Lt��[@똎oPÂ��p�r����P�c�kϯ�-���GĞ���Ҫ.���yk�>XיP���4��jx��(!S2����p��YlaB�����؇x^�_ƭ���6m2��a�󯹺h*��r;m�6pE@�l���7	nc���&�C���ĕw�0�g-����hˑ�J��ԛ �p\��'_H��;}�5�q�F� �1��IֺU^���;�K�tS��W2�� ���(�C�t�i�5��GP��,�-�z�u��N6<��6W��%~�x1�
�����}x�И�x�
��x�r�M�=.� �t��h����CD5auj
�`Y������e+?R)�}R�f���Wߌ �������05j�g&�<�L�8�W���6ш�� �r���8}ә���k@-/�b��~�B�9�_���3)��緋��w��a�Y�#�.Dٞ��g�-�v��y/Gˠ����:����k��Ni1����_;��Mc��s3����oE-v�8ҊGI�,"�95D�H� C�����4�O����g�x*ԡ	"t|h���� :K5�_�L�3�����yB�'$#�#&8��)*%{%I�7.��u��K��={�NsF9����11�L�˚��O	8�cmu)�.����ʩ7i�n��$���M	��*|=>�Ȕ��g碌��9"(X �������[�tT*]٥�U���̵�6��b�1m�_!�LS�1�.�ՉB��%��Ag/T��ݯ����h[>oܩÏ[P�����;�a��m��K�>f��W������O�u��{��N�.�����:F�wM��||&���'��]�Ex\a��x%6U��ݠ8�\:�q�/#r]�h%�[��)���ܴ3!ݫ��s���d -$��<ao�P���xùd��n2�8�O��Q�]a�����OL5kl�����nz�9��Svn�Z����i��œ��p��#�E��@={?/�:\�7Hsf�"�+��������δ^��_�৥�bfQ�����ܫ�j.�#��M��v��	������.���t�� �;}�=���?7'0����0|�xλ������'�zX��Y��=�ѯRgQQ�'�b4m��j0�7���%M��������8�p%�Y�k�*2VLrǀ�d�RN�6���!h����@��XV�H�#$9�y�q�-���� ͇�G�"�1=;n�Y.ǰ�oF���,˽�+H�u����>�3i����t)������"�6�Z· `�Ҽ$��g��T�s�>�\��0�n���ƥ�?�8�z�k5U��1�4�p�q5��V�,�Ц�	�{J���V��(� MxB����l��*G��.�G��3ܲ��nt��o�Mly��*^} �ʙ��,AT8zē�E<���"���a�vg7���M��cI�Rh'._.�6@��,!'�Cdiëa)J���@�Ӌ�����˅��(<�k��RH�w�\v��[�����=�;Ü�y�b�a|����J��]��u��&�?�y/=E�?�R}@�Y;�}���]`�#�x��"��6�G����pЮѳc�2��p���W8d��$�U<,��ۭ4,a��ߣ�?��ݘ�J[�x�G�+O���k�|�qO!SVސm9$���=v�����o�q!�у�~��\��r�R��]7�c�%�;��7�8�8���(�7{A�v�g\Z����!�l��j�dP�m'C݁&���>��S������OU��{߫�[@�C�-er?�n|^>�W�Y����'gO� �=ոo��C��i��)�ɔ-x�k'A��[��^4�D�������z����ʓ}����#�䞊�eH��'M�c����6=�d��c�$�k4v���l� ��е��,�<wB���AT+,��r��z�
Lad{��Ayx,��i�Y0ۜ� %]B>�Z�f��Ju#oQD�r(zG�;�ތ���.��E��rل��A-�R�o��A�W�i0�f�*�(�W| et��Yb�HCc�I�	��� �4O�~+��G�)s֣�}<�Bw�x�?����" ���^UQQ���)�#K-��=cd4��9���cę�if��m��71�wPf髭�X��ռ D��z3ӛI<���	3�%��]��	�i��/���h
̞?���e�l����h�As�k��\��Ej�<�!DM��l(Dׅ�0�ҥ-�ݟ�F?�7��HO�����/������}8e�9Q����>�Vq�C1)��Vg�td>��R(V�;�ϊ;a�W�ٴ'�T;��ڏu��aE������ݶ��E־��,�;P�B?{��)���G�Z�wy��?Hv������S���T�s�ln�K�"�J2�鹌�|Έ�uCV /�#Qe��r7�_��:h�L�+wڹi}vI���Q(���jRcac^��l^���av/8k~�G1�^}_`1_ZR1�5�����E_��ZWmg�{P�
���l �FJǘv|&˄��\��;��P�MsT����mc�9H~-�b&:�S���nh�(E�8���l�D������%R���_ѝ���#c�b�𶼒�4[Vp�^4�>/lE����gv�׈'�,�v	g�µ;ț�nDE(@d���ݬ�Hxh.�E���S��{"���`��#K�Yaa��*�6�z6�hFs��C�tSbM��s!qӂ�<AmY�@2&F�0s4����Q{̢�ʣ��u]�'���8�ۻ�j�gC�"�{����
�8cf1�o�[�C�_�I�z�	���	��'�6�Q�~�/��zP�Y�������g�`7k�h�]@��ui
��!Ϟ��7Yv�T�M�!Zc�v��8�T��A���2ޟ⌍�q��R���ɫ�u?� ��~�C��~ �uZ�z�M%7n�(��4�D�=��d _�L��^��S�H��\��wH���£��$��Ǟ5z�v�7	,SX?�>��e� �\�\���'P��Z����]�P\�s�����_��l���|h�Ƴ�MWWh
VR��3�Ԑz@���f�K��(���-��1��Lj��i��}F�#�g;����`o���Չ����
�#�)�����g��b�'0:�C��7p¼(k�P쮰D3������퓚sԊ$=���8��1�c9/��p�۟�:2�-yT@|�� �,��W���d�2Y m Ҷ�na @Ϳ���6q�}�j�1���d� �>����ݧ�3��m"\�G�G���u0��S��|=��ӔmB�(�7��lʜ�R��C7� <�.�k4���j���6��ο�dO�797g�
��;�7��Z<'��L%w<8�k�U
A��bI�_c�8���M��\�ް�Jج,9e����r	��MyT݁��`6gςAMŧ����&����ׁ�R�'���u�v���H�W��/ů^钃�t$��"�  ����F����>-*��P)]����~�����"�vPHfƞm4:��Z�_#s`O�m[�X�|� 1v��/�!cQ����`�k k.��6�Z�!=80w�P�%���tc�C���2?�����ק�o�n�=õ���ژ�l(�R,I�G�[=�4:cm4����q� �
\D��	���ɥ7��tv��)hB�4�]�
��ZBS�ٺi��a��Ht�)�������4����EZ#��H&����'|Qq���]���4�>s��R�܌��g�%#�w��6�� �Gt�T	X�bx�&�0�:% �j��a�,�Td�%ࠂ�p#r����C�����ܹ%�.�]��(�����M�_������W�1T��|�����"}Z�<�"����/�ff%�ΖII^�ZzʦB�.X��lE��5f]��,Ŋ�Wncü�n���5��W�u�J����Y��t�O�l{kp�n�|�s�\B:�R�j�����³�v|{�C����Ez�xI�"�zܶ�{����f���m��t�!.��J��?�4c ���lm�Q8UU�w,�hL����Wܲr3��zq$09��"���w���T���!d��X�� N�^������_(0m�\� [e����Kx�;�����B����"��5H��C9a��H�%��l���	"8�W�eم}�]�g^�4)O�~�'���2!�<� -!iG�?D,f@�	_\�A�IXe��z5��|�2�������J��l���S�]�.�kK�4���)ħVM�W��A�D��WӋ�n&t���r#��!��h��@��!��k�흟	>kU�@]�{�Q4{��g��f�+ɣ��5��;.�}������a��&'�EQ�%���X�x�1��*�p����O�m�]���68���\@�Ƣk!�̵J5ċ	���9�1t�ı�:L����L�׮��B��Xtsɥ�O�FKyF��?�J\�N([�j�8�%�����7X�'��vᢁFa�`�=���|ޥ�������N,�r���j�7�귞U�W� B�32A͚�;�����zV���$n�.w�[/�P����ߧ7b�>w:Ԍ��?|e+����l�T,m�Z��_���[+>ڦ5��]%s_�i�zX%[}��	��u3A|����D{��Y�w�� [
�l��!�aJ�-��|����,����0�������_�v+H�W����{�]�O�K��mj���U�7/�n���[0�Q&����ߺF�E~]ט%4SM'�X�u�S�&�s$��k�D��*7��᳕&{[�;�%�ۦ�A��Z%=�U��E�p��Å����_���uzV�\¾ZY��y�I1qs_O0d�46����$�Ln�2U���aWQ�p��;-��h����\�e�, Om�;�ρ���9Pi�����4=(��`s˙X�E�Ɯƪ��qܗ�V�]���Nh�t������R�ZT��]�q�� ��D�nV�C��l�{Gl
�G=�������������x�^���](�P�v�grK:K����˨��������0{�Δ�UB~�o�
G1��]�<�,f���2:�t���B4�Z�t��l_�<	3�(�Ǖ2��SM����l�?�����_�;JK�C	�Zn>TP�iQG�z/�g>aTO6J�`{�/�`�G���gz��jEI�%�
�I��U�-�7�Qf��J��a�K��0=�� ��$�q�ⳳϞ�yS�/�-�o�gw���s�2��pP�F�����~4���/�fR��U�=ݓ£��=�p�Yӈ��e�\��#k&�pWK̃��vIU�';����yi�w�if|	�M���c48Sᢻ�g�gPޗ�f���h��Hc�Թ��rnx2O�b�ƚ�j�6�MT�������~�t6m��Dǽp6v.��D\���y���0z^�X/���?�3LN�B<�Ө�/���U�2��\Y��WW?H�}�.Md"��-�рD�����|Cd3U�~I]z�ǉN�s?��HG�X u��¿r�Yö{d��$ز��ڽ�^�hrW5���F���c�oH�$#��aqϕ%� #[HfrQa�M=Fv�����6�q�<I�����G��ӵ0S�ɝ�l�Efr�A��䖂��rx)��5��m��Kdi�>!�[�k~��'������4	�ųX���|��XTo>5��T�:�l��V�S��ZP�(���%_VN~���R����S�e�<Q�z��g���>s+�#�ֵ�	8lG�UA�J=��� l=�dPV�<�y�P����ջ��u�[��);��GN8*T�J���m��k�L��>���"�ٙ/�5�OH���z�d�b�7��;\��1^���;~Ji��R���V:��F���-JҨW4�H��X�����_>8~Q�ŭq8���I�uX;w��/���8���vF��,���C���M���fo���'!�-jZ������;W�

s�|-�y��[l�����h�n5������=�_1�+���/zvН���^WE�o��8Mm��k=+��ǒ�@7n�wȮb�Ʊ�O��E��a"�W��X�/��~�N�&�j}�e�.Tu�~IX|y�e�S���4̏���:���TCp��#��#�Z��x+�u��$�'	N����~ZdN�%� ����־a&L���i>.q���?݃&U��.���uI��G[���d����U���(�O�㷦�ܾQf!)��c)N���S�+຾ r��\���D�
a��8/�-�[fv{��V������ι�_a����D�H�fj��؈��z����	�j���&���<�m����+�nr;K=ZԖ3f g����")�	l��,��:����$"��z������Nc��2[n0��]�T1ͱ2(�aA3X5K )s$�;��P�Ev#Q E�g��Q�?%יT��*��e�ws�s���V��k����`���\Hy��h
LP��{Ǒ@�a2�R=�xIqU���fvgXL0%+Q�I+�����K��@D=�!1m���#D��.�pz ,$�9��ⷂ��`����Q�/��_���6�0^��6��s>j�b�����R�� ��,��Q%�u�s��=A�B@���j>�!�-��#w�I�s�����Ψym��ݮ��Ͻ�ne�4"�"CQ�w��:��@�!���7p\�[K�LaI�i{��` F��e�����=�3aF��b^����Y�����_��H\�	�y7��� X��S�a�!5��/�\,+ ;�ж��?_�43l�:J��"p�'�.N�*F��u�Ͼ�{�E"]��~���>�L7<e���E�(U�㣷Q�YN4��	YN�?�2O�jàp'� �� dI��� �AK��,���Z�v��8�eԥ~��3 �\Y�jv���&��C���D>HLT���e6��i�����ΡDg��N��y��w�%e�=^C�-q�Y�jC�I�s��5�N��6݅�`�D��k�ݣDZo�Mh9�>��R�%xrJ�ĲU�;��G�2	S�#1��d݉�����2�U6��Y�3��@z{������|$�o��q����91a�z�$6�������V��~D���`?^Q�kWh�}�[Gؿ-u,���V�S��}C�]2&���8k�e�����gA�bZ@�<Y���qkZ���$��$җ�� P5�ܕ��c�[�-l�@s�$qn��$� =���z��Odx?�m�SO��*�0�����$I
��|n���O�ں5t��9�P	v��3w�(_[���#-a�t�I*� �����c0Ei�(}Lg<b3�E��H?'���;ֳ�ⓀK+<E"$�-�ᠧ�|�4�8/-��&���֦�W�i�y�h�M�I-��a�ΖAg��) {�zX䊂S"6aI����<V(����}i�dQ�"��)�N6@+�y)⴨*�E�J���c�C�d"�d!��u0�<6�Qf���.��h [�`�mg�Pm9����.>����m�x|7�JuVuj�D8N`6LJ�v~jO,�m����o� F�io��4�T�9ql�H��X3SL�5�+ޯ��+�'�6�P/Yw���{�~��qLW�D:P���1��S��QG��+�9�Bd��YIO���5�Nt���!e�����#�0�Qjb�;���v�d)`:m#�׎ڜ�M�kC�+������o%�:�0�n/���9n�[� X�����L��P@5��npm͗ԉ�ۤ��ɟ��t��
¦F?/;٢\�x���a�
�#�y�͵��m��@(��
h_&j�p\����P��^D�v_v�ϻ�.��t6��h�_Jչ���D%�I�»iFueH��c8�k�[�0��3C7%��EL�?�{Z�|w�.�0�����:,v��+��˕R�z��Vz��{8���#M�/QY%�:���^�,ׄf��/�1���q]��q샚�����{�z�����з���֫;� ��t�bGM�g��gm������I.�$4�g����rQЄ�Q���Ln��]_{z�t;���`�
q!��iL�;�aacU}RD�\�l�*r����*�X��	A����O�ģ���W��G�7�>Y+�yMZhjd��j��������M��u��鳣'8N�y�U�Υ��/5��;+d� ��ڶm<��~��>aDA��8P���L��wܼ���ξB�Os�Ǝ��Ԩ	��G��8*��=�eq� {�N��k43�����k�h(+��wdACӾ��th,��J%1�dE�t��lc�e��J�������oc�C$��7�V��a�۹�3��D�9.p<���X���ߖ���}V��]���ݒW���8��H��pYX/�Ǽ�����5PE�����,��w	N'����|��x����|4�Ӏ��7Mj��c�q�y?ߡZI�tQ���d��R�Αiy���F�I�<{�+'���x� ��7@�$��:�"@B{}|�Z��҅
%4*t�%����X�祍n>!�
I�D.v*u |AM	���e�Z�f�P��T!F�eD����`�Q��Y�s�78��4�ͽWr�ֆ��W��������\���۠0v��|Xjy7C�s���ܪ�h�[�}��Z$�����"ӛʀLs�+��I�7��Z%�5��-Q:5� Z�\�c��S��Y�HSv�^�x�P����SzL��8@��<��Ic�pY��S�b�	*��,���F����r�`��w݌Ͱ��cC#M��I�b��6�ܽ���$��i���Xf'jMv�qJ�7��x
���P,T=�l]���?�R'-R�H�}ρ�>L)��fE�`�
�r�>]h�@+tTb(_��}��G�9�53��~�{3����[�Qi?��+Or�;��)Y��7�MU]Ao�r��_����:v�79��V^�n�aW�j��ݰ��ۺ�O����2G�����z�*F��k!>���8L-�%��n+9���ٜጬ*ҷ�D��@��~��?|�����hd�@�M�Y�[ \ �����al�'�V '⺘�s��8���&qm�g��|O����CJ9 ��|�|��I��c*��[��Q��3
�z$%��J(��jXUk+J��?��X̖��g��;����$���F]<'�Δ�;W4I1��)�
y�Ѧ�E��xSt��Q֞S�^��8�T�b��w�%����2Dz��HNx!��%��3*���7�{y[T4�������٩��n�6��M=C�r��4X9e/�C��u��F����۵;��(���H��Q��1����@Û�l1������yv�_�ϝ�A:�Z�W ?����PC9h4ZѱR�������C�;�=8�Q�Td�/{P��њY���Fz[�r�Yyd��Z�����/�r�Iٖ�ʰr��4��q�o�������Yg�	C����
�}�F�kD~��3�Ci�H�@�r�N-��>��gR���ۉ?��^&��=���	�X�K-u>���F��1#<�ϟa�Ł��J	Μ�`��mK��
p����B���D��X��7U9���E��?P"�^�]�����K?�dd*A���BP�k����*KA9G�t��S����=*�cH�LJ�WV�o�X�"cg,��o���Z��m6�/�~/1���gR�P�V�U
�}́R���܀��K���x��8��!�'�",s즙��9z�/��x1\��[B�CGUPE�L�����5FqCE���
) �H��-��j�~��3�|� S0mͼR�g�D ^ͭ��h�O"}��jgvhah�T|"��Hg*�6K�^��Xp��؉T2�6��{ G�,%bL��v����3���;?���nMM�B���}=#�VH�vV��˝Ԝ�]�ǿ�b� ��٤݌�q-�(���2�U��ꔒ8�w0�XF٧������Z���~�=J9ks��gx�x�NH˟�}C���S��һvFk���T����S���j�~�|�c�o3k(0���K�t�QuB�lǎ�������i3D��J�a ��BO�(#�d0�bO:H��_�\�!���ic����	�KШF��"�=H0DE7�S��Ó.Z��������)WM�:G�ԅ,ڳ����������7�i���] ��@�H��,�^W��ή��X*�C7����Г��t��V�,�vŘ�C[��vO���_\˧��j`7xn�	�k�nz���ŰdWR2�$�u�!��O�-���G����k}Ş��)��.q��ȸc��HH�/&w�92�5�N�%�6��.��@r��ji]U�vV׮!��qrAdax&����nq�[j��܏Rt��vf�����C��o)��V�z��eG��=�uj�����>��b�fTѰ�IRk%�4���ˏj���A:c�h]�)f��],<Q-&��V,ȆY+ǚ��,�}0z�Ϗ�[�,t�v�ʡ�F(���%k,eY��Ŷew/��/�PQ�f��L��d������W�W[��~W�U�����CTq�X0�R�t����K��q}e�i�팂j���#�l��9��@6�>3�h�3���Ӛ�9�1cќu��v^3OQ�*��C��I\a�ҏ�s�~x�	7�r6̹,��6���s��Dc�ӈq���A���d�:�9�e��HI�Y7jd1U$If3�r�I��� ��0���ޔR[�u= �S���>.�d#�G!�x�G�~�L� �_�G�D��^UҜ�����|��S�Ѩ���1U])�%�OY�T�1�eB!%�CDj��Wg<;����V��~���/]���R�%i�Èo�&���n1H |-L}Y�r����z�`��+�{��p ���Ⳃ��re�x� ب��TeR����J������w�l�T�F���m�ӟv;	>��Zo���g�)�}KR1|`��<�D��aQ�?X�k70���xu����5�H�?v�4�m�I\5���uA�όY����O�w���Q<^AܪvQ ��Dt�w�u�sl�yy�E�7�Bxl��+�ш.K�-�/�|����a�S1@S����R��!�d�
����w���9���b{���Y�Li�]�,!���5�iC1��V����)�L����Ū �����^a?����-�o�w+��#�]� ��x�؝�oZ�Fdq�7�(��-X�)�D�h��Z(���ϕm@��QCԫ	��-Z`���.K�H�q��<�3m�Z��������H ('!.������|�)cH���e���`�>�5��;D�)>H��n��$#���������Q%�.Sh ���K0_76	�v6�]�fD�n�7�X2��Fz��b���a�#	�E����{)����mt>P��YE`4��_0v�H��5�^�ñ��a�v�{Qߣ�Sj��T�u�eX'��T�Q�Ko����C�ūZ/3o8�r���Us��L0�H��=W�1��:�+J��2O�UY�/�o�><���2��3����B2�f��v^�b�Aiʜ�#=V�p�b�z��F$���t�ҟ}�-���;>"72�J���&B�$N��������Y?���ii>��� ��<$~�T�8��e�ˠk7���W9�zF�X%ML����5D�ѯ�sKu���>ռAH�"�K\�#CE!Wj��>��bɌV!b �h��K�b+��h�4ؙ~.б��עn�pφ��i�nQD�(Z��i�"���5��l�B#�]}}&�^�� ��jj���Fg�?��N�h��}�.35Y��Z2%�%��
�Wo7�s*��Ծ��=9CmC�=�p��V^�H R�?�"��d����ݐ�Es`�A�b���IU�<g�UO����ն+Qަ�����P*E \.�ۡ �s�$+ p���~F^�S5�ogq�L����0mk�!��^�dY�<Ҕ�VH��'�x#�z$*񘯬1�T�/�1r�0!��Y� ZB�Of�Pm�����8ŵJ�6F5��� �˽�v{����"�`�ߌ�����i ��Y�O� wnE�f?xش:�0�+\�^�r�V��j�cz�%}"H���CA����E��b����V�P~�O�'�{���;���L� Y������df�ߨs1�%8�?��mԅ�CX1F
%�L�m?�j�����m�J$ź�KA��'Op�!����-Ma�'��v$��m�t�m�\�c�t�<+I���$�AY����Æ\[�z T\��%�s�n
N\�=�V��X0��F��n��fG�����T5&��V��"���F�*�ƥpp��ъ�U��� ����� ߙ�X�O�uqZԏ�k�����x�rx��F�1a��)�x2@ol�8�' O^(�[/S�bT��9����k	��T8�O���Ԓ�c�L�N&xZ�G��P�˘��K����I#�X���E�N$�St�>�^�?>����d�eу��J�ܒ�KWg�C��^�tʹ4F��^����Ɋc�H��^��Q;���7����1S��<�bOd��ψaq��3�s�ʅ4Am;e^�7����αt������>�퀱$�⌘9.+�%Ԏ&�[�5�I[B�@���{T�X_��Y�ڿ�(F���j�DEel��^&�ji�.�>���Cѡ������&]&E2�o��82��׼g�ゝ&���:��ڝ�Oc��}���'C��\Y��%{#|�����{i���{��.8.�0zp9y�Q�x���Hȑ�=t��U[��A��,(���Mv��Y��9~^; &�Kw!��DQlR�@*�i�}/L/󯠧T��ŪZ�jHۍu6�ybI�SM��r�-_���%دOY�R~C�R	�W�m�j؂�Q��8s��$4�� {S�r�`�����H˨)�7��m�X�v"�
#}_
΀<�,�1)�p�m������y�5�E�,c��?�ԍs�ulx�E�-���[kw�5S ���n<�}��Zc׆Fm�b�5�S��X<.x�蛬�ߠ�o��8m_�~��$0��D���`V,EV�/N��(�)gaZ�f��FC��f��[6��A
>��c���J,W=A+�\�㯇�"qrv
���Z`�D51��;f�M��^�ޕ��+K���#�$m,z�7�ž�׹�7آVj4|��,2#B)N���W���ev�٦j���u�Z�n\��5��M�e/Db���Bݼ ���05_�H����)�{��+�j+Jq1�V�}�c,�ݴ�tF}#:���V��i�;��g�`���ae��E$�Pv�[�QQ@�"�Ar2L���+�����TL��2�¨%�}C������̱w0�W�-U�Y�sSv�_?��L�?s*���iu��6o����Ļ0��������6h��L�����~d)���9!7�izmA���s��b+��z2��K{���е@�M<�)��S� w%�s,���$�/bX���|�)={fx�S��v��fđ���/}���2�YM����d/�?�g$]!��^�G,d^�J'���
���0[���˕�P,V��s�j)T[vI��Y�ޔ��Qoib���ǻYd�Y��3���^2���B4�b�k�n3���#�"�X<�^A�x��p�#c�n��/�-�g���e�C�A����է^
@��1�� ��?�M���c'�&�Lx#:�%6��p�=��u�-_Œw��1�7_s~3�mg������oLKK��w�y�P�/�Vܹ��i��?��o�u�$T3t�7�L���P9�䙩�at���
���xC;zmQ̐*��9�ȵ�{M��?+�d�l��Dt��[C��q��Z�8�BĨ�dq����q��Y�m������Oa0!ڼ8 ������MP���bBaj�,㈼j�Ԃ]��Nm�B�"����gbX�
V�hG�(3],�� ��	1_:�'�Ekq��"s�e�?h֭ �:G_���x�`,�S'��!	J�� ��Ԇ������@��7
���68��V��	ߥM�ѿ0�0�u��4�j�z�~�"��Ù�F&�f^�u���/FU���е!ubo-ݧc�*���� 0!�xL������	˨�b*��e2�}t���5�̉����b��7���~��k0wL
��LV�X�+�����w-��䓛�OB9FU��hi�$j�'����7�����s��]�sQ>�8�q&Ș�ّ���g���`v�v+�ɑ�q#�}mP{�=�c�"O�>M�mhgs�:!�`L�N{D&oT���*�Ok��l������S?���� }�;ڂKD�UѼ�e[����^ p:{S���ڵ��h���O;�`�C.�T��ɍе?c��n���D�ve/
�J����(P���	A2���W�.�����Q��B�'���1Y�zZCBB��"�N,����fn����*�!Ayi��d�lE�(���@�Q��$rAȌ��1�{��o�F�r&� C�vfM�YBr��*�j��PZf��)l͍ �oU�1�d'"A���E��W'�)y�)yucXSM�5ٺ݋��Z,�����i����z�4�x[�)�=��m1���R	�u�u�`{C�$>{���l6�����
�,謤��g� g�Bz���-��,c}�3����-��1��b��*l��f�,�����]u���d�Z�T�a��)%���D7�tAO{�lx
{�:g��r4㝛ޑ�gd���o]l�&|nG2I�[@@��0{T*�]mT;�/����-�m9�Ȅp����|�t�#*��x[��-Z�<�����Rf�W�%�O���h����i�������J�زg�<�^��)x˨t��/筁��H��l����k�����Kf��?y"�.�#� Ѻ�+ù&�����Q>���D#^֫��A�E�]�n��n?o�vM����f̼�;y��T���('�I6 ��4LD����FA/�X�YF����~���^]��4�.H���ߞ�*�#��3ѵ9?`K�8Ւ�F�?�9���0v�4�I�8�@�\$��!��^ἧ���W�jtԯ*M7������%�7������#�[{jWy*R����*�*M�tׅ�v��?�u��N�JW�߲��2���O�[�/��,��?#)1�f�
#�j���ث���ʭR����q��t��)�)������˷%� ��%G���Fi�-��_�a��Ѡ�fK_�%@��i���I���ĝaf?�Eh7��G��{fA���9i������b�B�ʅY���4̓�o��$�S�l�fRrL�4k��Ȣ���6%:�P�!��x)A�?��>RJ��rx4P�g�e[#���qB��g�Y����?������~I�zH����и���]	�qc�>�v��/)�Lg����^�1Tx�����i���&�����.�g�s@ٱ�q20�0��1w����]����޳�7�>� }�Rfں����`�����N@'��������p� ݅5�eW�<��n�^ #N�gS8'�~�E2C:�GG�Ӌ?�L���!S�_�MʒZ*.$��)�I`�t�X�-� R��bҝMY�>hDOGs	�X���@�+� �����hH�H����1��!�����de�bR�O��}<�ו;�">hA| �����x���	ye�HɉӞ���o�t���L��=�X��p�i�����1q�\X!֘zY{Ě|{�~H�ޝ���6�v�� �xFƻ��4���N[NS��`���
 :�Gź�0/�s�;8������
)`8<=&)X�kۆ3���]Y��K���l[,�\#�f\/���c��u�����m�]�9&��H��m< �l���;B8&���#xBcX:;u؁k�&��U�{��/+nX�<f*=����_J��.��e~�X>~G:c�dM�+F��"#�2�՘=�1��}\��ɯ�t��ny+I��h0)���n�YO��͌w�o������>�'�g-�n0Z��3D�8��������4b��n���5�V�Mi}��Z�H��E�B�(�Χz�����tD~�p���u��]]-����ӄr���v��*7��_"GՉi�ZW���O�|�dҒw����T82��ϩi��:�^��{�ۣE�'_b��`�&�9���0"�RR�D��%1�؀�7SCc���<�R�*��@#i�i�����fϹ����#�Q�:#��n�� ,V�����i��y���)B��w�gk��^i�+��~ZBĻ�W����f�Ctd������ba���yR��U��.����b�������̫�R�"�5��E)9�5�J�	����[`�ݗ�YRV�A B!�o�7@%>��Y�?�7Ҁ��@�(]q��Jw��W�-5�2$U d��{��D (<ʎ��{4��f�	J��|���Ѝ2䩎�,����<Q�z��3ύ�_(�)�h1��5I*�y�_q�Xm��(t��8�?�[�:�҆�!dJ�;p���{����~ٹ㩞>���B5F"�� N..E��*�gg�������V`�K(H����IAr�3��m��*IIaF�^~%ad��K�6{2�sW�=���ӘJ_1,�zF�&��pK�-�?4��F�h�3�&�$$H*�<CHŘ�N�
ҍS�M?p�P\e�
V�or��Ќ�n:4T(����׹l@�*��ә9.8�T�9h�}[���f^҉$\4�/]7���8TʰTTP��,��C8���[�z���\�f^���Rذ�{[�w���͠A��Eu��(١|�MRFTWLO�
�A-��d�4����􊻝 qֵm��u�Y�9�&`�C���T휊MT��uZ���Ȩ|�)�
��Z���z�ealDM�ma��Y�Ў��q�4���m�r?������ćE�H�ˡۚp�?m�!.�30������[�RVf�vm������w�5�(�`�%=Q�N������W̷��:�nʀ>j錝�c�X�����+m
����������\.�ß/Ӯd+�T�C��(Юj��U�P�a�%{�+�,�����s
�R禀����ˠ7��i�_�J�IŴa jɽ�R^"�Z���GP�Y%���	�h�S��� �v��-�Q��R1�-S�lС�Y>������Ӧ�"@�^���TR��øA��z��"�1Z���_��i����S݊P�WU6������41=��J�%���g�$�l���ݍUF���A�B�)5 BZ���5&ؐ�X�e�+z�Ңk��+��x�R~���\�`M	�3<��"5�q�J}���7��m�([�ԗxn]����O?	�����,y��r;Q��0sO
5����#2����q<��U�[(��@���#F��2E`�i�"x���w
54w��}@:�h��ZAbWq�̉(<H�V4i:w\Q�a���u{a�Yk���n�Tme���b�X̭̉�`�e下}�K5(6Z;� Y��5/�(:]�k�)pJ�$�$��B#�em�'�>�)�s	+T$�Љ8Ԫ�h'�LZ����7Ş��U�(6��mH�&X�"&b��$���#^t�=�%��;k���m�F��^������Y(.!������E̲/�w�	D�p!W�O%z���=r��UI�mz�$5�&A��U���F�8�QV�h�$S�OPM�t��9�w�1C����>��u=��y;�5��y'�{ڽqE�T%�p�'jS}<]��" ���S�ԙ�A��������4�Jo��N��k|U|U�������`��g&y+�C����
�x<n�q�ŏ�~����[G��:!��ď�w�Sʴ�}D��n��r�a.I������Q�+��e���/����|L<Q�[�+H<F����鼇�L�D��2^�.�ə�ft�@9�eT6g��}Z {�w6Vۣ?�_�.�0h�j*�vV�Tw����Ѿ4��`ji.e,4���F����, �F-�Y�O����(t ����:(��c�C!:�HS��\�X��CЍĐFI�[��+XYF7����l%��ƇJs4cX G7p��1ң^Xѝv�����֌I��R`��U2
��̥�{m�/&�|�q��S�Z�+����gTk\߁<�;k@k2TȈ������.u3���z�2�2M^
�*d��4ϲ������4,�"Y^?��t0��E)��]���je�KÆ���}��ʔ?)T-�&F��t��o�;�(�
2*ُGR���IB��^~�̓y�����~�j�HZ-J�����c*��n�.*L�������tD�WN 5�,^u�������U��gujB�m�홋9��ѕ-���1�RvN���,������`9X����J���5�菃u �Dz��B����N��Ǝ�I6��RLVX����|@{��+��a��]�>�^Dz�:�,�i�䄬�f��|���pѧ׆'�{ z����-K��y�dOl���C�A�JV7�.����P�rԱ)�ŉ��������[*�w�֟�nd��F�3�l��^J�n>rx*�/�7
@�"�)��G(SD$b�n��l����;N��(�F��UTY2����246^�ǧ¿���^qNy8�B9���K�.Z�ۦ��3�(.�).������j�e#���%,��W2�n�0��O)FP�����'�Z�7�8t����u{�N��n�l�+iZ>�H쒱�������k�S�_��a^��mJ��rj�/"j������q����8����fY���#4c8>��� �k`sS��U�ce�wг6Ep:S��?Z��˪���c �)E�&���*"Ȑ��~W��Jاm���\��^|�m��sxX:�}�5�c�d�qz1�s��y<��(���J�D�%)�E�"@��`���kƍ��9�X[S�+���"�c��hOe��Q�
�{/O��SY �M�=ϵ�5����R��Q��V8[w��A�.���o�ŖS��(�����lvtxR�5�����ԣ�A����%��pNU��nT,:�����7�|���OCK]Ѹ�r��Y1i����������G���w��M=��Xba�r����%U��]�M׊�\��Eʐ^�s` y�fm�V������|�����nܥ�q�&W�R�q�ku�$-�*��,*�l ���/��}�QI|nz4�g��Qm9��%�B��a�f{�����3��R�j,a�:���z��s4!�qQS�Y��`�Oɷv�$2�Wǖb�G�I�ᄘ�@:b�T�2�O!G�{j�Fż�Yq[~:C�P��4�D���v^1�Ԫ �O�7�Gb �3��+��>S��K�5�ڂa��07��(����hh�4���<�j�%q�+М��i��L�sp��*��6?t*��v7ٓK��L�L��j�X3���-Ƚ�a3�@=�Ò�n�$�.n���GZ%�g.��S�e���Eq?
�J*5��M+�U%N��3�ΘH��q��%h���GY���n����))����>���x5qڂM�+L?Jٯ,|�H�N�}��#�襺y	٬�F*s神�����`���@���TvR�:�w���,��������bi]�B���d��Brz9�$`��0��t����>�]��W1��X�v	�Q�~�&�!-�/��>O�"����k�C�����K�@�����?���0^v�B֩�i����?y�v\�ߞ�_ő��	��1���v��~�	iՖ��nj�.�Z+��?�#<�Y*W��[�hz���;�����%����@KW�Q�*oDe+�r�yk����=V�	����)w9� ��;���&������e�U�9��(�tE�F�UY;$C��6a��;�6�7����o�@��45
]���4�)�;%}ӹ�`����+�j�zZ�T�7��"j��܋����7]Y�b?� C����up?-�dD�x�)St0;,{��8I����9���
��7{x�����4Ө���a2M������E�1� ���@��sx�Y�o�ȩ��֡�h�R���e�*'T��4ոjk�Z�j*��n�6��G��z�������o0���=����S>��$��o�+�OY�G�G7&���!���Au�pW���(�@��rE �\T�^���6-M�uq{|}H���ޚ��4e""F���~n��c�h�Cl�=�W-0ƭnE�tǁy֠G��J���-��tX�U�-��`�9��j���(���(��Q�ђ�o��}�0}j�+`��<cv˼B"��LR\��<���N
�+m������r}�� ŞY�����t ]���Pn�֜>s��	K��	5�Aч�D l!�zpa��´Y��A�`��?s�xڂ��R]ΤA��TK�V����@V��a!���25����NL;kFW��K-�[f0��g0(�)\F�x����W�t�_��^"���A����������<�0�d�r���&��t̑�`�x����k���JЬ�S��}@�����htjແ՛���j�4�W�����َ*�=NP,��TP�'�ຝ;S'�!�]y\��;P��%g��ϼGd.�k���A�J'oN�-z(t ̫��#U����,YЎ��S!_�DaR��k���i^/@��>V�b��'�R�'�83�v��ay��wM7&U̮xt�����S��5d3�u�[c�Rv欶�PG?��'���f���vn�3Ľ��,մT�������-{ԇ ���i�J9��Oq�h[d�m����W�:.�unB[�F�n+ͤ2P� ��1{�o�$/�0�\O���J��F�On�`�K�Ӷ�P�0���G	˽О��Ĵ�9P�?Nv?UҘ/��u�6!O�-���Ca���'�B��������M��c�n���=H�:��D�� z�|:.����@3OW�⪮R���	TJj>9���ĤG��r	<Ľ��xgv�z2��n���E�����z�#"j�{�= �W�������km)"u,_h���hSK^�%��k�x���Z�'K׈l!�[���a��!tV�L7Wy�ce��M���n}�b^|��H��b�0�Q��cu���?�͑����M��gpS�${�MpZ��/Ug���d`3�� ef?�7MZ-	�yyh&�_� �jM� ��#��s�6z(�+��Y���B>��|���Nx���V�CH?���/]���_��5�S�l�D�U=�DMv
(��p����᱿���|zLQ���c��#&�>Y1QI/��Z��*?ߌ���,0�ެљ�>O�[��AYb���뇷8m7�)�,|
���B��Fq����n��p5 Rlڤ�<�������X�44�Ɣ����hA�}1&�r�y�����a��~�����b]p`i9:q�i����	�p۲.h�o����M��p-���sG���u�Ƅv�33�4a����;B$%�ڟ�˔�dj&d���hG�)̅�s�ko�6��g���:�ϓJ�w¤��{�$�)�0�@��>5K3Jrr����ҏ3�1!21��{�Ro<i��}��<��wUI&u8ֶ��3d=�E��O�ř�9;`+':�R+�"� ��>h;6~s$,���爂���k�t�X�^YH,	I�A�7Ik%`�V2���!�!7�`X����8]K��.o�h��4⺖\���2&�S�T��h���.�k��0[sD��ilJك����Bd�5gq ,�(%$�c�oO�ɚ�ɡ�K
��[9DZ�����badż.9,گ4���I��y�A��B�P�W���]ʆ�	Ƴm q@�$��s�dX�ș~�<$�6ؾAn����P��U͵�8��
^��Y�sm��ވW�d;W_�[߬���օ�%l���s5]�S,���w������4���2���,D��Q�cb<1E�Cp<�=w)�=Y�$�A*��r6))�1�f�k�4�{����+i����QRbg�?E�퀦*�lHju��K�8�׿��m~l)-�ּ6�ߕ%t�V�Uaq�o�i$
��7r���YX��DV\��K��RoT"+V[��\MA����rIb~%BQ|	�r,�`�J`z���(�6�]G�N��Ψ��B��!��`�2y$~�������^c�JF|�N}��Jvbru4��E|�}��l]�6d�7��بLs�<;Gf Ȱ�MK��qX�<D��0����-l�Vۜ��)��[�l|Cki�?��ƥ��Mo
���S�x.Qκy"��0@G���(�yq�3�d���Qr��0U��8�<ԑ�h0H�T���9�eX���޽䨕ӫ���/��/k�[j�ӡ�wmS�������׋G��i��\�T��&�H�c"�7���87M���S?���D����C8�7���/zM���f�0�"k�7@/k5�-i�`�5�A�q�r�2��&�+�b������������㶸�\�9��#S��Ȩ����C���j�B�ey�C��^%��HY����s������a.|�aP^N��a�QNV<�v樂����2m�٠���#�xj�_経ޗ�������޼ �}�ˈ���,8�/��M�?�{����݅�v���C ��$LAd�E;c`����c��U
��~Z3܏b�g�]����;�d~��l�'�m�ϣzHÑ��R[J�v2d��F
Ս:#
��u��O���Ȳ#�C��Pr��5X�s�J>M�Kb���S� �_���fc��C�Ði�=��Z�ǰmKT����I�$�I�����i�Iŗ��:�4�����?�����j���1�W.n(��P V;�!��,o��<E���Nl����ƃ�� M���"�xᢧ)W�c�`|�ݘ�VWM��SA�R��y�l�K�#o�~� 4ı��Z q����Gݡo[Bu��N����=�S.r�PDڊ�>.*#�S�H+w�!�x�=L���\Jd'�Y�l���dH��%�.1�(h}l���o)j�o��&��c�ц�Q>�8�MUZ��cX���),� �<^d�k��
4�'��cU�D���F��S �5��~��A�w���
(��ܷ��O�Kf�B�PrioJW�-~����V����L���CX]|���=Bƈ�|Q@�3�`R���8H��re;0�M�썃C���p%�J"��:�����j�&'@$龡?���𪖊����z������3vxd�+8�J7,��S��kLZ��,*�(RY>�(�U�?��[�����pbp_�N��� (s��'�ߵ�-��%v�<3�ܺ̩4�$ʎY�C���D/�O�FW_�� ˿�����â��y�n���Qbѻ\�`������<��A�v�ށ<��dy��U������DE�Gg_8�i"s�f�u� /�%x��^��)�Ap��-�vr��_�����)��)P2r*	J")�?�e�Ip;G���R��v���,�z��'F��Ip)����v�2�&m��Ha"�L7�>���`�t�H\J{���M�QؔDQ���s:�HA�u��E:��4��E3D������M�
5-"t��S`�8㪣��Z��E�f����:y"(�檿�h�\~k3��S?0�2��ߙ�6~�&�/9 ���š�j�[�\Q	��u�?����r���R���F���h�	PG.C���61�*	c����a��.a����^�ApzMC�r�Xc�����G��j�د�����SzU��pE��5������Q!����G����r�u��A�˝�\1�.�� a�����E �^E)ҳ�^�ћ�.��VU�����_门z��<��߃+_��on��A"��M��4�m�v���UQ-����i@a��3��N�[YA�yO$�'t��Nh�B@�NM�f�#���O�VGS�*��l����SN;�طA��Z M�lzd�<0�����	�X��bSۡ�bC�5G�8"Eʵ�bE�yQ����9��J�;Q�c�H�żN�F��;��܆Y��ij�0�;�� �wl���$����!��u�V�kx���K��s�I��t �:�x`u��[��Ǳs�p�^>Ʈ' �t���§��p��싮�b�c�p��B\y�Q�� ���dn�ϥ`{�|��W��|�Y�ꕟk�Wi��%�T������lF�#Z��_��:�ֶ����&�:�M�L�L�HS�����h�0��ÏŴ��6��n���b{��������&>CQ���h���۱�%���@N`�&:��{���N��XÄ2�@��KhG�"���A�b��3���v]�.
�b?W��������=��}ܬ�Qd�8�Y�� �x,��������9�H�.`4B�� ���E*޻����߂N��t1�由�Їf�df)E�r���<HnGT�X��,�B�T�F�D�I�iSG�(�k!}����i]Pd_���nޒ
����kS�,j�CK�5�U�k�^>�ǘ-@���f[�؈�� ���sKB��1�?�z��v��el��3d� ���Q�<&M��됤��_e����"��ӐB�O����,W���y_�z�}��B1�[��*=��v��eI�q��u�V?>sq�p�IR��_&r��,Ue�ŴzQ��\�4����T�*�^X��T/5&��V'�?ā�������>��2&YXQͨj���A��=UE���[�g�K�M���_�M��OL�X������΋��'0=���+����:���]_��+:�Ls�[޾�X�1����h�����*�D�n��$|%�+���J7�%�����V��d��MM{ۀ���5+	vU���E�r�_C����=���zUƄ��|	u�5�D�I V;�_ߣ���'^��6�m�Q�@���xH�Y�cS�e�)�E�ۅ�
#���XF��L�ے�B�-����h(��ͱ���'w�>ƫk�[&��**6�1V��6C�Ӎ&�c�[�Wg���&�� ��j���� x�b���Oo1ҥ���}:V��[�>)ؔ��9���-�<js�#��[[�r[Q��L�if����z0�`���9E�����bF��I �&&�99��PϬ!n���Ks#Q{�<���닩Ñ����)F�LB�UƾM	L�+��߹N�ku��3�R|/k �޶���\��2�H�}��>o	o`��S�T���r��Pd#�zd��z�5c�`W��Rt��?��n-���Hw�X�n�i�����/��D7�(��,-�̝Q�)9Z��W��`5]e�3JQ�M��H\��궴[�V�������=h
�(f"S�]�4
���Ǟ��~�������ɀ��\��`���u$�~!4�gM\?2�`_bzf|�(��K��^��:l�Z�7�iݗ?V�|�	b�Ӣ�W+L���O�z,���j2f?�``�Ċ��v)�8���Xf��mk
~UZ�Ӑ��'#�,�=y:E�D
(`�Ӥ��o���O�W���	dj�AE���`s�@���j�,�k"y�IR�AW :j* �k���� �*Ъ����y	��T���0H��a����ֲ��ϊT@�TN�`�kk@��N̟ΈV��g_�Or=�sk�_�,<���).FdB��C��YB��6��y��8�淚�Da�Q,�_S�ίt���.��I�����<v`f�v�G��0V�7!�
�ʚ�J��?&�v�UF�J�d1R�"���w���[���w IY��
!BA<3�o��/f����6����l��b%���GEl"ƶ�5��Zl��ئ��	qL��� A�i`*��t�o,��AڔE��0淴�*�m��֘�U��pQ���B��J�G':Tv"f����WR����$/^@-�۽Jc�fv�'��3�kM�Rp=����\��k�xB�@��7&����-_\�a����]ҳs
�zҺ7����u�$E'�j��
���l���P�$�{�=?���w�y����]Q���!0%�d F�ԩ8�;���	R������g��\޻�k��c����IфV�,زs����!'q�>ڐ�Vp�2/�UF@^8�A�q&x���*��Z�#��_xN�yM�;D�ܪ��=fFT�����27���qK�^� $�l��x�;'<�E ��%�0�P�Y*lJ��(����m1ޫ��c>��L�UK��97bV.����ym[���d{D?����./s�?~,�0�R�Ƚؗb3�("ׁ]y��2rߘ&*�/<-�|�e��A�u�%�
uK��'9bb���%�^m���Ѵ� ����啰|1�2���ך��zD��6�� ����oE�cg��}�Dw{(�SH�y0��RvA�=�Y1Y�݅�ĝF�Ƌc�=
���pE���ݫuZ���L ��R|��&�#����9��5�)w�g �ϫ�˼� RC�h����=������C�헀�I�h����E�cjD�L"�o�zgt`�!|(���(���8����pb/���@�C`�d1O�����j 6s��+j��X-�v�oQ+pCv�Q�N�Q�>|2=J:v���E����f�O�v�L\#q:+�a��}���2p�v�q�oc~+�Haw���ccy.r%<���W�%���������-�23�p�`�k��i���Ӄ[པ^O��PI���w��E�@�r6�BW�ơ�����Ӝ��I�{��P��?.D��L����&�ǈ<��~������9C�hܚpL�m�x\<2�6� Zg�^ٺ9�
:0b���sf���t�۳�Ǆ��o.���@rz�f�D���N\u�Da]2ׂ4����ˣU�V�FĎ_�4H��`W-�@<KI�'��LıJ���X�4�M׹�Z�>n�4Q�m��'��Y�~�(&ϨU�M#�����v{H�������I�'��OP9�L��Y*��E~r{�t���'���2�U��N�^��=�h����?�#{`������f�?r��[�b�FA�ڽ^󦒉������O�,��%53-�Vw@Wr�󠁒q@�v��p�3v($�P#�I�jDm�}(u��e����[���"�!�0�8>� K��#�L㟛�ɇ� ��:�'F	\{ P���g��4M�PH,��ٹ^b�x]�=
��P�~�
��V���Z~������q�Z���c $�r�ħ�i�0�_�d�B���#}�}$��X��=<�"�4U�^We�X��)c���忾Prn�*����gu��Ĕp�{?���&衢��&� F��������䥔W᧯� ���^�4�/���갈X���[4R�>Afi�,�̠7�X��'a��&�j�O���-�%(��$3�U�x1�
7vj��n��h|)����Y@w&��Y���CtR�cIR�>(�d�t��Av#g}
'Ʈ�Ə�����&�����fֈ�͑|�yC��ݭ"m���`T�.rT�I�s�o:��s�JW&ց	��b	�w"
�e�J���:
@����܉q�9_#�m8�	"[�m4BkFd{E��mН!����ꍼ����,����4��U��͢�ӷxEXł�kzZ!��0��:բ*�8׃��S/<3�b����YG@��_ﾇ�$M}���B1ׇ7����k�$Wfr_�DyH�(�<�^2m��}����m.&l`�)��]<J*'��2�I�Mq�� D�Xp�?	�R;�U��OLW��>���o]f��OQ���4�7��S?��s�Z�(��/Q�b��Σ�%��X/B�R�;��e1�	�{L�u��Ǘ�dW�SX�kv%����H�S��e��OD>YӨy�2��A�z�+����ǻ�Jd�)*Hy�h)j��a)��{^�@Kz�H�q�OhNj�菉���ے[3��]�e'3�L�ţ�9���H����8�G�>��s��R��T�ɽ��S�D�L��:ۦ3��]��
�op�^��o�Wbb�f9s��'��kkr�F;;o���Ղ�N�N��<���V�YAN�S6`�����W����}(���! �c��]�s�%O����o��L�u�=�XZ��>'�<$2�����19��I
����T�W��5�
�@;_�"ti���t�D�T�� 'bEeft^�D)U�:�D����e�F"DZ�F&wK��r�̂����I�h�gYX��)��
�h��F��D�4O���{��ia���|���Soˡz��N��� ��L{Ľ�D�S�#`||���XԺ�g��k��?y���Ӵy0iP.�."o6��%��Vuԙ�����d���D��RЬ6E70��ف��֟��w��x��;q���4�[>�"�ic�V8�/�eQ=�B73�˹퀱iY8�jv��	��.��=�k� ����^��F�����rM�S�g�=t����6�=�T7@���Sy٬�d����s����%K8�(��K�Ȃ�O@w�T+��{�v�G~u80R�'����G���0^u��[Yh�o��1�h.��"Y[�!�o5Z0@}�]`��w���ʹ0�����K|�,�-�q�˶��^M�,9e�P�Ԫ3�M�$�%Ao{�o�t�v�1a6Tn+�29����g�=:ӂ`�^)����s��?�*A� �^�� �Z�G;i4��������vu��zA�T�Ɇ�R4{z�8ԢMS�T�}��}�:�NyI`�n�+��2I@VV�=
:֝�8�V[A�Iq����t�������sh,Ϧr����J��#��Y@I�Xb_t��:V�S��L4,�����Nk��w(��թ;�	bXx�Ͱ�I~�S3;������'��bCn`�ntgL�r.����?����
���Ũ��A�)k^� ]�6R1>B���:t+�@����߱�����i��`!:F'	N�˳8�3,bf��U�u憴�)��\�Xt���E������������
�*�k��Y��F�AZ 4۱�'p���yx8ÀaH�,<~_���Y�ڐ��KA��*p��ϧ�#'+r���ŕ�t�I�t8��,'~\u9�Ω������Gˍ:��y	�"8�<�Bc0+����u)��NT8J~�E�]=��i���<C��.v��Ӕ*�N�z��*2藰P��/�i���H�^L�}�D`�9?�=<�©k[U�D'EƟ@�*�7_7�tv0���Øk[ns��1RLcr�b���?�#)f0�.l7NgO����/Ω��������;Gl{?&��l��Y��r��l6��Xc,�:��T}��t,.�:`���<t�T�0:J��J>>�/�C6�䱤D��h���H�)<���P&,��C׀�V�c��G� P���G\��A�z ���&���ZS@D`$-��n����~(,1\�Q�!_@�a�8�g����=p�+�9eK�d?V�j�z"�w_��@K��IIr"�) �ަG�H�s�Ǽ;�˴����B�G��lAns^�c2�8���s�huS��n5o�F�|�ZϝZ�I�N��<�,�L�ܳ�JK"���4��F%$�I5�{���rY��ŏ"��=_z'^a�d���^zW�M��uQv���(��j䑟j�3�_Y�AQ�!�`(�L���t��Ͱy3���J �~��������{�=-'�,�������u�b�I��80BԴ�>��X�wr#�d�Bm�Ij�ʄ9����3��"k���~���������rXPr�p4,8����}���JU�D�R��t� q�fR�����>ވ̑�ݻ���kڠA�c3���]ZX�+�cߓ=�IKW��=�|K��CP�!Q�K6�rj�`���w�u��x>?b���>Q�"o��z���8��8ˏ=Y�؆Q֙P�B��w���ⱗ��	N���8��,���sѳ��é�I�EB1�Mb��ۊ�2��LmnW,^Ps��{�Xf�B���#�>Á�W"Ae���]D8����F���b�1�/@S �XHF�[��Ƭ1�����[��LapGӐ�>�ZS89����$��W�j
�����Fk����;���t-k]�y,�Z��'�b�εn����\I5{�u*��ӞG*��o�2 l )������;�]�;G�I���]�<�6Y�w�������ݪ��@�2{���6*Z����T.�����5��+����@��  8��'�]w�&y�d��UP�da�ܢ���8��t<tL��L�N�l�G��ňi��dc���H*
/�[z�Wob�5e�Je���a/�낉��6�(�:1Ē�jg�_��s�|?�D���M�eZ�D�WoYs���n�`U��Υ�t��&��"M�a�N�&�Ĝ��ţ�uS,��^���4��HAmbc	l%Bm�@RCA9g_������W��i��	�mN���ZK&�|CB,�}�ж���
����R��vH
=G��M����!|JJ|����(�R�����o��{�g	�^����X@��B�1�>��	A�!�B���ܜ#�"O �z����aA���R�T��Q+P�0���ʛ��l�}y��@^6�X�����]������p��'7�������Liw聄xI�d��v�($7Mwʾ5��`#*�i~���>f�,�{����j�XW���~���avH�2�a Bu�B��	1832^����Y\7ٰ(�8k�G�v����FBH������_ԗ"�+cC���W�Y�h՞O��خ�xw� ��)�CD��&�X*�'�]Ԥh�ԩ|������� s!��j`!E� ��>�.C"&o�ӹP�t�ZMwv����QO����f�[���j��"�U�������9ԺCz�I����g=f��]�I�x�.�ǰd�A�s��E@L�����[��ۯֽ�TZ$ه������p����Ĩ�������Y�n��ŃQ����8��'m1�����Y�����~Ւo���Ku=�eY�:?���i�@Wx�l��v	ݨ�pRUP{惲X7N��+�?+7���TH�T�JI=�}Y����rq`��rhz&�� �1�\L2��?��R٣f]�V,�?��<z���)�\vK�=�A,�8ߖ�ra">���%jS�S��
��͞ϧ^�'B�z���$�jb�F�3��|��˫���h@�Oܭ��(PZua���V"��mZ�٩���]����sެc��B-�����=^Ķm��2����p��T�n��|L~�[��O�.�06(,���̵�k&��xS��ᒰؗ����l9�c������W����6��qR0ik0ȭ�}����n,�R:�j�z��i�u��k��ƚ��y��I��R�n�kjuŻkߺ��e8���OW�<��9X��.m��'�_��oD�Pr` Oid��B�Fj�@vNS�R�a*�P;:����OkU%�)�b�������)���Y�2��C[��)����=�[0���I���y� 54���g�����Ժ5]��Q����-�y
dV���2�6��L)��ȳ��`�k�A�u�&W�[;��E%&.����m���{�Z�q�
鑇eK؋�{�����.���D�U���G!�����*�g(cB¦&)Hy�&�ls]�d�4x��B�܎�II�wg���<� �A!����Q.}�'�UP��S,.la���|�
CQ�	E-����=��FG��h*��Ǐ�9	�T�߁D��:� 0���M ��8b����E��g�qBn.�cj��[�լ����*�Q[3���EK�@� n��������mC���P�D�0�R	�^��
���k��y�I���X�ʈDWn��p�IL�%�+<E��kM���^�=���=i���ԡ6w���jь%w���|��A�`� c�'�,u�1%��4���w��K�	��t(��`�Q"�F�#��=�ά��;�.o*�X�<Y��?�ua�]v���[�x�����p2�,�{�Ц"�%��D��*r��[��c����TTJ��z�J@�V�c����<��yj��9ֻ�֊^�_M?,o��t%�#��l�q��_����͹���2O\=$3Nk7�V��)�H�V�8O�F����*�c�Ŷ��;Ahۓ�N"���!;�S��pT�-�T�6r�i�X���$L~�����\Dru�P�^�ߘ3���q�"HU�L�`�q�'pG�;��s�\$-��(�7����ُY�icM{��ȻT��v�/���X�sR��P�FC����$�ı�3'�ڦ��!�^#�_m��n�ӎ9Zh�++�xi��[�\s�wp�]J4���͸@�C78U�j\#BsYCW�d�Ǐ���K?�}�^3�D�b�iy�2�Qe���.`���mm����Ky�?��A�R�&��=�m+��Z"OBـ�;��+�h�����B���k>PÅk��c���)�]������&��N��9m�(e���݅x�
 9F��B��t��no(8�<��k�3 �*��8���6m�q[tm�C0���U]���.��VA�

%|P��E��\i��A����Q��IR[�Ow����:�3����b��)�W�\�'&-N6.��gm!j��ͿO0�%S��b1�K%����e�?�+���]�����ԇ��y`���u|X8�^G�"�u �!u�D�k��v)0k�hn�q����@{_�i�E��<�	�U�f���T�b��q�u
��=Zi�?��U��Q�e7I5O�V�2u~ ���Wpڏ��M��6��=;�=�!��{A�*Q�ZH̏&���[n[����Q�\�� ]0�yPJ8�nL�!�a����A�F0�
v��B�V��vV�����W��hb@脃�'ɮ��D�q����$}ph���@��L\����Z-䉭H��_���\Zc4�O����̞x�cT�j�Q�Y"���ZD{LvW�g��W��D���楺I��|�٘�Xr��'#t��/�e�TXh���ĪT�\	�Wa/���/GI����a�3t�Ḃ�&@�_���l;!�����pZy�}N9�$i���
�����\M5!f.o���8C+yנ��~`7hf%���!u[��=�h�	�����Н�SZ��j�V��K�c6n�P��#F���N�B�i��������߮W�.ZP����hNhj�id�q��ĳ�cն���S1�F��������@�%�Dx:)ze����4#1�L��-���Rŧ�x����s�Rx�dت4���qV��(��Xm��^n<���@z�
+��ir&S�����!��@�R�G���3��G�ك��Y_�*/�|�MZ>0�\o�}0;�o���	V<mf>�1,��T��J>��2���=�ݿ����ȓ'�5Kјᾩ=c&��$�%a���-l�.7�]q����Ŝz=	qJ��2���K�sC�ێ �ɬ4������	���z����$&�C	I,�E)I𚡩I�ap�_�]�~k��hm�ʸ]���VH�	��p
!k"fr��p�Q�=-��x����Kr����f�Z��{ʦ꠯�Ndא_���Z��y���j@��S��j�9�A*pI� ���O�t��ʞ�ޯ��ײ>��Jơ�"��w-��Q�}��G�Yۡ�|_���41Ǵ&���C�=|�r�܍ſn�`=RU���b��uzj,��m��Y��K�*-m�[�iriM&��|���L
c��<��3�W�`�	�}���tC�� �	��2Qc�xFo����qyJ�{��gb
�ʌv��m��1o~�l˝�W�{�
�،R˫��jzĐ����2�	�3\U�|z���꯫����CJκ�Aڡ�{܃(9�'jPG�� ��YW�ˁr���>v`Y�F��|S3��x�q�z�%9*5Q;S~`�Ԡ��s]&9M��:ې��'f���eA��eձ�u��ՙ B?@�Ϭ}�u@�5^m���Hp��7�Q�kL��+;X�������>IVr���(3M�����!��zSv�K-']��0���.�e*��U�׶�߳j_��ǹ���<fo�]����mt_[N'��� (�?#�J6�m�20��mQf�X�7��9B_�J\P�,Ҥ�l��#�"�_Z��i1��i� m�F���N��W���s�}���6 �*=AH�5�nmeE8��O\��p�N;jM&�x�N0�3e����	^@�2Z��}������'#����Ye��Hl�h���['�[d0�0�4/Jg�,�SFW�Uk��J(jh��>��p���@�F����ӍY��[�(���_'��0��u�3�.��<f���π�c"f�h�פ��5�S�6@z�@��a��G���Q"*&�k��x<A�8Yy��9�Yf,�aڗ��2�?r��Ho��:�~%�w�@�/&�A>-�d֚�f��!��>S�W	��VSt�o}�L�������H�u�j��`@��x�mdu+����x�8�ٷ�f���c'~����6�M%]�CQ%+�^8C�F{7�{ߞJ"�˻O��㩩]!_������q ~Umj�.ۃ��e�t�yL�C�p�}�� m1ܐ���r��#瓽����Z6x���qd���5]�!�)���Z���V�hnT��8Fܙm�W!���'�T�C�x�����Q�F� 38�bϤb{d3��U��զ&�Fy�I��5"o�*�e���d
�ݨ`I;l	iMɻ����,���*<��s�����v�=Q_#J�#��=�jy����Oɲ���Kx��o�\ovg�Z����t�I~9�L/P�����7ζr��	(�ty�,̸�f��fI@J}�ම!����Yp���O�Fz��kY��!�`%M96��l!���9(<����BW���ܷD��9��3U�i����c�,�������"�p��_�_X��P&Y��_��q
Gè� �~�d���*"f_��	�kt#��'�}Ol9$M�z��ߘN<l�6�˖Fy^���y5H���M�0�
L�"��GW�{�r���w��l/�x���(��ّp��P���FZo�ؓ۰��ʖ��ڕ*��g��N]��)�I9ґyTʋ)�5���,�
W��{�$�CL�əC�q�*�֠1����?�=��rI��2~#l�Ew͒�S4+��@���)ڪ�/G�x�5S2���!E�x��I��I��x��(��^�o�#S>�R�u~�k>��7%��{>���<�7qr.����:�m�v��gع�c(��en[���-�dM޽� H�����/�˺���ݴ�&Q>Ɲoe�1���P
>��"j�߁�!���Z��O�tPo��|1�R��e��З0X�ݑ�Y�i��D`JZ^��9�8=-C��E>�Ӷ���0J�`���V���1�����ʜ&-Lp��Wq�o�k����I�[}JJ����E���y�FV1?��r�X�ᓗ�8X)J�颞w�~t}�2O�(��>�6۠�D�k���a'�3=j���
�|��u���������yh�ڡ��w�ɝ,,ܚ@5[�o�p4�$��̱:��v������w��I���(�#��Ȇê��h���Qr����?DX���wx��G��f*{Q��;a���L<0A�a��;V�T�Ba�<�2��g�!o^�I϶s�?��:H�R�W�?�#�4��3U��Z.�9.B��K�X[|'����tՄ"�C&ZQ5sK�O��}~��O�R"Mo]k��	�mg	��] ��'�J�U�Uv�����.�쇿�=`W�v�l����P��cPRa�7�Ν)9u'�����H�׈ �e؛��{�����e/��y��-�e�EF�Y����>������7ç��G���2���͸�z�m��WU����C�L5���e�ӓ��ތ�$;� xaсFZM�7�pg�$����Ӡ�@=���JZ�H���#��3Z��ק8`iZ��F�47�{ǜ�b_�۷���#��[7�=@p��*5���,S�� �c&> ����A1�)�2>�nu߁�+�i���^�v.~�Hz�ݶ�ƛi͜��c`�`v�tt8{b��J�n�e�<=�Y��Ԫe����;|h�KS�>���L�}��]�����ǜ��FnF�����	��W�������<k05��y7q�Au��Z�]x_aF0��4Z����.�s���7K�Z�T�%��JN.Lp��&��J�����!��`�&��Vk��#l�a�HM�*��"��FFDc�g������,2����JtX����@���Ci���|�m����(�?�g����,z�[@�$q�EK�E(H*�&�9;S�`|C9Pƹ9}������B^t���0>Ϥ?��3KW�X�H��ǁ�� ��c���l�����=�����h�2�m��c�!Z*�aaN��f�v2uF�I�T�!^A�`������on*�٫[
`6:-aK�Q�������d��H�w)tϩ����GUrJԒ���1��X.�6GI�&�������Zi%�(ѶQ"΂?m�U���j�(���a�����_�W����7���Ϋ�d4k��l#�m�C��5��>T�3�2���&�,--}1��LNOw!'�b�z�^N,�.�n0_���GZ�"��bQ�ia�x󈏒�}��t{��!��8��S��U����H�Xrw��#Q��[0���S#Hج�-�:�q������{^���YY�$��f���g)06�����@�8b�H�'M ��?���LK��Ĩ�"f���X����-�y������A�S?d�D�I�H@G*|]�ޡ�K����
�����ۓ�ή��'�*RPެ�����ǟ���t��Ki��H���"?��}�O-�{G�M�e�LQ�(}��{� 1����lQn�x���s+O㷯���Z,U칶6ўs��E�K��!��:�iH�E��T-Ƅ'���D���~}�
����`^����ˉɤo�N��M�G|�j����Y��&>t���)+�m~��ҽrє��'[q� fi�b߆J���߻;#GF�Un%x�^��9`~�j���J��5@���h�k<.�Cɥ\pܼ�*�;}�B ��=T��+qG;���F�n�mN��F�w��XͿh^a�W#V�)y�ΨW:
�!�ՠ6�)�"�B���E����#�k���\W��t�&GDW����k���v�Y
<��,���:$L
�X�N�֙�ǠK����E���V��UE�����9�6�	��?��[�_��:sA�~��Zť�˼���v�#o�-��2���qэ��2ťzl�o�u>�4_���רB���K���<��G�j�d��T��)��k�Ԇ;Y�r����4%������m�Ĝ��e���:a�S��&�g&���c�M�j�=Ι�h�Z�Kj�21�Ǣ�D�▱��A�-Lwh���<��"qGCB��.������:AR�G'�6b�Ack�IYx��a��n:�M;B������/���3<i�����w^��d����[ �0����:�Ƞ��$��:;�tl��Ѕ�ﶤ!_9	��S���hu�ȣ
R��eCI��n}�s�6�g�V��Q���x��[�0��`�UlF��"1#~�z��Q���Z�>����� =�[�1!�py!�RZs��#�avL�F���Q5[/�ns����Z��ع�D�i��{�d�D� Rk T��M��/A{�U�|k�XG�%)�PBEх���t���V�n*}��S�����%H"5Tԛo� Z����c��,-Ѷ��l��^an_-3��*���������
�獋A�#V@�A�$h'��.�2q-��ou`�"�1�|�F�	+����!mJ�Xp�j��&K���cGv�����Sу�E��^(���9o�p8��,�G���%l��[jn�V��9�j�D�+�G(H�`*��U�c�eo�A�
��S����6m		���띑._4�S9G�����UX�W�.=��_��L�Rgz�@�u����j��ł��Z@fW�Kn���ï+!�}��]� �SB��S0�# ^�}����3)E�W�mRL0cM�׊;#/����x1{_����9���gM��N��ը x¸g�|����O9d�i��1$5��z�x4KMǁ��s���c��}[$�)g��`8����b��Q��3L�󌶑)�ҎRo�xS�wIgG�[T����r�ð���*?�� J��&�,��]u9��g�ke�"�K�p�l|���]���Tqd3P�K��⅛�����5j����xeR�[|b�cja�G�
�H���H�r��|8J�?G�
#'�EǂX�[θ�pdyתw�PVu5��֨n0�Fk�2�u���lU���V�`-dʮ�����������c�L�%Z:Eo��w���D��ѡ��`@.�Nꫂێឰ�.�W(�z��*�6Rשc���
L�8̘~��_�3��\j�:k��3S���.��^����o����Z����>>��\&7�8�Vd����B�<�b�@�_]���!P�jqU[��~}	+�>�@�fc;R,�/u��:�����V�ݽg�r1t�r�\Z$�^AeiQ�P����5A�s��X�����c9 v�11� M�͋�ȴy����9̫�#�9�d�ꈵ��C�}+�oT|V�EJ�� 
�aC�[��ݜ���Δ��p_DΟh�2��z�z���WKɁxF��y Q�v7*Ź���6|\O�1����ޡ���MX��'e����~��t'�t�87��e�`-���
d ��'VơG�k������5P�繛&�m�(	�]�,�@�X�y��4J�R�uķ�zQ��Å�X]��qm�Q4/�����B�~o�K�� �������"�~���>������t�ڕ�v�k��Djj�Y���Wp����Iz|!)1����I��\c|�>㱅fz~�<�3��$b;l'�����5z�`J$U��ƕ՜�E�Y$w�#�
�vO뀴�?����@��I)Y북Qe�|�á��� dG��ˍ�!�/�o�����$�U��"�	����˄�F'��̈��,���劥i���Ԉ����Ws2c�G�������rq�c�m�j����a�$�� W���y[����k��t*�A<(��������m��������9fi����Q��(���ZӲ(J�ڐ�!NW��mZ0�t�}��D�Eސv6Dr��Sc��f/U��,��).؞xY�����E!��np_E����7ܣ�<3���2P���J�3̡��|
��̀�E����p�fո���:S����c+(��:^M�ڴOM�YJ���ۃ��xh�����QBQ�nk�@(
�_?h���$�X��~TQu ��B��9
��ZY���݌MA��*8B!��fve�V���Y��O2)Sag�D����on���f�vg�]O3���h��Y���v[�!!# &���Z��=7�Xܩp�J��sc����F���^��3v�1=A����{� |4P��^'�(��Mdv�|K>��7R���_u�V��%����^��h�;7�Z	#�W7��u�3O� F�#i��፟p�-�=�
�����<�����~<�����{�̀B���m��_�>yK�^�y�g�0E��MX �no
o�IY�/�=����{��W�(�~�xZ�Il�<�&��C?�ML���'�z(�x��2C��?h&!c�{���s�Bͣ�I�K�8N?�����a�?���p5H�i64?��oo���س~*���"�8U}<��j�W]8���lу�$�1��Ves�R�"+Lƕ��`?m�>������7����o]��p����[�oL�D�������8���JfwF�1��f���|���4dA7T�o�+�IV�q$���K�HT�F�F���& ��5�z���ϋ<u� cd�f����Ӈ}����:��xx-���p���|�}X�Z}{ܪ�l���w4�G2<���V��
�*?��
�i�x�<�7ߏ���
��r uG	���\c�f�K!}tf]@�ܻ��E��w���5M�f��E�ߓ6A���ܚQ|������_=���A)߽���(���%Kv_?��p��첬��yΪm٩ל�߲;�;$ى���IՁ��"���ף � =�`�\��NƼH��xP���Ზ�pk� �س^��1m�u��5���&ӧ�C|2�4�C���"eL\Y)�
�Gß.	�!pɇ�I#
hW ��1��]��3S��>x2|v�_�P���/r�/N�b�o�	��PDB��Jw�o$[������6S�ɵ!��Z<����g�ʿ{-�[��.L4O�[1-�v���*����aS`8�nކ��%�< IbH�J\�v�����J����w���AB�Ǡ��vxl��W�J���џ�B�Q�"i;B�,v�Nf���4���_��fJ$*�g��p	.�����ͺҟ�\N��A�2/�V�
��\�wK�.yԎ�N�|i�a{�Cm��u���o2��h�ҥ��?r�>v�b�z��c��l~J��:9�`?h������0d�hCist4�b�<-\"�fE�2���7��Y*`��Q�cq�v0~�؁M��3�q�hY}*��W"o����r�`C2Y|��zwm���[�B�VGR�آxN%{d�N��G衘c�`T�7-�*�����i���B"�eC)�cN:[Go��,J�er7�[ca�i���blf��#aıi�_��ʑ�@Bq�"d���r?��l0��z
rF�T빼��!%�;e� ��o�~�Um���v����] w�L_�@ZA��E��O$[��
�!6�̝�Of�G{�.<cI�ArOkα3�|�(7ȏj�E[0����+?�N��V9�b�KcdM��h@9���]�I�,�eix�B��L�
xCGq)J�*�)*�D����M���/b�?9Y!$B��ʒeO��Os!���t
�Y��ld���k�K�&<���դ*�#'y�3DA��=%!tF("��'��I���(�!�oB�q?�<���[G�A�8
���lη�J���_[�5�yZ<F�ԫ~���TS����|Z3�q����Wļd8w�����C���6�|�8��G���/��2�/?��� ���à#դ�Y�BI`�Ϻ���Ɩ#�Q�RPw�}��◥-�N��k`%�����-�\�6��a����4+�k������2pq��S�����/�[��Wr�8*ߟ0@dkg/�!���X�<�Gv@����&�[c�� �0|��<=�
p�@���H^9د�� ^��k,69�5qNH.����_���B�on���#ԑ�� V��^�iX�^���g7�6�\��6dw)?�vnU�0���qt�ɒ�*�E/�"���+B����y�(--���4�>39"�����1lB����B�c]t͇�P�JJ�{� �$�xhh�� &�{�<���j�r�vW_i�@�i��|�_��V��y����a`�w�����G��\��Q�식u{*��r��Q�*�y��$�?2�-�s`�8��v?4�򸛎��î��R�@1�M4ź^xR���z۹�"�q�Vf�콼�������A�Bף���>�a�^?=�e�&9�c��Zy�
c=7���_[�~e��d��?�t�`�ePe~
!��1.�̷Q���S M��W���#�$�#h��/�e{}�-�d�M��1��d#!���ɛ$�#9���9�[O��Fl෱���b^R���R�����G![���EA6���>g]��!����L\�H�!Zy�0_����>0���Mm����& �_�k�6p&�O&�UX�XB�'��4��*��+�'ayn�ٖȾ�����J�]�])��U*o��>�֭F|�V	��$O,CA.���\G5�g�:e5H�9��[k
�,��7�7F���途�)��3b����:􉃼w՝�X!fNJ���Iцӄ]Y���C��$��"��R�%�t�5�!죨QU_	� ��S���t�����
�v��[���ܯ}�� >|S����o�^��#60��V��n�O�� ".�TM%��*����\d^|=�Vzf_���mz���{ʈd3��}�zx�*�U3��om_�BH�����Ǌ��� �:Ƹ�x�y���Y���턭�L�i�qQw���YTR�9� �6�6�^�3��s#n�,��+'1��|EU�6R� ^�I��H����0u�6̓���#3�����/�mՙ�?w,C��Y1���������GK�n~[�M�ޚn��6�:Ҽ��S4
��'���j��]�ϣ駓���~Ե�q,,	�F��L�Vv�\��}e׆$��>	��U ���k�\�/1Xe7�wF�EC��ui�?PPP7I0��T�/u�}��/��:ȿ��ٻ&#� j��O�h�q��s8v���֜����Iy��=��T��h�Iǃ��tX��hf�H���B޿e�zY�N�6H�Ou/,�t�m�Z�"����ePD�e�	B9�ʃ�E�mj��w�J�к�Y��ǉa/�G�L�Wm�߹���ǋ2�/���}��x�6Y1�pV�|T�/����z�ծ�߼�d��_��c��	/g���  ��ùj'ΉM���^�,�����p�Jߡ>0`
�i��>��=`YK������ͷP�t����]�����u���v�/�u�֝nJ蓕�k���Y��E��G��{ �����GWx}��,k�`��/������u+��k΂�_����wBZ��ԙ.9:�Y㵭�թ6��n]��d;��AH��i�v�P��g��y�
��q���k�����=x��`nq~�`P��_[�Ң�E0Y��y$�Σ2.�إA!X~�D�G.R�� ��[V�6?K����W�ܖ%�<���M~��W*
pT��QX!�����������#TН-�LBu�3��6t��|î>z�������R�Q2_3=<�����kA����K�/�f~�JYȞ���*)�"9B%{��M��R�?l�ۭ�!1hT:�h�a�.�������u��.�ejh�j�A:'�~E��Sd>�EQ��B���0c$�R��Z87�3����".��C�9�����ۜz�<��Ƿ9ݦ�����"|T��dB/��dVZll���ԝj�M�]�.��#�@8�7EV�?����K��Ϡh���Lp�]���nt�Eq%�x&�/�'#�S��:NSV�TT=*��x;s��.ِ�\�:;Ǵ]K����6|�-��{-���'�ib#$UNd�~ >�,�������Q�af�|���<*[���wF�W�*��0E�;g�Ȍ>�`8H�����gQ��I\�>u��=��k���d�|@n/H7��k��M�L>辡:^�q^z>�U�xd�Y3!ۼ)m\���ȧ�@���$AG�*�639�gz�J��?�L����;(W炨�����T�`Gv"���8��~�>l.8�E^��\���[��7�z�y^{l�*VM���Ê�+�J��4��[Zw!��#8��|&
T6�"�0i,�=ʻ�K��(-��;�۞����0�4zOx~%�E�^֧���;_/���5%bZ�/���sɑ�=J�.�����<r��3����/����n<�����C �xŢ�MD5�����q7��ȩ���Mp��5Nj#��1�AR�/�����_)�Ӭ�"W��Q���˥���L�f��"yi30���^�)m��;�gu�_���$nzk@m%��ܗX�O��nˈht�$�a�$��Q��Ӥx�薌i�!T�1Y�����=�3�v1�t��)Sٕ����ދ��t�����%d_�H��6Ҹd�;�\x!�H�U�]�Uq"rs�*�%�Y$֞&��8��I��]4��~��n%ʣC�^8���zȓ���L�2�*iM��7�m���Mr1~�C���>�p�ʤ̅�Z�Ԡ����e�5��]E2%�e�ϡn�Yz_=�W�02�ۼ�|�ڀQ�8'{��诤��[�c���/����烊T1�D�戓U�� ��^�u�Xv�K����S�t�u��@�������=\N��=���$��J�>i��>����++�N�+�G��ǲ{B���D�|�{�s�ZtC,��XA�ߨ��O��S"�`��	�=�[�GM���L�N.��Z0��d2b���p:��@&���Lr�@	����ڡ���L�в��b����8b,=އcdI	�,������L01Q�Y�Hb���;{�O�~wyћ�8��!Ӟ�J�z�"DH`� 9Bl2�a���E�tc�
�T#�P�(�;���*��<��GD^O��� �hbn%p�8�#HU�~g<Ai�����@\_����!
@k�*^aڊ񼎰.��oY!1�W"�F0ޣ"!ov��{fvXA�ĀMQ��i��}{�����^��j*p�"����A� 2����ew�g'����Y�[vb[���a@
�E� X��Hq8�2�|Z��e���l���=�&l>��<���X���l{�zt�� ��$-#WK��u�����=�z�B��k5X�Ώˡ�;���"�D�g�,a�u��o�țĭ�ṤD����4l�yy_�Z7I���H��L����@"����-�Ǖ�d>S%��IR������l��!�υ2�� ��_8���I��怡a�+���l��K�cیL%��QTX"K5�}n����oF�T��
�}o  ���+��ă����(�����X�j�����b�]L��TQ�ʢ�&L�0u�M� 2�B�0�R&����]��{,<*�,npYaG*|�G��@��K'���D���|R��4�2�^�x\Ӓ�H�(��KX�QJöBA�1�92"�����zhJ��A�I���f�~n��dbԴ�J�)Q���{fD/QT�4���Cn�%�Z?Ox����F�Y"h�_ezK�iOP��]E��a0b� �4�x�Шw�r̈Lha�5\*��,��L�w�/P@Ʊ�=69�ͤ��o_@�y�~�gA3��FҎ������u�9u��f1)��5<����c흳�q.E�w�D��Gv���S@��JY�?-F��R� �~a��/�-�8f��4�0qp�|���j.d�П3y�0e��uъ��#�h90��5��4�����uNj�	�C�X/��t������t����V��z��Eé�0��6��Ps-r�BJK:Nnf�9�*�U//�C�9L���l]�N�E�QQ�D����q��n�@M�x�JT#�x<�Qԫ���j�ȥ���c�+��:C1�K�����cK���.(��p�R*�X-)��M��ekz�L����te���@����5�BgpJ��$q�+����W�F�uEi����b��Mv�^��O�:t��+wį�(xo9���M��I��4'�������M���[����q�X��4 B-�X�f�GL�����Ŧ��B�?Y+��{m�K�Mj*]|b����|7[�dK�@t�&4�'\o������w6�I<q�Q��5�J�8%awq�r�1��Zq &T��g�y����E㧥�[����!A����c�{{"�T����D���q���F��.E\[��J���s��ŕj�P�کI��҄f�䩺�	ڔ��2x/e42�ٹА�����"-��b��d���[x��D1QV�;�hD���)J�e��y'�f,��c�W���9�����9�{�/J�Mrl�"a�h޳#7�c��=H��Iw�#�T����c�m�˚kڨ�OXD�v��1�,ڍ����D�2�G�J�چQz++��N3*��E m��t�`����az�|�\��p���TL���a�� �R,�^�Y'<��_)�3�����	��NR�ue��b7M	M��_"�3VL� y��}�}���[�������M�Hg�?��U���\�Z�ӽ689��0e#�O���v�@ɖ U@�!�q��߲PЧ��`o݄�@p�J��NP�� W�X�����{̃AN�����y���uK���� ��F8�D+�WX;r�U������unQ�D�a#�R�S�:�CTA�*沖ei��.�<� ai^�PP-��-�9�oJ�u�}�=��	.y��ъh�^�>���#�(�F�+2p�H6,Ǆ4#����଱���/R�3��TK�����ۜD$��h���	�nY�3=�".Ɍ�54v��.:�w�y�6�[b��$G��������Ք�!��;��C�26A�T�H�� *�(�$?�rIփ9���g�O1�Il��&�bq��U4�M�BI ����sͅ�!#E�yt��00@�/=����:�z:���x�4�E�Xgt+�?>)�����t1u5�{p���H���'Rpp�l�ͬo^ a��	V�7���;f�T������%Y'�0	(�=�]7����U̋��_�wY7�s�b�t$_��^+ ��X;��%iBbЏ�޻ތ��ѥK
e(am9��cQ��ҍ�*v��x˪�c�N1�X�)#_���ͨ5R���ǜ�z�MH�2�)|9Eg_K�)jM<�m�)K�i��}}�1瀒�����nm2��P��(��(��T�j6��1F/�bMG-���ޠu=9����Z8��"<�[��i��\D,�@��H�RHZTg$�sU�(��rp�aE�W��C���3�C����.�y*�|Q<�g���P��X��u8Il��t�>m��L��R����(� ިI��O,��"<����n7{�{S���k�i����u	���Hψ(�A:�g[o�%��!@H����� ��%�:��;pι>��h�{��su���-��Z�� �ڛ�[��̯ii�Nnv�I�;�<�h1��ל�
(�5����t��6��|�fd�O�;�x�@�|x��'�Ę�:9�/a*oDC0��H��F�#wL6�9�<.L}���D)\��拉62�Rs�Ro�J�{ໃb�m��e�},�;.�t�ڽ��^�C��5F��\ۏ�O��j^(j�۾K#���C��2����pd�#'����q
V��S��q���Q��9���M~P^�@D����i��3m�h�6�	8�&;��M�)�#'��ܙt�4��=��I%��%e�]& n�=CK����0���+R����o
3����>�g�v[��أ�:���轁��ҏ����G{�Qt�N�����@G<�:M��h���KE�� ��t��D(	�7�������i�^�JlsN�8"~�9� �U��os�K4�����(6s{�(���_�P�ˍ(c[P2`^��Z@ļS)�y�q4�P]l7�؝N��O�%[c�s�7� ��*.��D����Rz�VjD El.�5�}i�|�x�L!EGA�@��w灳�P=���|��%|Ki#�;���* �s����u�ܣ���Z*vyo>�0`��\_�v�
Q��T��wUČ���]/�$�O��ܭ��j���̥� t3le/���0�Yx��^�i��U�VK�\���\g���S5�?s;�V]�DQ���m�;^�5�D�S{˝�.�0���W�h���{��`
��^��p`�>|�m*v�	 cR������*�ou�B)�Oc�`r9���Ju�~��Ik�F ���U�u�TvMH�y��"j���\8��2=]�Nh��KL�6���� ����ч�p����tD����oL�3�s!��rQP���0�v�'F,kr*��� ���ۍ�e��~ۤ�jR{�@�]�	�XJ�x��_�f���9�&k;�0�w�x�U��k�N���!>|ڽ�6�Bl?�=3t7m>��DJ~��H�zX� �����������ȡNw�r��N��;����^�n��0����)`�� �����TVsS�s\5�e�[hv���Y�k��5����b� '�����+6aS�8pA��;ۨu��xOH;,���A|��b���k�2�A���3ACh�������vi.�R ��T,dpك�/�`��}��}k�������0;�^��i΢���oN_>&Oq�ON�0�ӴP���Qh��4@.�&�`��7~I�F���������3�̕��|��1 o�'[Uzar�$����>��o��`
�N�]�Y�6y��Ũ�Ĥ	1`�Ν!8��{��;�JC�g3���r���P܎���%�,���<����bk�� �	%�(��U�NX��Xe`�h4sWa���.Z��a;�Z����gړ�pG ���<,����З/=�'פ�]�����[���E]'���|�UiJ���Rߕq�%t6¦o���O�w;Q����\3zݷp�ຑ�~��yNM����-_Z���c�����YI�ۅ�-��>O��-�� �ַ�Y"�3�*��Y�G��2\�N��Ȇ��T���S�{�����Qְ;�"�K
ʊ�8�4��@��� �{�5J~�e��m���MO�6��qM�&;Z��k�!���ZPPTe��Y�BQ\~l�~Ky��8Ѕ�c��+I��226e�fCb�"��P��,C���%΍�8G�5�l�XB$A��
��A(��|L�BH���$+�7��bξ�#���ѡ�.�T@���W�)��-�U�O6�/��;>���~e �9z?��*?�nG�-G�^��8T�@\P*3[\P�^1���^3je��-:�����>HqZ :��u�,ub@?��9��_w��'r�D4�?�6�ZDQF��t`�5`~E/~/&��ɶM0�IX�Ԉ��=���M���b������:�	�w���8��-�C �Ӎ�y=<%�#����.��u_B��ި@Ĕ�e*G�i�KKl��:=�J�Nisl!!|���m��0.>����	,�ၬ�J���<��x�X���	�ARh;B�H�A%<���: �'6��3��(�|��Ch��2��B�j$�x�Qyњ�jfX���p#�u�v./�q�i�B7=j-AҌTj��㼴�_�x�.,ͣ�����r�=V+댯�Jz���F����<�σ��r�V���:�3�M��a:���a7�g�I��u�[#D�b*;���/
��A�l�Ѿ�{**�5�JXl��*xM8��^������Z*����F<����矽���`�������8/Ƙ�d�ZUy�" ��f� ��rJ7n6�������"�����7A�D�5-n
	��U
,�%�k����f��;��F����ޓ3G�-/�?k����)��9��i�]� �ն �~c7s�����<8�����6bv�7�i5�l-{���a��`?�2�")��ھ�+�x�4�~ӷ�S��H�T�c�L>���/�`�����/-������5�׺�����'h�	bm��Bb"տ6��]j�[|�P�a;�=�7����bQw��-��#l�(�}�	R*����ldqPB���yo� .�L�G0*(F�eƝ�6;���A���1��L�r�R�l���oc>���Qt�4��KR�V����0�#to�z4q���y_c���2�r��op����;��
Y7�U�������?��r�ƫ�$@�'������MqG���K�*��&O�N1�i^���O��y�)�5C9cu���� ܫs��a�1�"H�Iӱ�����T&��S���C�||����ݛ��je�UYwbId��F�عE�0m�����E(>����W�k�󺊼�������P���0�Ԃ�H�9�Z�[�c��ubQ��.3�&��#�]��-@����U�N�&�12�����g[l��"���-�Zu�q�Au��&���6h�8?�x���<�
)^�,|��\p��A�?xŃ�k'�q��N�딃�gg�WE�'&YLD�2����"��2Q�#�I�]��}�GO:^X0����N��(���i(���9�-�M<��1k�n(t/x9iP5?t�<Ʃ�T>���ߍ��
>���ls5/DH��@03mB�����/�t�?9)v�yC� Ϭ��2���$�1��@���%����>��W�[�9g��}؝����X�eH���=�DK�嬘j�b�cw����p�ْЉ+�=�É0A��Ò�0�{޺	n��]�<��M���/�pV񨧟���Ʉء�cVN����exg(",ұ_;��8áJj`���;�\41�zw_V{��׷c�[2ei>iLn��à�Gj�FU�z\����M)'�R3^MVS����\^6����㛱e���1N��Um$���q{�Hw\�`���� ��GmD�5C�nh*�\x�Iީ����$m�Gٜ��7߫��&c6��dVp��^,�s(��3��n��w��[�a�����n	<:G�@�b��G]9�}۝�/<z�*����M�}���k��o�u�=��� ��n+��-�m9�g��I#X%�������6�Y:��]�#�b�#��I�5�&;�O��}��A2k؎H��4��c�O�Eqc�����qXm���VX� X�#{����� !��F�D3�gى2 ���`��y�Vdg�B��?ÞHO�Ul��f3��ܡƩ��jK�[�	�\]\�:u�˕ܯ����]�?�i�W��U���j9�(k�PH%=���bO�Jv��D�7�� ���Gbs"<�(�Aķ�DDEgXwZe�����+�|T�SN[�D@�5a���L3)�X��3��Q \	�2}�XZه3�kN����j���#��L7����5Xa47{6g��qX@�:J�6nS����Q����	���%߅,L=~��r�C2�5���SVn�}\��RU!�ӔsN�l>6}�ڻ�Bl��0���_��j{���梲�n���h����sK�U�ΥI��2E��j"�9A���33b���@���� K��::���S��3���)�* �*�P���ů��0w1�}U�~$����Ǥ�+j�7{�B��U]��֡@�g�֕��[U���-��22�gV�#S�k/����)a:�G\Ҭ`��,/��M�,A��;/����Z&ahHŗi,��Qu�����2�6f��O�*�=3.E��}Q��.?�WV�Z��ԊcR�W�`�{�"=
v���'MW|��k�!�ֱpUH+�c�=�+r*��^�aE�)�kK�6@(�������Y|�ԠiBh�j\�I��$�ǳ��q>G��1F�Q�^��$Ε�Ńo��/�[��-�2��It��]ɨQj@����A�ʌ�P"��FS���nX��DgD����ۿ���<�\���B�x����t n0k�K���#ЯmBr�|�j��I��76��F�[&���]�����v�������%Д<:P8>��)\��/"�56�� (8�8^���Jz����������=5	1�ճ0��(���]��/QJ;���!���A?q! ����g�ns�Ƃa]T�ìf'��k��)P5�"�F_	O_��x�ω�A���]�W�Xjֻ� Z8ϣh��D�[�aljwq���
r�Œ���|`N��v+��p���/F�FDJ�����vd�/�Jȉ�/? ����^�iNR�&b��Ka�%^7�}�T$��Y�Y�5=�3T룂�ڨUa���W�k��z$��ZhWι�z��Ye	�2���(I�V�`0��ڢ�(�;(�с^��A�ւ���+3;�����\E����vX���t�	�}]m���/��h��1&<�E�7_�:0h��]̜���K'S���J(Y�,HV��=�O���Qz�Ug��&M�)�5!$O�ыˠ���;@�-�7��QC��S�g�ke���_? Yu��&_W��O��*��qT-�,~��۔'�S�_�~���܂�9��帤cbC>�Վje����N���ڵy��8ǖֻn�������7����~�jY8pJ���J�:�vK;<H�w@y^�K8s��ㇺ:^ͽw
̍�����0���g�+K�M#�@P��<����V�駰�#����Y!!���p%����=�u��!��w���Hx$��Eⵂ��*g�$јq��"��o�WR[�����	�λ��=�xLp��15��'��6x�t�e�_E�y�Y��I'0<��w��&�t��ƹ
�{�,��P?>>����ro3p۟k�a������?�Sz~�c�Ƞʘ����mg�+8F�����~Z��~X�s��S���O��l� [�D熡�Y�S6�t��c�v���/+#E��<L�l�$y�^�Z�AUgB|��vL�Ŷ���Z� ��{�w�P�ܽ	�L^M�I�m� �:X�C�I$̜;qս1kb��Ñ{��Ċ��4�+j���1Y~.�S!43"I(l;����a���ZG�R�R\i�Z
D��u�uA�z�8U4�)w\	~�A�oo3�z�|�J0�i�g�� ���;�Wf�{��M	:z�s��k#�+��˸�]��+��wAy!�v�����8�/�^l^/���
�u�*(찯��ϧ�*x-JbR��3��q^��>�)�{�����r�7=��2�-�pT�S��E��v�ܵƄJM�K� �%���f-j,��쯟wDmH9�
���+>F*�pq�����hlSr����C�PI^���e�@ɲL�s�Ğ1u�;s��Q����/�}����V�"<m¤ ��d����=��U�I�b�w�x��M�z�4�����w޵��,��ȸ���r�L��E[r1��p�0�@�N�~o^�O#{��z��V�����(��٩ߝ���q�n���&���2��8��G����@�y����:�H�fJHtw�P�H�~(u����*�~-�'�5�K�&�|��"�-�(^1�A��&@�}DJk��W[k�S�%Z)����[8�茋5Ůe��$�T>3D��=/��Td�P~��be�+S�*�Y_l��Q# 

���	�u����'��\y{a������rl+�{ȝ)_�@(��;8t�ի��w��|�7d�!-��+Ы'�,0�d�ھ�}/�k��3@n�������"Q*c��Y"�b
�$&l"���B2��lb�(���ѯ[Eߢ����~�6�?���P��C- с�י������6�ZP��!5��!�@Ӌ
KJ�zN�a��4��a��F��iö�^� ��Τ���Ǡ�I�(YrU}�-I�Wl�x�i�k�*�$�'�Cp��b�'F����bgk��u��RZ[�L����;��Mx��.����N%�u�=�J��i9vm�傅~����/�v'�0}_,�t��SM�M������EuI��[�8�<�EOn�j7��	�L�,�K��������Qlo@���7<e�$��n�ӓU@I��Z��i�߰���z�U}1�4UTY�_�D�b�����Q>81��w��W���A��q�i_�&�}[�E����6#E�e�P�(���c�_�8X(Ӟ�u� V�!�<!�xb��{i���q]�-C	=-[�U��"h�LM� U���=���J,���Nz<r}�|O�h�hӦ̳gs>	EY�i\]��"�-[�2NF�+L�?�����2��1��n�?��KU���u{Mp�q)��Y[[o腱Q�dc0������ҨK�i�	\0[x�������F������ #���;����GA+�p���M$�C��P���)�5���)l$!��3�ի��z�>�����";�L���!��bd��G�y-��c�q,vfw'��6F�D�D?Շj�C�?TY��v<�]�U��43��%�qy-J�%�c�^�|��s�[�P��D����3�6�fL��rl�@���~v��d�xV^��6�	���ث�5�*��6��/�R���6~�e�-(���Ga���U4�n�7SI-L��Bo�1��ɽ��$ܠk~y��6�ۏ�i���z�-:�S��hM=_�v��?GǗm`�6n�~�F䏛vY)�g�h�[��5B��
����GW��귮��0?�ާ>*s��G�'��%�#����]aq�(3�̐��t�R�����H��ֻ6�F����,���S�E('rG'BNHO� v��M����AF��T�?�p���&������3���9�sm��3�d`��B�Y������ e<��u�t�����@|^����纭"�V7R;RS�a�Ӡ��!���3�"\�A�F�CwQS��4�������#�,�T�:�t�:#�p�q��2������렯?��{g�u�x��1H_H�� �D�;쌽�WR��0��E�&��N��`#3N��q�U�3�.���9D}�p	G40�<���J�Ѱ��W+#�����L�,����u��6E��8�.4 }+�})�}�P�I˿t��'q�wY�d�'�V�U�(g�$�\��xmvs�&(J˷껾j &�Z�c��[U�]	B�C�Z.����� � s��/�/g�c�8_�E�����'ҡ�n��"v�����Z|�k�#P�W�(���lM����\bcUMpe������-�Uo�ư�Ӆ��j�5SaUL~�G�Q!gi�8!�p�Cblt>
��sT+�v�4��냚t�u����B�������iE'$���$�x��Ԥ���-��A�hAId,
dI��/�kq����V'a�BYt3��ϕ��ad�5�(���3��ݔ'^P͕L��3';�"�鎑;x;��]���II�ʲ��qOx<�����a�A�*��\�]i]�����ŋXl�Z1߽e���iҹ�"��h?���O��ȼ�1�D�%P��>z�2,��.E�9�s�V�i�h�/: (Q�h�w��4(Z����@��wp��r���ʟ0����]��_�W�+�`'�����F��`+�>�;����A@S&R�S���$j�؍�+��"=����e��G,yB��x�s���@�ػd� ��/�����:�㗏�3ʟz[Ҽ3OƎ����A٫v�p��n�@O�{nyWS�,���}��@R�q��oh�j�!�y�e�O$ b��˕n+v��G"�B ����./`n������!2�{��Cs$�wHL)�A��ܓ����N\�>���3�9��wd���z��jɧ��
���H����q!rP�� �\�wG J> e��i�Yd�gY"&Ft���|t��d�v��C�*�����㗴�ho�i�![]AZ�c�6(�"�·����4t)_��T�N��t}@��&�a���u��.+�w���V�0a���= \��}��cXb��x������U=^U�����S֏{�&]��s��K�j1�=zl|Џ��4��
zJ�o�܅�Y����x�f�Bs��m]�<2"��Z}�lb��˺@�)�}�;�06��?��7oy�[�g�Y�څ�
~>�bs ��5 ��Puy�nM��
[��ޘ'P��d�i�@��E������9d��+��_�o���f�;yr'��*J�OF��q��Ħ���3P���aPb�h2p��.�N�R�ꖐ�2�W:D��WAڵU���8��x����2y�S����?�����X�b|������5�����b�� �1�YM��,3
���]�r���u�{� K:�b�`5Tv2���3�ۇ�uan,A���QOjeã� '����Jx#����%��/���7����uw2+�K�35K�v���-� ��䶐�]팍�+���.��X���k}+���B� \�et��[��n�.�cT�Y�[
!|5d�x&��T��|ы�9�6��HR�4`� �.H6eh��"�9n��d�ck�OaR������~����5���D��1a��h$����ð�7L3>���M �Jb��0�	_ٍ!'�T{36��P^�ql��H�|��Mzy��?�P)�7�_�}iM��;�HE�O�B��"�!	��i�FPy{�8��3�TI�<��b,�s��2_��<R���_\ x�C=@8f�}I|	K�9��1H�/�)�I��S�{S�g_V鷍�a��
`t�XR����q�K[�Q��̋u����q����=;��r�&5��O��$H�G�"���y*��G�4�յ�@�I˄� ����2������zc��g)³$���!`(�X�z%[!���g�3*�kK�{�W1�R�B�qkȭy���zi�T�0p�H(�FP���ȹ��{t���I�/`뾫��'_Å(����pl?�/%��_m�"hY�v�� h�̡�g�����O����V��UB��ڤd�;��Ҝ����
Q��zv־��r�HĮ��\��OKP��uu@t�cw*;qUp#D޻��̺�v�2���+�
-�=�]�a�ɦ��Ԙ�!z��� #�T���nw~G�d.��Y����}���������]������>^�gx��x����&�99�o��0�8��0���L�Ӧ<k�*E�>MA�0��%�����Ȅ`o"L�4��{9���Ը�"Q���ǀї�.Sc�i�yC)fu/��r�I�G���[�Y\ӚJ4��Y[2=DB�=�2�X�)ubwZ�K㿕�:���s�e>�o75�񖓔:']W�&�~�"�C*����d+����R�d��� [�K�X�y.Ih֨s��YZ����)���>��h�dNNy�\���K�t��0,ql���	�}wcC��zPq��P0���%��uQiLw����c���AN\��\p��@9�-1���聙� ���M/��u��Z�k~Ks�Df�w`�m��^,�~ѓÓ�iv�)u�n���
-��b�ݶą��mC3	�'i��X���O�t�Q~��QyT���!T�� z�j�s�;�-["qa��X60f�|c�;X������ ��$�Ȧ�1����F�I&��x�Ck	\��{[1���'���N�C����w&����
�G�h��2B��mmL�۾��ʊ!ȏ�L�%m�QW�fn�'�N�y��\?g��Fp���KM|Q!�G`>tb�24"�_{9V|�a��q*)�8�X��h�r��AT�F�ƀ��Q�l�j})A/U']	�çP)��9k����Z�����*.OT��8�"�0zme��?��[�`�{��#A������Y�)O+/��+��G�_�W:�]�H��k���0H�ZǢ!I�c��a0�7?�Po����~�{��z��t��'�
~�=�
���v�S�|.K���,�'�L����P͹����s�M��Flfr��t�����K�e�|�;|q��m�J�[YΌ9l���X	��CW�-9s�m��d����"PF���&i/��u�q��bV ����af���϶ʷ��1I( w�5�)@�U�4���������B��v�y.Lc���c�v"�V0���'�;��ev$��ħH���M�׍�a�G=)�Ծ@��M#�酟�&k��4�te$�?ΚI���G��+��ڳI��
��VJ�NR���?,ª3?^4Ӥ���3��?�����~v��FJ\ ������B��[�B�)�5L�Ft)�a<u-��%����4��6�AG�5˱��e�a"�]�I��</DV�a�q�F�g��.�ݜ��`Z���x
�L�g�����^Z�j��QO�X2XH���i�(Q��`��ȭۭ��8�d�$A��)�����,%�T�׿xl���,ɯ�wF(;�*���Y�tFv�[���!B@p�{3*��zK�||��W��"�l[}=j��i� ���q�5�9K����}�:+����|Ne��%��Zӑ��~���`B�����a2�V,��MP���fPН��	�Fa��n�`L��0�h��|�§�#Z�
ݮ�����Lm��`����b]��f������O]^���F����(����H�ݑm:��D��Tnc�� �nR��w�$o$E��F"0��"���c�����X��o�d���S�(��'�H\���t�t��5�t�,6.�&�X9��=�kl�>�����ago�K�"3��]�U����`�+Fյ2��y�`�V��dU,����m����!�)x:{>�y.��1oY&�t%�zpx|�&�#���,������Iأo��lq��sK�.5��D��7�
st\X�d}�������7C��*6������e��h�����x���S�5��\���4�ϴU?g�r��OS�q�����89��ք-�Y	���.>�����C����$N�&�-Q# ��S���e������.9E|1�Z��i����!-sM��Ͱi�?}O��<]H�,l)���;ɂP��XI��^wX�f_؉��*�����l� /�k�#��p�@!��D
:��R&���.�����l�Cʅb֜�՜��9����@������6��FL�v�P�~�?~���a���ċ^]����.es5n/'����� ��=�������d��!?[�2��%)v:���#���nj��>�-��)��.�\{X�@ٰ����υ�}D݅��V�(��;�o��N�iR�gzE����~�Ɩ�tyf�8+�ue�렳�7���?�M,���4N�!|y��#��/JpJV���ql.�N���Je�{��(�B�[���r��w���V_�I����$My�XWMg���6A}��{pG���q	�P�ϗ��?z�F��o���
@5�L�u��b;ɗ~������i�`8I̢��Vn��O�aռ�${"1���l������ⴢF�UL\�l%,n���[J��C�-x��
?�sU�m�d��W�����ñ;�;N��R�ՙ�?=YZ(XZkg��6�M��a[��d��`���y��~�m/#S�D�I��4R5A3d!�z�)�(6�ι����ͪvsiCIe�w����H� �5�i-�����)WȺX���2���w��ҟbkzc��!Cq�����x;���q��
�\��!��d
���rq���RP��5I�J��U3�y�Fn��ٕ�`6��^�`чQ�ܿV�@�"3bϖ�S�H����f�_ƶD@���v]��i!G'V%�c�u/�@�f��h?�-���ѽi+�����K���������&���q~�S5�T>�%�CS�.PK�g������Z1j��}9��6@�I: ����V�n1>�W�/��KT�#j����*�`�i�s�e�� �Ox���?L��9���e��z�I��%�H�;|����ь���z 2���+�����&��+�I�����;�I�n��_F�^�H�x}�n�����k2�hƗq2���G§J��~`���HM:��KW6����Kf�v)�s����V�űSK�.� ��+}+-�kW���x��BAe��@�78$�5P�24-��CT�k�B x]�q�ԇ�K��R`��tק�Їb%��;r7��%�Z+�0SM��\-�g���/���O��&ܔ���p 3#�J}Wj�*��r.�^3����=��f@ś=ġ�-����*�ad)pSlK�K�m~��>����E���ˢVLP���%r^tΚ�g�L�uc)ϭ�/��)���a@��������73�J��XP����B%��D�� �V�\��dM$��W�/� /UU�Ҿ+%$�u�����6���n���]b��׋��1��2�FUU���ŕ�~�#�7+\L)[�w�Օ���u�EdAL$+�=
�{�Hlw�߫�m�|FJ�1hYHG*���f��%ƨ+�Bqǆq�����%�\iE�.;ܰ�@�^��=�g�#:Q
�m��>Ұ�-�����h�k��S`A��j=c`����$�;VqN��e�[z'[�KF��,"f�6�/�/��"���U��(�M�i\����{pPȴ�O��u6�9��0�E�n�'j�&��Ɉ~�jń<RM�vXTwi;C�gw�I=���e�b��� <�������}�����c)��jq�;d�pM���Qʍܿ����=�P<�����A��^K�p�N�cE�?q.��R�7� /_w�[D�3F$�{�m�,S�k�Lz�:�
\�,#�A�,Z5����-�������Z�'P-��g?n��y����]�Q|d=k��tNq�V������}�U��]�(�N�N�Ԣ,?�6�	�d��n�cw�E2�D4�k*:V�5G#�v�9����D�a��!)8@�sC}6������4ł�<c�����#�J=l�x���YG����v%we��e�T�Ld����UIq%�̼�O�F�^��%�9a����W����\�l	��V�Ȇ�ߘ����27���]uf�y ��m� G/�`K0�׏�'MvyI�Y�A"���.qn�X�@Ҵ���cb}�9���pf0���/���c
��F�!��y���F����p�&�D١� �P=~�`�4�9ni�u�� ����vn%W^�����h�;?�b�] ��ڋ�v˕����uf���V�ϐU��xa�t+����Oh��˂6[X��A��Y��%buu�p>�N�q-�fd[��S{��~�9�cY�{*_�Y!�G���Q�-*�v�Mu���-��ͽ�մ�I��g�m<�0`�J}�aR���% �_����a�?�B��'9U��ce�1*�|�7��1ѕ��4���u�ӈM葲����nP��J��6z)�{��~2/wS����d�Qa(��C"�K���A{t|��QO�� $YS�X05,3�����i0Cj;��q1�ي�F���4�:�����5T���nY���	[�-�+�s�L�W�F�0�Y���8��Q�|L�8Cy���l��}&�Kn�n�ѭ1��]�3i�ה*��?@�6j����(t�/~���@ �NU����xH �d�Z��}&AjY��|W��c�FB�}}����p\6�|U6,��ڠc���&x[�/ϑ禘��:{P#�|�[t���du&��Z83F�sp
���5��a�ZF��ٴGC��u�Tu,��qK�m$��	D@C_-���n��pWǜ	7�`5�Gݐ
�]k�o�>Z$��4K4���zT���.�oZ_8澽z�d-rz���R/oAj����T�[
��֓�x��g[�Z�uS2�m�ga�n[�x� 1a�\�Z,������$�;H�<i�$�����k��iƅ ]��__��$h�K酡���`�M�s�G�2��?�:R0@��kK?3ɩ���Xg���� RD������i�9Q"r32�r#�<������$�{���8��E�������M[ޘBl*��B�C�T��riSA�&�t��`�?���S-���� _���p5�j0��]D�ؐ���\����O�sS��j�o�f,��:F�=�E��U}�o� J*��[�5偃=�Kڎ����~�	���H�#X	L��<[�a���Dz��,��p�c('8���t�Io�������� y��~��(Ƀ�!0:uc���3�v���b*$ӎ�]���)�[�[O͆a0G�N�AN�<nZ����Xt�g���?1&�ˇ����"�|���E�;�N��B�u68S�0�3��$� qo�G��R�8�L�k�	�CN=����赕9�����Յ�QU|�M���V;�S�J�09�ǲ�z&>�>��Z253oo�h��`�p�=���z��7��j�,}����|Y�x��y��u�ŗ�x�����[A��n��.[����>����/��P#Ziw�0	��\V��I~�Qr�X�B��oE��V���b��<�������r��1ax��07__W֥a��h���9;�,���U�"?�.��t	s����h�R����E�B[V�D��GX�N,�]6�! dg�ji�Jy7�Ī����d@�R�wjK���b�4���o����;��l�D�45Sx��y�~R���Y��(����{�i#;JU����D��/l_���P!H��ۋV��6��P���ީ��+xL?>a��S��q�Xga���V�+o��v���Ǚ%�M�4�g��_\��m0ƛ+���]PEH.rY�
Ӕ��3W��&��/Nޖ�7\{T�t�筮i���ߴyc+�>2��=��!m�YWf�кx>I���%��_i
e���ʩS��1ib�]�{�%,[�X���v :0�ۥ�'�&�y]:ve/���3�ٲ�#��UD>[��wm�u���3P�X����)e�-���^�"X��>�MQ��h��p���<��u͢F��-~�u
��R��R"�]�׀ꍆ��m��7���$g+ ��|>3�7r',�t���: dE30Ytd΍�d6��k�yŝӔ�����Zf��/ٜo��qR��K���b�X��J7��!wë�5Rq��LA�[p(�4�rH!h?$,�C�"��ag�=%|xS�}�kD�1�L�8hm#��"���@_�f��\���C�X��-�2�s�p���z��W/���ٝ�m��Q�y�݅�e�7�/��jX Of�F�ڧ7A[�[�Ki�����,c�QR峝lW(���ؽ�Kܟrt(7�T=�a|�~��=W���.���U.��y�}��ҳ�N]�į('���Jx��?�5�K�!+6P�Aq���("�������q��������Z�Z8�J�BC�������Yt�(`���@�&�a�o�
|.4���u��2���Q.U6N�QG{���!	SHV��o�8�(�����֘���EW#���v7zʨ}%�]zvD�q��IO��w��mP�9~��,4��:K�$Wyo�fUi�������=��\M6v��X+��O>ѝ���NN���n���c���'�FI�t��J�.��D�p�a��\�`S�sw��7 ��D7���J=�אIs?_pQj�̣�4�q���E��ow#D��� ����K��8V�ۑG�[祆PN�\��7f�jkNW�� İ-EM'�D+Q+B�E�X� c�)��M��� ҽԮ���Τ<Mu4t-L<�=vk������0��v�+Q��L7�b�2dgˤC��됩�S�������	w�Y��׊N���NL�
�KЍ���%����⚨<��h�V%���C3�֪��*���h��Vy;߇kx0d�
͐�Q�.D~�]�j��~��lR��o6Cs����V-^o/���x9A�xO������껝.ً��uy7��A-?C�{��"#�9��Z�c�F����_y#�X�k:ONo�+�j��"gU� [>����z_#�N��vͥ'=�0�)�k]��#6cm�`���Uw٤{�&�F�WC����~�iBY�|�2�IC:��>�&n�	�_�C�L7�kY��X?Z�1Vh���d��i�@}N�o�[��贇�>/7"D�W\e�~�>��=l����]xʋ:������NI�0�r�GCO�)���J}qrO�HKΙs���5��O�dGxò�NZ?�E�~N�/F��|��%��!Jˈ�ic1�f��7!���	�O1ƤgZ����Юr��~�J3��$y�����O����:��q�� D��V��}�BȘ�S`Y��e�<�L��Y9ㄘeS��e��~�u���B��v�(�m�_�*R����ͪ��ߦ��y<uQ�H��v����eG��P���0����!^��~6���~�qlʖ�y�ÿ��M���'I�o�	Ph��|}=�.r+�e���t��:�48�C'�D$`:�CI5������D��cFUAG����_�x�b~�8T׸���������R��R-�ܑ�W���i��!���h�]s�o��F��dy�������:�X�f���歉!)�����f��5y�Χ�15(�='>y�i&���� ?E{�F�l�
����-��N��} ��C�I1/+Z���mG~���KM�~�Y�p��l��M�H-�
����1�b��p�~�t���?��z.� -=.��@��u0C�L{TY�y���l�?�Ji9YP��­Eqx�l�b�T�~ 0Z�G��E��ҫ�AN�զ�Ҿ�Ђ����j���|�M<���*��}�u9�*�n$7�f�憤���XT�|k7�%|����}<���z�r�+��m�ݻfE U�	����J�+Bˋ���n�}�`�Dۈ=�Cۜ��^|�D���W��l�z4�<p�t�`�ܻ2A�pLHI�o��@I%�B����
>?�B+G���U�+�i�xLA�l	��؛�@7��?��O�G�k�� i_�g�C$�d�놱_F��_�]L��g����t��Z#n���_��͒��B�J�A��`:5����"�����5��Z����k��ؖ)0a����=�</?n��O���A<�B��_q��VR��ɂѵ���Oh�`Y���c��.�Paw):�PyAφێ��\΢���Լk�,+��}���x�2Q~`�����JP�O��H#:j�%;+�E���;Z�o���ah�Qk�32��v�k��P���
<B�t%!s)����zO(hiዠ�Sgl6�������s*�kH�} ����E�m�=��=5�W��	y�6���'n�ys�7�9�6q3��Z]�����HB�Cw��rK��\6ٲ���^iD���/?�� ������O���0{�jiPt������S�q[�LGw��m3#��^[%�w����Η(�i�f�P/,!����0-����/v�%��h�yE,c������i>�@�O��g-��|~�� �7S,G��NZœ���WLޏ���ŋ�8gu�����U*��΢��Bc��{P�w8,��� pY��(��lձu(��]��m�gz��}e,Y����7D"P�UK�␃@0|)��U���j��*��w:o��od�gg��j�z/��78�S�g��A)� v�YC%��=�NMYS�<��������[��7:��^.��I�}>2��=@�����e
k���:�xf"Gާ�؈7!������ʲ| �.�����1�reIum�����Gf8Qhtcy���n�<���,��>wdT��
��9�����Wn�+k�� ��Z�[�����џ�Q7��S�=��c�m��1�$"=@\��8��E&�e��(�i,�e����>Z�#u�&�&N��x�Q�������C�?)J�C�	�J���|��w!V�?k@���R��8c����J�����>	Y��}͜�?�jᎿ+c�im_��@��uN]?9�B�Pi�u��}\G�}�n|Y7��*tr�ʞ ���J?�h�.�Z��;�{�������(�g?�����VUI�C���z�&�1�8�G�Yշ>�;��H��m��o��$iG�tQ��
�)=���$� �J7���.I��SR���Aob�FL2��%4�X�vS���ܳ`���
�#��:k��J/�:D�>i�QM\����Gz[���tqzo]M�4��\�4]������Z��	��:��y}߄�U��y��g��,�4�U���	�@���!нx��	��^M��� �=R��?7��M��RǍ}}%%5)j�����v��	�5�Q!��j�t�
m�Hq��O	lT�L R~�O^�r�&|P-;��� ��]"��}.��M��?�ڀ^'��{��~'T˷�c��e���at���R���@C�k��Ǧ�M�����4�qڮ
m��M���
R;�tѪ:���%���<r��0�`R�������{�9�A;�iPxH��fi�� ��<�G�?~�kv���?/�OlpM1<,:@��C�Ŕ������ G�u,n@ƿ����,�������#�}�WVB��iН_�
{
��*�/�쥤�7
'~�sl�|�ٞ$�07�/h�_�m�-�+��7��3���ׅ:'i�u傜E
�*�<~����[���"W��@*�}�-a�17�t��FY)]�P�@{/s���HFI��Y�!0a�:r?�z�e��������N�oz�q[R�o��1M�]�O������@N�	���͊�_[V��9'_�xx�,�?
�P��8����${����J�y�x�LF�D ��2+��\!s3��!��؞��t���r(���(�ZO'K����w����˅dh�Ɇw��`lD˽-颜��{I+	AdM��,N��T�
�g!�đO\�}��]�cڎ�Ǳ�fvp6?pG����+�1�0���w=�s��hD�[[��w%=�CD��s�!�W�����A�xb&O�� �XB� \6E
0��;_���T�%��bMHP�ޓ�����]g�����҅�S}�1�{Tg�$�6��2��d$�NK+9��Ƿ�h0�0N���5c����!��u �<�Nz���Pѳ&���Qjb`���7֢擆�x�i��S&!�.ˣ\�	޿���Wę��͐8B�6Z��R"��80���u�o�+x
�7�S�Y4�1w"�Q�f�3���{w%���0nC����� ٺ��^��oVt�Gb}��n#|ת�0�ީF�uD�J�E��^K���3)�9Qb���QZg���+��VU0�B�������·�"��F��LKw��K�dR�� ��/�+3��b�I��(��8����q��}�m+;�>�}s�X���Y��jR�^�J��c�����GGA&���_�e�F�e OTS49v�ذꔭ�y%�CTkh�N��b-��y�����:�k�e>� �9Q���_�ײ=�ӑۓ��g�bX�~�;� ~1+�x��$�\�I���Z��M��p�o��3)�hq�ocI ��Ù��1�mSV㧏g� -�����&-f�۝.]� ��D��08�[!\���3��0 �f(Fb�����?�(��y:�՝�m��f�|̿R�Ѩ��7nMך��s$$����=*>�e������]i��/C(�+��*�7L?��O�����1#.e�H��(�+،�^�\0��
��+qһD�-38���[�q�ꎨ׽���WX��62K Q+w��h�+v`7�#��"�^Ï��$�雁P}�_�	��/�=������X�4�2oI)jd�#�� s�Y�Jq����P�9�ԯ�x%��ɋ���,�}���|ސ���9~}}�`�S���|���9CH۷p|w�FgAS?�i
2����>b����-V��B�#Ϝ�s2 ם
�lA��p�(����¡�����5N���ܨ�>��i��ĢB��@��لC70�<��|���lq�2Y3�o��~�P�P��a�,��:�KU��ˠ�V��K9�%
�Q��V���i��E?�+���	(�ls� �l޷�������'��mI��� �T]op�$�%�uXKpʅ� }��_����sꏢ�ȎU�5cX�P<` ��L[���2�;ˡ㜩�>[�э��g�� "�m����3�?_*���d�&vIVY��ډ�*�9]S��"L_ã�0~�����L�!��ɰ�����_���G~�x_��ϗ��4͋*5w}�	;�F<�븄mT�A$jMK�����ź��2啂~�j���!ْKj��|_�"�_���.�+UC���)�{t��䆴~�i�W�zЛ�lK�����-�-/��\yT����x���
/��GE���g�a3:}8y	�-�s��T�%#�n��٨-a=�*�ۄ~��D8� $��Ǻ��\�����ps����S+�_�<p���pE]��N�&8xL�=�N �-�gf�s@Ɯ�mX�΢t>��w����f�i�ǂ���D$���1���"�TbL�/Yy Ni� ~�fq,%:U&�������5f�D7m�ʊ!��@{��Y�zOمӱ1	E�M1jć>�C���<�$wa2)$*x��������ޭ,�𚉼��%�`ܖ+!NX�A�Y34��f_QF��Y��$�k����سF�w<8p8c�����t�����ԙ����B�Y0�׷�B�Ծ����m��F1���&����t¥���7��٧��ü�,{��4T�=àE�V��-�\X<)u|]@f0v��z��`�T^����S^�o��+�|N=n���mC����St��}�r�ߵ�3aH���A���,�Oc��V�����7���KWHN�ؙ�Gԙi�`�)�Q��H���7��dHG�C�Ϊ.���/t��;��Л�*#�1�(G �Di�7�?��,~
s�\��� #�&Y6�R7���E��+vfb��ʌ����C�jqY\�(i[͋V����(���9Th�h��]�_? �ƀ�6�F��t��#4j�b��U5Zk��IQQ�9�����=�I|#�t�ܡ[���;�ٱ�k�c�ٞG��hr�l+2��to�P��)��7B��;=��Bt-� �kw���x�(7�a�Əك}��"��3��d%�b-��ʻ������r�6<�%Ǉ�)�R�|�ۉ��!��J9IJh����]�E��Z�Ib���,|�Z�7s����������P��k��KG��s�emA��6��[����n&Q5���4�u�P}� ��{)b��i%����f�nO�\b���G�>	�k�~H��)����B��@��'Hܠ��������C�ϛ�����Edl:�vo9�L�8��'���sB�Enq�(2�V����s'["�}c���~}a�3�޸����I���������3���d!ULd�\: Ƅ&��ʪU�r�$���"K)8�̡O#Z���	����M�
���5���H��椞_q��p�=���3V$�dL�H@dB{MEv�̛��7�� �j(� JОXFFs
���'E�K��q�C�t�F�y�I��NB^s^X��uh��	��y�6����F)��w�1��CD�z4��E�����ez���g�>�p�!���#/�X؞vb��g��@zM�ŷ�+Xk ����2ց�)�uZ�Ud��G;�2g��WG�0�+�yGz"�G��"��P����3��߯�efާCXlڂ{�V��
���W�d3͈-3
�S�Ʋݍ��Q���:���*n�٪B��������Y���`�g9\H��N�Q�(��P���Q�6��vC� g�:�J��D0I�v����9΍�h�:I�ډ	���9��c�l�J9��At���T=���Ͷ��/��*%	�W2��/���"i��	a�{@��@���%)Y&�[�d�\ac����M?�?M�qj6����݈/�^!tf팒\>3������/N5���?"�-KA�}�N%�4X����(ϼ`�!���a������~��M��z(�30��V��B8��O�Г��@�h�B��<��E[ ��H��)�vB먞b�� �
,L����&�$"��U�0 O)�u���w��H���A�]�X��-�<p����Pl��_g$��M|�}b��P�\�(t��!�)�S�ّ{TbcuI���K*�
B(E����m���%�a?]�n�i�,�T��s���W�͝l���9Í�J0��%�&���Y7i���W&l!}�XZ+z}��)�7��N��I�ض�}�m黣G~4Q��ʤ���5��Ncʹd�� �"�������<��Oz(!2�$�����i���J(���e�+���� �EMFK
A�*��s��bZZz2�)�ч����y�V���½�&_Q�3���/"���GDY��-�Q}��נ�;��)+ؙ�,ǚI��H�:��F�_��ޯ�����}��l�* ���`�e�,B��8?ꛩ�f�H�I�J�����b�nr���4z̟�]��f��^�ͷMPC��s4�ќ�.��AZ (]p~�Hk�:�� �P��ͽԁ���_j@�SX�Ϟ��3glأ�Y��������N8b�8Q:zE$���9?���x�j����5������,1 9�/���k�X`p�H��z�߈�eTRI�6���L[�����C��]1Sw���sab��8:��ӈ��Ј�X�~f���g�J����|�}�y-��a�DY\����	�a�<��������ZD�����Y�y���瓃H����@�����XO%�D�b@7���u�gog�����3�ԫ�9� �p�`���$G��>��x�-��)S9��= h$\F{�ս
4��� nL�^�t�[�������߇�<땪
}�?	��ʍ'㑺y����j�� P���*��"P��M�&RV4P��=��m�Tҍ뾠6V��g4VZk�,�f���j��$��<k�B��`�4_���F�ٔ��.���y^$���m��cK��)�$l,��v96߹���Y�����p���tk�X�-�=?��dM�4���'�߅Tj��ڔd�88"�}��9O�"�5��mtd쁔>�Vh��wbݜ��!b�����υ(I:�us� �L����7w�a"�RcoO����lF�Z(�֚����+Y�s�=���Φ~]�&)e@���#kڌB�r�(/�o�s��ݱ��b�Q�<��d��nSo�k�4�`��@K>F3>�#u���i�w��u�]pSq����H��0��e�4��x�}Gܶʃ��
�'�|�T���3���h�>�3F��C��*�����,7Q�`�-=&�R���������$z��i*� �u[�3���#�$��	Z�I��=��ȑl*����L�?�����/�E�JG��/_1@�F�����3>{��?Z�荃�d�z�2��
�(�Z�w��H��I�2=�5b�[֫�7��΢&Ͳ6&!�_�Ӛ���hI��K�R&��Qw��Wk.HA:+���L��,��y�R���ЊX���b��O�"����F��QT��R�}����L���&N�װ�:�!�4B��Y�+��=&�� �H9wL�������G�&����:�R,TA`�޵s�LL=��<s��ޠ~�}'F���_�%�����.�"�8��0�ɒ�� �JM�����T����l�U%8�(��t����+�oR�(���e>^Ʊ�|B�v�I6%
E�"��IL7Q	�RJ�S��X��|�4�t���IW[��Q8��g�~/��n�GZ�N�;{�zFn���B.�z��{���ۨw�,��������h>UT����[��Z����~�<�^Գ+��z�^q}���4w%DE�Բ�Ԇ>P 4C���ҙi��)�oK.�}����jO�̖8�����/��Z9�hi_.;8�c�u�������*R�C���m8�g�#Z���Wq�����H�,��b��h��ˠ����(�f�u����(L8�d�ю�ˀ(>D:��������O�z8��mHY���xZb�|�d�{�C�D(�E���f�r�f�JGֈ�\�!L?�a9������s�K�&Z(����q��s%����F�*C$�c6��#����j�ٌ/�T~~1��t$�g����1����q�rZF�1{6�U�Ţ�-8���w_N5
0�#�����~����<������X�()^�qw�|I*��Q���O�V����~z|O�)Pǭ�������ŁJ4u�<��%�t�@F�S�4�!��H⧤�1G��~N1��.f���fr��ڡS����|�^P��P��v�� W��_���>s7�65rv~��\2��82��Jո��u�#UeX���� M����K���ɇ�2����K��ec~�8���%_M=�U�
	�_i\8n	�kVQȊz����WQ�۪�=���h��Z��"����[YQ(�<x���z6A�dI�T;FԾ�c]�T�e���tL���ت޴�(�ոl��q,�:qcU~�s<�ak�'J��$�M��Z�b�t��1��M�c��0ǉ_��:�Ŧ路�5ۍ`#8�W�xqrN�4�?pv���Lo�<�*�e9�c���Dgᵵ>@�!�V�Y����Ĭ�@ <���S[��ɷ�x�7Jgo�-�9���Hgs��9�N#��y��Eb�L���@��yR|9O���<o�ę�'��u�l���A��x_J���l�n�}2������! �^����%�@�����/;�x7��56���EX@�"�n�h@��TE��1�0��[y����_�%]�]5%���d�[u[��Ts��Rfw�
.|��b�:~t��7�L�#Rd
����u�8����2Z|�="&���)�Vk��}iGq���� �=��-�;� 3���)���ԉ�V�-�w$�f�#���6�� S�G�m(��*�9|��+��fN'����3N��U@�뎙<��0k���a^/,���4�RSeF���d��ϴ�I8�E}�]{z�Ss�L��Ff芋W��j��i댿�ӧ���q:� 3�[������ح���=m`�%9�� � �ϚȚ���L���1����a��V��w��� З�'k23��Mr�L-yDW�f����uܔ{�����c�������G��2�����+� �I��3I(�9�4CFW0S�zd����-y�h�/DWިT� &^�^w����/an�'���	V�ẽ�z\��p�-Q���c������G#���� ��!�D���A�>�i�T1J����5�B��ѐ�DtU�"���Ŭ�+9.��ob�(*
yB='���$�2��'I���� �J9Ӑ�5.��dm���P(���ס
x���	DG}�������-#�զ�p��҆��"���T��X�c'W��.���!�齌t
��D�4�p1�8 �h�g����%�I����ʷXN�RL6��.�3�y���ո�Uck�s@H9�����t����a��3X-��:w�7�0�\��n�=[Y�ր����|n�)���O�c��J�aJ���#ِ�,��0tW�3�y4K���緼��l��uS���>0������_d�y��)/��r�ŭ��x�11��r�~2�X�2I�	P�n��GGZ�G�!�u��
�16Ҙ�M�E���B_�.N��H&�*��uaS� b����M��i7��cl,	Ҡ��e�>Y; }�rƏ��q�XhD�	�9��>��Ƨe�JV.F�2oxԃkgC:�h�_������ &���4D��R��{!PD�)q��)�z�?�Nd�T�I7d���7�Y�Eۥ#_�:s�5�V��M�==���I��8�/x���ʾ��<�|�',E��;E6�v���T�V5�r�����=�ܬp��I��M�L+��.��d��*e��p�t��_��@�
/�:�` 7�P��{�&e��fh�6+Ns�q"�"�#�VV�F���	?̧r��h�G�� ����+��v����/��Tŷ��S?F-���E*��)���?����{^L��ӿ��u�R�Ǩf�^��ir�U�de�"��0��ʞ��Q��bw�N>�{��	I�%� �4"�"��%0����H"w���^D�BE:��X�IJ�%<�\����:>G���7�����
nz(�E�_`�D��%��[p
���y
�ؐT�*���zP� �b���b�|��VH�@�1 �w��uU�Xȅ�JI0M�8�9��QZ�T�ֶ2d8u�g5�=-������7���|�2�䗗�ZG��J����2�k+�F4�
t,l=iᐙ��2"I��f��<���X�"�Y�SS�w��)'��'��G{[aFMGסe}�:�:�œ��:1�Gݔڌ��I"	��:Lѿ���Y�9�8�I�X�ϧh�k��]�h�����1�C�Hk��k�ohN}>���ȧ4�-����[1��V"V\_�Ǿ�_=�_�4La0�i�U*�A_F�^%�r�Ё�]�x!'�A��ķj����&gY�V�8VJ��>�f�uꕈCoفT���җ��K-�	j%����F��⦊.<���l��lбU7�m*CRL�4��Y��5+K�N�-����� �W�jߌ��(���zm7ˠP�[�p�_k���ɹaKOP��lʃ1Z�L��b�D>	��ZN2���vY�$���f��j��Q8�JH|�gl�����{�j8MӔ4�q��s�z!,��0�����`�2���h~`^�
�W�eh��Ş��s9�M�C����4��"� �*�%,�{�p�;���8,о,�D��Ѧ�Aܽ�ˆ�<Q&="�)z��.�jR�>"��sEJ�����gw1�wƱ�x>h��/�|	ռv������6��qw�^��gSSrW;�k%9μ��1�Y�������2{\Qd�#�S�����/sA���d��	��6v���Q��L�L��d�R*߂:r�U��I���K�1����3J������)�M���¤��!��V�k9����d��5��|�p3��4����g7_U�%��\����G���k�{R^�8�'p�ƥ��x�7 b񊾉�s��i�9G�����0�M������RD��G���?3�����,_�d�bט}��ʇ,�N�?��A���6�^��pp&A�J����e�P)�K��Y�0x���f�,gԼU���$�#�`f��]I�&�;��WD2�����򋤎���P����KK�m�4M��"e
�	��J�(	-r�Ɨps��aM�MyP��}ѹ�!��jTR�/�z(�-i��)|�4�kj�5�:�څu�9�j�~;�X\�������]�gOK��]�=a��h_�oR@�Δ�#k�)���Ī�������߼���U˯��~jw"� /����r�e�@�a��|-|�g���z��{��b���Y*^��Mؑ��=E��VB_@��;!|���q25�p*l$AfkR�:����e쬂'�E��c�XWa@^�'��� j�iz,f_&4�q�6Jh�[~%x�4���r��]J[�e��|?q�M*�|�<�Tc��8��9�Zܓ��&��`-kq3v��&rA�V�#�'J�Ќ̀�5�kc�c�;�ʣWm���0�r��#�i#�3G�u�_IS��͝�2�g_�'���7�5*��O8 ��:���a�\�<��@Tԝ[Zv>g�Y�D��~�bO�x/o�]o����_ŻeV�O��$�� ȯ�o�L�P�T�6b�i"㗽�ϳ�q�Q2&���zܰ�s�z�V��x�H�����J �([������B)�ߓ�-"��Gm����Ki?n����#'-�/R0�zr��T�� N)G�^*��lH�
#�?5J	�t�~.b>#!�x�3*fO�R�)c��j*���S#��p~ve�hT�<���ֆ��Ps=�d6bΔQ�;�J�w֍�#�
$�`�|@o��*������R�s��$�$FI���VtѸ��KM��R\�Z/��Iq��M:yLS�OMTJ��xJ8��1�!�� ���9��y��ζ
�Or$��-=�8~����\�p�W;-�G��~���ܟ��N�|�2Ѹ����_���4�z���-n*����<!Z�>?5/J@#*L��I'UX�{�����8�p���}��]���_��Q�'�܍�"��5�u����uW��4���+N�k�0>~Ϩ��hpS�*����jzKnw��eR�vy���0����v��;���B/N����B�7W4�̂V)���v�c��n�W��R֦L̴��1��h0zu���!p�Ԛ�<*�~���y �
��3p�_����{�CD�<Wر䵒�	`�8�IJ_�B��������"@�]�f�w���Ne_�)��&wA����딖��� �����v�2�8�&56�?���wk	��n� � ���}����o�w�յ��h�B�+���M��KS�v[	�8���/z�$�GD�wo�
_a]��ܸp���`��&YR�����o�g
�m�,]Ê�	��pf���}
�2Ͳ��!Z�V";1���xX�xHԌS�5�[w���m,�8쨚h�&xC�5mu�I9�,Fa�<9�Q�jg`��Lh/Q�j?��j�c��bL}c��r.�Hwl۷:(��d�l�h%ii;e�?�(x"i���(9%jK!�M�P(���<$-�Z�c0��h?���-	$�mΔ�dn]��S��k{i�bzU,��g�J���م�8_f8Qh}�uP5�d(]�&B ;B��֫v�����c%�}̇G���1�_J�����}퐓��M��5��s4��U7B�<�Ww�Fn|> ����uLv�5��B�.�{(��y�s�tQm�&��l���n��O���X��X�ƺPI2�Q�^[�U�:~����iW�96��t}<Z@�#:�Uz3h�N�l���<1�e��Jz�u��W�~G��:�W⚰��!�:ޑ\=#�
(�R�����4ךAX�����7�8���X2u��W���?C�ξ^5���G>�D֭����1J�\�dэB��7��>�ri\������3[���#`D��V�:̜H¼�Q�%��w!#P�r�(�d�b8sP�&��=�@?늢/T54�'G�I)�0�U�(�F�(���A��3�}~zDo�uMTv�t,+�}��` HjnRx��m�=ֵ�b HB�v*:׫���`���NӞ�=��ȴ-����{���1�7��pPD���8��*��������<�˪I~�DaQ�s�´��IqO<0*l���ʭp����� ���Ĩ��pdw-���L��4�I�U?ğ�w���]!��mz� �.��<�6�B�)��$��'�6�RS�H�['�W�tz[R���
7�W�p�i֞]�M�P�@:��y��z��=δ�����`b���M�L�dTȼ��i7=K{4Up;�۳$��D��'���H��.e�f��m�-�����>��z�����@�?�X��ĆrF}��ۇ����}{��4�3�Qu�%P�2��K>c��ӦB��O�_��l[�<Q��>����p2>�X����}��[���>jBvVA�
�{M^��ă���������t%���m7&�:�}t��%t��a�6��<��!�|�H�#@�)�ݗ������p(�E��Ä+;���QmL�����\�p��R�,�_#N�R�{E}�j'-�ե�(��"9�LG؎��Ӏ��4�H�M�^��C A�)t8���I!����&�n݉��M�=+���a�k�2�Z7�ٛ��j���}�CR�N�I�.Y�x�&��C0�qc-<�d�,۩�k�������WaOO��/����4�ŉݪ4rZ~�E�gA��ee�ȯ�6v^����C�k0cD��&v?�F9-�G^P��N �C���ڒ��K7#��o�k��a�:<�f�����N��9��KY01rj��B��%p�&��O�r��]]��	h�9!���v��`_Q��T�2[�ʯ�aTqi�v���s�Z qU�;��v�*ڍ~(���uQ[F��e{nu޽U���g�m#����WT�M��V�� ��F��G�D�8���qX[�%e@���V�w�@lCM���m���O��g�fD1��#���6��%.��㭟�v�V�f��l�'�je(���F�z�}PE)��x�]�y����L�	����u@#�y}`�|��I�nU���̢c��Y�S&3+:�9&�k��!\�*+J�+H_�7��u�RsJ�Z�[7�t���z;�HlPq2u��q�\©97�w�j�l��J�Cx����#�[�k6c1��n���֏l�[((oT�:���V9���S�Q��)��Jp���b�<��?6�WJ�|��ū��O_��T�Z��'�Iz;`m֛��"��Z�Z���^0OPb@��T�4�`�}��)K&�Ӣ�"=O��59�J�dm���J+I�ηAT'Xʦ�0�t�Z��t:0��~�m0�R<����(P毊����G�A�J�Ж��Ia���G�t~�e�
����L	d�|��r��o�4lNT�^���vx�{����g���	5)O�è�g4̜i�8[:�D���%v�-��e�O�ybze�"�UVxl�I9[���?�[\�'n���sj,4�4#���ٲqƖ�q��bLv��v
�ܧBw�^�b�ĺ0e��-|nc����`$l�����a[>��m���e2r����|=/�~p�@y�b�^�ψ���ߋ�<�I�iu�
�1r$��r㺞@��j|*֮�A���Tm`w�O����]���>�0���ݒCn��e��y7^�`�6>!���&��@�*%��y�0{x�g�t1�g�d{�}��d.R!=HJ1�K�"��|���>Z[�:ݶ>�ْ9"+Z��K)M��Wg�\�����(+�E����G@Id}yˑ��V[5b�x-����?�����H�90��g��U��dLM8+]ut@� ��-S���\��2y���]�g6�l�8ǝ� Q�'�r��	��#>��v	"�����zH���ELl�.�����Ϋ���M�S}�N{��՗��:�]�%���\3Z�0�jjn�ڗ�X�N��'QwT�A�� {f���p(X�|tѝ�y;�8e�#�K��fG�ذR����VP�c)֠��~^�⟆�KS�i{���[4�ɳ�.�1�`!�-݀7lp���?�,��?:��|�;��������$��	���$��3{sI([����r1x�}#�8��G����������4��Y��}��@Ż�,0��Oř��ur�+��L�*�,��	��2mY|�;��.��
�?#���a5�A���_x%n<�yAx��?p*ϑ0���o�E��&=�{�|�Y���^W�sULp�]n4=$�0Y��P�+ރ\CB*¦�m1A��pO�`GļL*
��'2t�&8������������Y���M�>�>O�4� �H�� b�̋���c�q�ǈ�n�����
�kߘ@���x�>1^�7}�3r_��}�����.L�{vB`�?>q���ov�<�m4���$��ؓK@�}w޸[O�Ǖ��<[�8_Z���U>)8v�����O�Q�ꃪ'޷u�f���v� nx���CW��u�C��MdB��Ⱦ��xTm��e��;V����.At|?l��׆�P��!g;��.<�#
�Y%1�`"�
��]m���r�~j�]�q�ӵ�T�6�14!��vf'w��S��tb,�0/�0#�6�ժHL6�Ö>���gy\�����M��?T�gM�Ea�E����7�hfQ2ĝ��X�/���w �����-������wbf�RB���!�{���9�C��M�z��,o3�`��IY��z��cπ�Kړ�r��VQ".9kT?�^���>�8T��S�@�I;r��ٗ���!�T�M=�{N]t	��6Z��J˅Ɔ�aj?���(�3�fQ��M*-�Γ���4 �D6�t@�0[C���L�:`#�N �67��S�B!(�IA.dM\��]�ȅ�����H<����r,�7fbY�%Ӈ'��ֹk�I��cCk��4��>��gj�2-�m ���L5��-���=a�Ęk�ɮi�'���h��]CSc�A���![��⒎�?�Tύ����.�ri�Y��B���S������X"Y��sA[y���s@_d
S���*͚���]����n~H^E��j�����9�h��%w��"�=�zS�s:0�z}�;��t�G�@��_��5�zpP�A����7 X��ؚ0���:=0�.�J_�b�x<�N�W��k��8��ػ���|�\�T�h�nN�����w�Ϧ�q�ޛ/�߁d.�yu�sg^�H"[�C�	�ח���7սG"m4T��Z?:v�{��o�,0	��X�PdI��t�,�F5sH�v�1���/���&E�X�t��HB(
�M���>�qǡ�] �&v���F)�hlY�&��m��)o`��ڵ)�����kv�cX3��rC��>y�6m�,˖�RKhG8^�5�|�N�D����(�'i� 
���QM�֛ZN���5>�H9A��~��H�\r���+{f��S^]�7����k�)�~�#U�{im.�/��z�)�T�pu�rₐ�c{�%���g������wI��B��2w��s��_'�T@?�JSZ��Z�Z�gO�)�9jk
�UVR�6����G�����g5�ya�D����ۊ��_�Ȁ�<b��I�c�=W�r�EJ��� �G�I�C����|2��5�AE�2�;ܢ*�|�}�����sT���Ure�i�̆�7��k���!��#��.O��%�ffw�L)�Z�g���<x �W��z��-��dR�ƶ�d�o溹��k�|�K�����ŌgE&�ފM��r����wV)�@��p!�b�=��{�CL�c6�P��sZ��M�q=�W�c�:J�~Dg]7��Щ޶G����E��&�5��w(}�<�9��:W�N���<.x��	�g��f$@�{!	��E�����%0]������j�?�M �N�M�A�j䋀�1�`�U{N��[Q��&�r/+^c�mJ:A3��l� S�)��Vg�#�'@�ݗ�q.��s,π� =��z`���m�=�Hy":�ǤX�'������8eN���&D*)�0��~s�s�aV�Z
�ޔ'Ե��}�3Ҝ����ǁ�t����^���֔�!��[ڍ� s�6tw�����Tm_6L)��5e	��P\R8�yYjXX�*����?�bcf6�{�Ϧ"�iU�՚2�Y����At���`(ڤk���PF^��I���Le���{�����J&��G1vS���|0Z�p�cKq�3�)��W'1�3)b��z���h���n���E6�m[y�v��I�pYɫ�3l���<b#p1��`��Twg��2����Ji(d�&����l�5 {����ʹ}{B�V �\���,�%�4��Dc�^*��˧tǼ�>���z�}}�P�oG��K{O�ard�t"��5DT�P�a����a]c��S\M������\+��CM�����a?�*�)����5���x�(昏��\|�)~Ǟ�9+Y�,��<�]|�����nz��NN����E������/+Y}��j�~�}sx2���S���`y�y�,JJp[�U�c#鋓Z`�g�L���Ջn��K!����)'�84���>θi:��2�������ܗ���P�8j.G�`x⧴HF�i! 'cw��B�c��R�"��D�k����?��+V5Q�֖�l ��9��Z�0z�[��	#N#��_|�u�υ�k$�4M���e������q#H�[�	���V�[Ѻ���~��z���x�dS<]�1�[�� +�������qǬr���_�Wx�6\�\�����@U~����n���k���$q���<����=`	V��YN��VQ�O�N�Gy��8c��	i�>���$h�UV�t2~��p���P`�)��\����
���e�TUԴ�.���8_eG�%��'\#�?��,a{v)Mi���#�����t�`H�-�S�1�ݠ�z-H�n�{5`��)>u-�\A:����H��G�׺������Ш)q�1�b7��G�, Vޡ�O(R�u��]���;���.W�QӌKoZ�Ӝ�$( �B���[���J��}^��q��B�Ѥ��DY���hD��s~&*l^�Z�qeb+ZA�(�k�Z�Lj0Rk�ߍ��\|o�%"��=��hI`(�#Q';���6���%�vM��z���{ׂ
J�촫�:�ҝ�!6��t�z�EL��XG�p:�~��>��l�<lv�R� q�1y�ڏkC�X�M�Jh���AX��R'�B&f/�ar+JPX�
���H����}P*�#�A(���N���/L�_(���5���w/s���-����k,�Y[�	٣�d�Y�U�k�,1�����˞��7�P��!q���G����+��jU�:�籟jZ��l'y3�QIP�aTb�]5��·�|�چ,֎@C��S��끇jǿ�L�i7کs��Ï֠Ο�E�, ��Z���]���YL#c�1�Ǆ-�CހH�[����ο'l��y���[1V�����O���k>���BT��j��������	�V��s��zC����4�T?'0h#AG���o�F���������R�A�Ӈ{�3�3/���7�zH+Cb߇���^�O����cT��%�OOh��)��B�h���iY¦c�݈D3�����3���Ǣ�哴o��4�4w/���m�g�c�x�8�s,�d0�(;1FH���c8�`1�A��:�*EG9q���9ӯ�*[y��kh�������`�'���.T�A�F��o�\A1�0�3�?"�6>��_�~��}%�������	�#_�d4=�!�b"�;����,�����pz�t�/�����C��k:�"{!n�/)���\J� 9p��M8���#�i
0���@��]J��#�{BdJ����ų9|�!29�1�2����v%��I����$����Çm�������4�[�7Uά�QCB����������p�Np	�&n��!��5 ��.����֙��U�:S�t�#qU8M�+�;ֽ#d͹�Κ�7zk~[2���"������˃e��%'"�a�wu�;_:�7fр������h;~û�V�d��4�q�y()/S��?s�o>`|�:��I.�N��/Fc�����!��1��vcD"^�D��q���;�SnT�NŦ�pU��j�xh+6�sZ^�Қ�i#E/�<����X|'X����@�pp,񥶾�2Q�(���'~�O��*��jw�$��i�CW[ı��_�蔟�	2$&F�ʗ]�h�������S��Ϋ3��y�7i�%0Y���vR'��SpҶ�ӥ�E�Owq��=�u�d�K��'� |������hM�c��[�kc�H��r�UA1KP2�Z9����J�pX_���r�k]��o��^+,ă�@́,��q(r�y�m=^[�U2�y���ï^���:�E*Ҁ�U.�f�Y(�;�
��� �l:�^�HP����R�D9����O�#��v���_�.�s=���Zn���̄77<t�
���F����s���C4*� ���@���_�N0�)���ò=����g���n�b�!h�2gh�_���!����"���m+��6��F��P����tg	��F��������g�E{��V�,�#��ES'�wMI�ɞ�h�r\��� �tu�R
\	Z��� hp�k�4��#��\���%Z�ra�1|��3m���[�F��Oრ�e�~N/��/3Yt0�'��A3i�CLYLļ��- �n+#Q\���+��@�p���zQ����&�q@LU
���F)�V�˰�5{�/��+�onEG2_*9l�_.Y�o6�~���4�"�W-a������
�\�S�#ک>�K��B�B�<
.+R�j�)&H�Z��dh���@��:�{�;��>��&Z�!q�a��x�r��D�x���MJ����fJ�P������R���܀��y�8αޮ<^�GεK��^ib��=��I��vu�`@S��?R�a�ry�L�pz�P�V��ß�Bf��v��<����+��m���Q�$Ct��9�H�s��" _l��ɓZ��j�L͉z�N3Z���=�/���*�>�-���"1;nX��S�N��U
�v��������]���93�%1���D�c���Cr��u��^�҃��N��ڔ0�^�����_�]k��r]�~W���ƨ���D��4\���g���:�X������� Xy�frI\k�c,))#��$Ew ����_�~�4فD�E4�R�`YD��Pج|4��h�������ެ�0��HE�NG��<D��Z�"}��Id�W��'�a�63�V���@��4�{=��$�f>����S��L��%Z�׆#������4��XT�=�QD�y��8���k.����R�uc{�|�#<�b�U��+ћ�O���$gW�	Qo���[T��?��/ż���q��m�?>^b�m8i�&T����Ƿ1��R�Y
f����׽rǻ������:{����za$qFx�B�^H�=��W���m/����K�k@�789���ď�J��8r�?�R5��	��y�A�R�.�YQ�d:�#��EH6�g�<�M���ˉPZ���R��8q#�KȝpQ��D��ֈ��y˞��<�#y4�`����6�|�����S���)T���N�[h�<�H��B�Mh�hxԈ�.�-g��74��?/�%��h�L�{÷�i\��e�-KoGsDv���X�Ml�t���'�i�C<FYt��I�+5�5 ����__�5�����o"�2�N����Zb}�C�5��EH0�}��mgV�%��#�>�'��<�N��j�IT�( �fK�*\�9߿:�<���&n��?�t�Lp��YQ_�dF�vN�;��lM$�D�d�,/�h�xM��T>�$��C��yJ15�n�)]��
�t	&��e~k<���_s��y�&�UL�^����R�6���Ǥ�=p�g<	"�Ba������9���8��ZEn
&�ك�$����A�*Oݪ�UoWH��r�����z9�x�8��vT�(����A���z|��6��H}�Y�Xn%�^���7��L>��8�؞̖ޅR?��GT�▓��{�۷K�SMAk(��;�������z�3�Vי�Ov����W\�-f��k��Xm��Sf�^�����قL�B>�����b�=��id�*h'=���_d|"���h��n�0X�p�)w�~�Fk���J�@D��7z"ai�i���q�%n�zb�Ͼz������8-�-���b��)\���s!/@ �@��Η�i|���n9/[�4k���$�|@�̬l����ժ�����R6V[����?ێU�P��8��`��x��?D����O8!G �Q��[{��-��;X��)�먶@�e�ԞRQ�BP1�vρ���[�4�j������^ō
1E����I�Twe8"�d|]�9\Ō��㺕;�Կ��$��J��,왲�Z�!Ȭ�}g�d��.<�j�,%Y�i]UtSjj�*�)'�E\fQ�H��=T�7�w�&����8�_�-�ET�c�m��ۈ� 5PW'[���V�M\^�������0��q��#-��/^4�2��|���ŮH,X�D��l9�iu��˭fiC�z:mM�PX��s�P#��7�[Y�m�~� ��[�^�e��0����CV�;��z��}-l��|g*y��Þ���.��إ�|�6!"#Ji���+z����!��[�eJ#�}�fc�����Dd�5彣z�/��R>w�Q���a��3������D�~l��;��+����}����\j_2���s=bs<�?L֠Jb�E�l���y^��r�.�@�I&,�[d��*�����uǙ�e���&�o*��
�9�n�ձ�*/�7 ���1eT����9��ߨ�˾t)�A���Qфw��
<.br�I$�x[o�]z�b��x1�9�&��YWk�:����f��F�!$y�+''铒�5��n_
E�q��,�D��=��ub�i���nsq�e�b&5�'�c����F��$�σ}WX<�k�[�C$��ʶ�em�lZ����@��0Q������ֺ�� �K*��bXQ�ʽOr�p�l;�,i�w�T�
�O�K��+��]����eD8*$�+��T���b`T��.J�|?��L3k����Aj�u=o�yD[&�?��
�OPr������`�LnD��|���'���
t����S̜�b/��J��
T1�wa�̯�c� ܳ���j� ��� ���~V �S���*��V�F*�10�((�?M��
B\:�w�2r�k9ia�E���t�����t4`�a�d���q��$���ij�سu����?��S��ԣu�p�>Hͦ8�45\�����qҖK�1�]Q'\z�i���Izy�Wq(��*y�)E��� %e��ԗ�����R���e��̋e�Ac�������N�WU 0�_���p��U4��^`�w�8>��� �8]=�ѓ�:h���%�.R���yЩU&�HW�_�ү}��b�fW
�������=����O u�DS_`6Dy�਽��m�I�[����g��G<v��)��}�д��5 ����^�A�ڞ�p�T�=}�
��9��̡3h8}ɥ��`�Q%]��U�u���n�O����j7�]�Y�op����$Yaq�ݍ����}ו��w0�[Rs\g�ZR>�{���{ᗟm_�2v�Fd1?/I
�<��9)�n�y�La��_�!~�N�ҫ�R)"�.�O�f]��������ܽ�r�?4�'��H;��#_�o̮tT~�c�p�	������ 8�!Se^����r{���b10��]7Y�i���ԽrU{����ֈ�����Ī��gy-��]敀<d� �e�@�j��������/�/B~Ң�w�o��ǵ�4U�h��+(����휘_Y���ý̓��]E�5)!Qe�~�(|��;v�<ͷ%"�*�ն{,�<�K�)oB*S�;2<����$�����\�!:��~E���u��w�^���ȡp��S�d�Yvs6�Ԏ��/��ƒzD��R籂�7;�\4�bk��>]2�*K�}��) )&Rn��NqND�Ƀ�c�GZq�A���!�ۅR)�QU�|�4M��r�Y�>T�Y�Z-=��ޥ:�)γ�JZg���93���g���1�%�)5zԡ=�r7�7ۃ�o[��0)�r��Q�p)���u����HKFj��R�U��־a���j��0|w�8����x�z��i�=m#�5*H��A7F�X����H�g�Q, /#MA��}��<����A �O
�S�*��m�mGWn���W���x?U�+�j7X<��x��]���8ڠ��^@�LЄr���֕�οRm;r4�~�4��J��?D ���r:�����@�Ƨ$+�*����L�[�!XI�����,R�d�5o��v=�"��i/'݀��Ӄ�͑���'�^jGk8�Ґ#�.l=e�g�Y�X��7A֌�!u�|}ȷV����`	����D����p~�ٺ
��9�R@��m.���G����[�'�dO��� d!���_�d�w[_�"�	ä��~�+NTU˖ ͦ��/�o8�U��,T%l5~?�ރ(N-�X��{�NR�ѕ5
�P ��0s{�<콍a-	"�xLH��ǸI3��Xev�tϟ8�� s\XUo:��va��
������E�o�����U4I�⢢����W*-�"��zA�ք[` �R�!Iu��R⽿�"W-a-��XK���"�#_lO#s~��Л���"i&��\��VǎTҡO�0�L��)>�d��@o�m���/w�z����m����0B����&h,�z}�$/�S�W�b]+=�?��6��#���?
�<hݠ�۞����;tw��F��KH�jR(��Y����TaZY�~��{Q���wh��#)��̷`���Z5"�RY:nݩ-b�I#���t���H�ѯ7�������ZV1�?z53��/]��܍[ط �#�������m@�SX>Yk.�u�6_���D�N�Ƕcܢ���f�Wia�Ӥv��8U)�fi9tIz##H���Lזf��9E�L�.��꒹^���|�H�Ų+���<ϯ�((��Wz�OD3:T�?y�G׌b�tRR�MvJG�u�5�J��<��ƯϺ�!���VJ-D�w��5m ���/�M]���9i��������b�=BR6y��]�tD�v(�z7t��9��yơ���b7RI�� ���WuW�: ���z�h�Wd�޴U�`�)�&��	��J	�5�� )�q�da� 6����L��}�t��_��LQ!���^6U�:C{�i7��d>��>�.$���Wi©g }�I�4���z6O�C����\��9,1Is����K���3�-F�~j-n����~B@oS0<�W��ml��=��:/����p�K�	\{�|cBq���xm�#~�P�R���7�ڽ��;�Z6�v?#.�wuOztL��,��u�,�>��Q'�)��w��@���w~Zw:,�ME7 �u�j�oN�۶�N#�!�i4B�T�6A�Q�_���:��{|�(H���bI��<Mㄺ|ڗ��1�$��o�OD}�G`��h�j"�qh|5�B����8���-�����
���B�wz�gS���H�X�n)��ho<�w�.�%A\�[�ss]Pg7����B��o�na����?Q����V�X?6f�Wu L�L9� ��~�4�h/��Ѫ޶?��^\����/�%>+L�3���62��|��F��!�_ ��ڤ��޲� ck���/D�[)~#zao�j2ݦC��Ag�Hn���Ha$��#L��O܂�(-E��0I�2���$X)a@�;ߥ�j|��P�5ؖ���>s�EMիe[J����*Kh�̐g��$��%�Rq���`�N�%Wv>������9Bod�}�F�F^��@� ���Fv��V'��M�O򨝮"=�
�(��)lb��|�:�$!��֣��$��&��2�ֹ���	��_SOк/ ���L�a���M��nC�ۻ�	���c�GJ4$���nQ�f�Boqez֐��m�1k�*�
]��VX����^H6�����5���r��lTG��M������� U0�}4/���Ruo�DW���L�p|��|�u�T^jn��5�5�3��v�T}ײ֐#�#C��KdQ-Ѯ����i�*n��_����`��?��u�N�]>�[�������I%��΍8>�H��5$q���A����x�m;z$����0�E1^d�EFQ Y!_���b�Fʪ4܄.Ѿ���c���¬�vF��9�4��1�=.C����%�3���3�z���~|�ų���mM����ˡ��7�(�|����$â�����g�	.O蒖�v�q�##�"�o�X��b��[J� ��M����8�Y�3����������~-���#���|F�Ԛ�K/�� ba�����&�/�<��Gq�jl�"1n��"R���(�`t�����"ug��=��ȡoi�:��'��g6��p��o�d��1_jL9��D:��`K���.�����z�[b��X��̷�CO���v|�@��G�gr/�Y1�M�9�rK�?ut`�Ֆ�e����5����s�&�����o6�����Q�Nm�s�oGuTy��OO��1�)K��焥�؆��RT���Ž}�^�W��m������9_v��W=ϵ�^X>�	�^��5"�{��nV=b%X��K_lb���r��<
'i�pMU����n��J%��0�2䭙���(�
hF1�>V��Y_O(*j�N��z;�ִoܕ?�)}T1T�3�n����_���0o{��VU�c�v��x�K}��V��4=�i �67S9��=Γ+�F���B��Vu>�M��g��_�kc� I��F�vI�YO��{���"+�Ш�f5�6�|�ǫ<�;��!h])�h�utm�{�iG��q��/<�L�и�u��`5D�0W�wm����;;���\R�4X�G����"���{�6���d�m�������cG��`�=�aRx�O�G{%�<�	�����9���k��<�0"�{j�t)���I�L��΋<\>���yN.L�ؼ<���)rMlf��Xv���r�0�S}p\�Ì�W,�{�&���7��"��oEQ��)��K�y��do���.�H�ua�Ԓ7�x�gQ ���KJ1��[�
b��������I<�i�#d�i�\}������f3��V-��i0˭�Hd �(�o�=6F:�ю�lPP�Hڔ��n�� ��gÐK�+���2D�&!�l�u�V�<��p�9�&)؆3Y�J~Ϗلޫ�%ֺ�#�V�l�X�pȐ�°�~��ݒ�i�%��%R�B��O��cK���ͬ��~õН�����'�V!D�Öˬg��h�����%��E	�ůu&��N�/S���:7�ӋH<l��Q�愁g�$��C�p	h�3���V�.�S���ɒbu�=�5՞��7�r��1���:�wv��	r�G2��Gi@fh����(��}sn�Y
5h�ol�ջ5�1xپ�g�J3e�tʠV�3d�r}X
 ������N9bm�r��4ž]�f���(p���*�zCeh�������N Z�.G��T�Zb((���Z�e��c�m��p�>�;L��o��1�m���i8sҡ��#��I�.����A�a��EBM���f�/s��"���65r�[����^��V8��,Ʒ�)NhJ��U���)VM_�|PƉA1��x,���.�zV��ZM�$�=:��;��`lz��c$��=sT�qޭ�:�`C�*Яa�o�w�.�b$�v�kut���6��Ckޡ��s���o�=��Zc�<���h���z�,Ә2/���ƈ���b�8�<��q%�·(���y�u�	4/,���)�����" Xҭ��6iZFm#GEʸ�8x�q9�Zlq%�"�i��S��WO�ӳB�e��-�
5��Y���9�e�����n/���/I���6����9��t��Y�I��ubm�ɍb�(y8���H6�~�������E���&ǃM�2�Y֣��j��<L-J��k!z(���;���r ��>˸Γ��l=Ѿ��򺪉���^e���m�i�=�u��z�8lP�;��`f-GOwy*6���}h������w
��w]�9�u�^�*|�,]a���J�e�.?�Lz-˲��Y
�\���ӂ�[��Yj]	���g�)�6#�'��OVÄM�QM��+�w�]��.+��Ǥ������׀�|�i9<J�2�p� �k��CY�E�xūɕ 	Y����K��H��Z�2	����Ne�� 9�}i�O���^�&7}@qE��i(뫷ul둥14=$3�� ���,t�֐���Ռ�>ԙqe����I�~"�N�H׾�nO��ݙ�����y+�p�9��HE���\#};�1��K�V����+����`D��j�I��	b���	�wGe��XW������@i��d� H�"��D(�m�J槶#z��i�Z>��aA��۳W6!�Il��k�|E��W�+;v�}��B�QM���#�nȬ��=T��L�L�'D�{j����ĝ픿�1����
i�G&�u���NSkX��B �ʸ��7��^�l�p�Kv]�@��Ɂ	��^�����cfq�"+�Gr[���������q�{�]S2���x�����X6v�׶�fZw�$�p���8��W�A��d~0�l<�R��l���J�r<����X��|�ٲ� �?}��� R�t!fl;�&|+�^�o\\`)��oY�;�7�гh�O(&n�:&h�u��m+�I!e� ��9T�>��I�^��F������Q�PJ�y�+,JJ�x�)��v�-��+����62u���h���A�09�{�1��+m�[9��#~��|8/����=LKK��Ma��{Kūv6.VI>��N�hD��T�����
#n��1�V�-GUP�l���k,� `����Q��%ӽӞ�.I𔉡��M�����ۖj�F˦��h)[y6a��8�y'c���=q�|�����,�l��������GE�X8�j�W��QXlr �\�����n�����R�Vk����5Q���W��#Z�{	y,2*ļփ�m~GQ5Xr����GZ#x�=wY��=����疛���W:�b�����"!�� �P�*f�hxە�V yyX�Dm�����u{�}���u(`�6�w�63Z0�����o�������P������^>����bJa�`�/��sS�]�e�kElz+O��Br�SDs�eU
��`�уT�ɓ���gH�_jk���9�1�����W�%ȡ�W�����X]#��	��H0��n�c��c�hz��Hxf<T��L��=���ldҭGDB.K����5R��Æ[�S�f/��9�	��˚Ԝ�\�����z�Yn��%�4aڑ���ӎ�xónD�{�k/��]D��޴�ʻ���1�(�G����������[�
�ƾU���h��*�c<�����Q�F�3|fʖ6���1h�[eo�Y����0�����)�e��:�f����b�h�ې��~U�.�yX+�������Z��UZ���g�0R�Ç�zh�G")t2a����;Pp:�b������L��a���&���]L�P�6q�QATLKoo@I�#
�8�Й֎�n#n�_�X/�@��j��<ƳZ�p�tG[B X��z%4�p(�n�%�UEX�F��Ѕ�8&��u�@<,y�*�iH��[Þ��&���Jn��(��~����֝Z����Ofֳ����A�$����&���
Ϥ�ֱ��iy�B�
cF�d$xUK�n�Ne	��.w(�S��x�T��}���~�Ox^�,�>dO�4��d�dZ�%���Q��2��Ը���j���f�pl>S��o�G� �#r�2����/(YMO�D���W��I�h
ݼ���^�D�������1�>�I���1��]����K�4ԥh�M��5����3��D5�8���ݩ��ֿ����d�
#���y�v�t�C�� ���[���a�)�W���Y{5}�=��������JG"�����G �g{&�Җ7�K����p?���G<������&u���؃3l�"�mB1�3f��Z�4L��,�W�*��MG2�4��`[�2�!C�_���+�ú�����\T�e��� �.�6���?T��	�pz<���VI�.!�����% ,`=�`vIt p��2��6
#�����e|#�[��:Qn����к�M��oA�v2w(�W�E�Xړi�ZPJ���b3r�Z(|��m����s�'�-^j������Z�k���UD�fp��ڣ�����e2ob�qC_+�5�T!���v���Ua�g�������1����@�ku��\M��1O^���<����d��� u%��%Й�)zv-XJ&IQ�;fY]%v���������vM6הΒ��
�r�]�����%�f�^�ͫ�"7�9��rɶ[�# �G9w|���Q��Q{�'�z<��o@{Sdb�3��'�=+C~C� �z���^݂>���).kL��%�	������V̛�Ҟ��?)�gV�Z1�Чq!��Mק��=�n������%ÖD<�m���·"��ͼ���<j�*�� �Yi%?��)��w�v"&ƫ��e��O�9��R����bk��x/��Jf͸�����	;2�;�Cş_u�}K ��a�o�S�����;�|�r���*G�9k�O�~���o���c�:uh�@	T�]�&f���D�A����6�2��sI}܎�P��Zc>��z0"��c�)#�)��T��ߪ��+��g8��}ԟ�=�v���²�֝LY�za&���l-�A��?2����7�����^���irn�o�y�xKiT(�wl@�ʯ�S�n����v[�9�6�hZpi��O	�1�g1�Y��zx榞�y�L�;~�s�S���M:�F^v-�3���N����K+@8|[�����k`�Z�9W|î&�*�ZB�K]	k)ؿF���[n����Q�T��p>�n!�����;<�V�0}{r-�~��#��ӈ~�E]sY����>s�V���@b�����,�>Gֿ�sx~/�[�'y�7��y���2���ڜbѪ$@<��s	(��XZ�(���ԭ ����^Ȩ^	4����� ��!�����r��B�b���g�л�o��e6x���c	<C%69ɭ,s}�<��_�X�yo�T6��F�hS��6��K
��-��d��RH��\�?d�WXRz�3�g��Q¤����b�+�n����Q�U#�����g���(�1qA�פ �$'F@J��B�*�6��%g���`�FݹGL�TW��Q����e���=�,y�{Tf:3+�ڷ�ʹB��Ӊ����Ƃ�Z�#D�����	����ٛ�rHIꭞծ��J�g��*�?ʌ6�v�k?��8ےă��-{�#{�`p֡ł�c��6V�@m�jGV�j�Z6���%w�9�,�^�	�ж�鞶h�����N�i����(��Q��֔�@?���P�D3Gy��=5��\k�u�E���Wu�D��ݙ�]����/Td�(����@�S�#8mc�C�$ݕ�z�&�Q���/���C�H{Q@s�ξ����t삜S48�?�^0s�qse�R�Vy�T�	Zg�A��Ѥmj 8dDoc�r�w%� ���[�r��)�Ӝ�t�:JMN�[1���.�6gz�'���FNƯ���*��R�Ѡv"%�Qz��vKr������zH��l��&���r88Bi��`#�F���@�n��J3qTu�-��\�#` ���]��KS%K�����*;��w���I����Jp�H��ӊ��Q���� %�(��Jr��5g�C6���'m~P���$�I��	r�����{?Lb���ҾIP��[Q �#�%*���>BQV�aXH���R�7ض�����wq}8�)�M�+i���f��]l9����34���H�A^�`I�>���C+׿mb۾h(��5�M|,����貧����ӸWV�������212b{Q��˟����:#0zS[����|�ÞT��������W����x����D��ӟ�J�?$��Nw?���9JƬ��pReթm'/\���I�5�QD��,̜n�����e�~��"�J�%�+��4Q)|?�<d9��C�ɨ2��������b��	�xwB��cZɂA(�����Jù�0� �a�Н�q��C,�%�܊�\��;���h���ʑ���?dH����E��;|���rt%�[�nE�`�A썹��(cꅢ���z�o�0^� *-�n��j���X�h�;�K��<^f���(a�C��\#a�[h�
�@S1��Bz��!�_Vj3�A6��v�X-�zڞ^;�VC�d�p���i'C��6����"�Z0��o���c�E*��s|ϟ�|�;�#�:��K��´���9��F���/DS�3����r
�v�O���ԧ� I�J`�@�]����w+��J�R��X����G>��@zR�5�I$���X�/`��wP�����w�� R�£��.
X_���M��[*�0�+uft�ɮ|Ԇ�\��U7¼3���/�����WlVl��&��(���Hr_.��<4�ĕCO���e�P���Q��-ZɌfuI7�߽�#�@�F��; ՇHG#6ՙb&�E�Ty�A�*sR���Y5�9�й�ޕ=g�hNەt�I�R�xn�$UR�a�t��E��1��ߜ_7� ��/���u�C��Ĭ��ˬ�h�6���[��ڧ%�w߄���jv�kr4�0f�g��q�!��/|7W"z�+?�?zTˌP� ��,�^�r����	^θ ��H}N�e�d���mɽF���#CL���󳰌��
S8�99@A瘽#�+K��k��Uy�!�n8��`��Qaq�X�����s��_i��[eξ�:k�U�UYKg��B�_�3�ZZJ���/X[����z�"L�3���&`� $74K��Na��o��侰9D14�)�VY��L �6ݍ���ˉ*�|������M�`�Y��)׿�ȏ;���@��o�A�L��gd���xO񀍀�5��� ��q	�}��(L��~�LGx:w��/����h�Ë������WX�g���:��Q� �@*��ݬ�B	��0��%��?�[s�'�i�DϘ�m�c�E)��xEd�ܭ���M�� 3�� ����z�ڡ�-I�}��_��[�?=x���N�s�\���l훋`N��D���^��١%"[�B�h�A�9����̲��P��-&<DFՎf>���rP�S��ѓ"F��R�J6�b��W^��X�����#�h����b�t�µ�u��e��fh�T5��"X�@m��@Hw�T����59[r�&z�vL���d�YM����Z�����<�/Z�;� <���P�\A � �o�.�0�IG�F�%�_�CB^����\<ۇ~\������,�n'9���&u��w��ފͳ^�M�{�h$��k��a���4m�ZX
���v�eZM��%:h���>۲o��w#� ������6��9��2bĽ��4��oꦐ�ѡ�(�4vɡr��j�{94u�XN]%|Y<X�Z@���>S��u1�uґ�Q`�u��W7�,o�!��a4+��BR�wc��f��	X��5o<#��E�>��kљ�p��}F�PfEg^���Ы�rv�ȵ��ٶ��s�J��v�mH\��vl���>#\��Ay��^`t;�����_{�,�c���ښ�W=�^�Q}Bxl_��'%��_!Ы�銱�T2I��!<O�Zq��a���:�?J�a��^m$��:5�`R'aw��
��EЎ���������{I√&x�lr'��q�x�`���������P6�8^кF"�5�DحuPoL):&���K	��R���J���D�	/�>����:�tP����~��0��������@���k
H|:/mHd��L�>�橑�?��6ŏ'�����9�.(�� 5�7��� @5��S�ᔃt�C�3�UwZ�ג��s�g���;ѝ��!���u%u��^P�wp��C)�����i�d�("-�忇pn'��^kL��hq�<V�$!o����|�#�~��Rl�D��FFX�\Qp���k�%�#��5\��dMl����@��^���c@a�J�� ��.P��5`���~^��C�n3�'����yW��cC{��1��Ֆ�K36R. �δ�T�[���#]�/�c���P鯳�Z�A�����Knm����8�|{͍w�����_k���c}a��8���o�6hf-�ԽP��K��-�c��T^��v67 ;��g�3�Z��,u��7UF��p?S,�N�H��Ⱥ�L
Q78H�kI�
����P�4'�=Ҙfw`5{���߲��_r���]a���̤��n�v�<�-n�܁��y���5��|p68�^��-(�2��~���b]���X�A��xt��>t>("�e+���7$�ޜ��|�|��iGS��{�G����pkΩ����Y϶�/�
�q��������L�!���dʎȭS�̳A0��[E�#V���U 9>���_T�I��;,�aX,��e�t|�$��@�8\��Ƣ���n��o�ާ�!�6��P+���JnOyc��*�O���T.��\Om��Fn��RX2/o[ұH�^:B����A�	Ň0��FM��j4	wh�.	F<.y{�ɳ��7j�r�����S�����/ug*)�Ԛ1�K�U'/��K.��8�����Xv���$B:p��;�g�c��T��k�������\��詙�1y�֏�{:r1��� �Vm���!7=S����I���?��zԊ��w���FT;�w��{�R�ꔹ�;b�bbcv� �~��YNΡs�����7a�V������rMY�����zU�C�g/6��kZf�3Y�]%L�U死�e�/�Q��s���>u�ࡼ�]����ӕ�P�>��������`�83�HY�'F� ��G��{ �!��U-7������đD_�����T���m�)%[Eƙ��k�v��vƫ7'CtI3� ~�O��RG����X�Ғ��bbN�M���$�%���c���$g:��B��$�8҅9\�����f�l���*F%Eƙ.�)�р1����Ir���VKN����޼�I^(Y�d|�_#w
��d����M�9��raפM���bVD��p�qs�p�PyS�!��:N�R���� ����@��x��4�<��Z��u/�+�:0�V�����b5V6IQq���y��@�fh�1��S Ʃ�H/�fSh�����D����H�.W�����_�r�H0�z!�ir��PT�G�k�8��[����NWx!=Zk��6!��-�R�֘���9�Ӛd	֍?���|0v���Xn'<�X�Zܧ �P�m>%n���.���T�0���^t���[aRߨ�Ed�F��WGOxe����L��p�,<I�`�^���1JȲ�z��@��2��h|��L\�M��Z��n�De� ���-D��A_;�6~W���x��@�՞��Y���E�2����p3���"��o�\?��E"�TN�Y�ę�0?7����ȺE����e��b��!��ǵ���Ib���Q�!||;�Bv;�.�O�s�KY��د�:�m�l����h���=w�x\[	u�{٠�^�-������)w�
�/l~��B��*��j�y�MjE�z��a�'�R���6D'.d��i���u���X}
i=��IM��p���y��H'�A@w��m�;,R8a�O���9������ֆ��|����՞����Zmi:��ܣ13Lu����8Q:p�k �F��qE<�m���W{g�`j9@W� M�z�5:H�c\)6����թ����z�03��ڮ�d�mA��='�`;�e~���_�o}�M[&G*y��B!�R�~V�S�{�uL�u�ԝb�qd�g��0����n��t9<�/1���H�7^-���	��x��%�6I���~�kuށz�����d�{�5�'�|TE�}�h�Y�t`���+pj�R��C�xG5ג��,�m>!`7;�mɽ O��V܄�����܈ψwqۺ���#i� ��d�;��(ut�9T)ǻK�Heh��o���D>���CY+�餏_P�lWA�Kd�+�(0�t���+A�q�#��T	5bcc�h���@!7��%l��4���J�*eB�w"?av���_5\��+�ux�����L7�7s��e���~���H���a����=��(��.V$�}�!�9Mh��×�l{��AB·2Zӥ7�;����T�~�5����9t^}x:\9n ���Yě��OUo��R|�>�S�Z�/�`m�8��4��,y���.Z�����J�['s�]�\?�X�d7��kȬKt��mq.G�3v���&)M�I�p��^:���y9���z4�Ԯw�b���Kl��ܘ����
�չ�	�n�'[V���P'�z�:�B��?��Q,�d�?
���!����<n�f@��ƭ�������A��\.���8���������c�E�!�R|ć_�:�ų����laX���w��&���X�^�Db`��M����q'�h��zGͪ�u��9+���t^b��a�D�E��XxL���w�rN{�)X�6�f�Vm
�]�%���������������NX>�L��R�[I2�� �@���D�:�"R�¾���0�p�g-���gbJ1�!?���=�i������)R��a�5]tiԘ�9��s�%�����O�k?ێO�ȮC�%������,5Y)��gMb�}�2�7��� Wpf�J6�Ș`���'Xo�W痌����r���2�?z,G��)$Q�l�>1đ�BK��m ���ڱ�;CԘ*#
C�B3�b���������<+���va��H%}N�=�)V�L��i��D���?;"-�oY^*�m��:�~~ݼߎ�\�n�ݨƹ!:��4��e��c^8p/�����-�o.���Zf�5�$��܈�Y;�G/����7J#�L'�$Փ1��RT��G�<IKu�����K�P8Q�֑��դ��f�\J�:��L�*­(��È�0$d3mQ��_ZQ2�'
7�ӿm��<�{RW��g��ӎ��ĕP�']\�/�Qd���(�1�~��K�rkB􈨁�7 � ����X�S��U��[�C58���A�v�]�db?:��ɦ|G"���VŊ���w�j�3�*�����3���3���-�j��,�hםL����A�q���b���/��f`�,�/��2A}xs���čV
��ω��|.nƔHE/�5p+���W�����_��讶�2����_?4�L��T�Aw@���X�7�j�ɦ��N内��uez7r+���fۆ��ۓGm��*dZ��呹��Y
+�C;B�W{��Go��*�(�ʤuZ�(3�a#����I����'���IZ����\���I�7ȫ�ͽ�02�徯Đy#{���%y�	��H���$+چz��D���"�n���ڿ��ye�&A�1]�������rm���y�siG ��W����hj_]���E��p��ȝ���`P�^)݀�%�#
�an�pp�6q�t_EIn�g��ÉE'5�5}�s0,JA��ާ^��&T�ȸ�I)��R���C���|3v�qM8H�\�������	��p�J7,?+��*��# <c�#PUFa7(	�lx�������W",ľ�89��nƏ��)�����)�\�a	�t�ۄ�[�@v�ox�la�WA�m�%��\A�67�ex$�7yD�%�.��C"�L�-���L�������C���@֗t55A�hE������o�Q?�J�:�`]>Z�U�I�'��5~q[��=k��<�0U3�?q�zӽ3��Ռ��ں�H����3����16*�0q�K�ɎJ��x���Fv�}�N�l�G)@DW�F����z��V~ߓ|T
g���je�6�������A �2�@.��'oۄ7I�|v�U�U��DHG-e0f�=Vi�;K
@�8A���o�+#����b*be�6�7=U�_�a$��X¤	�>���?�^g���ӯ"�a�C��u�E��aMTX΅�'�?�k4��H���|�0͋@�:�R͜�U̓[ViM�Z�V��f~��3$�01���x���S�����B���t	m�:���GA�@쳎/CWC�6�Ăρ*٢[1�G�g_�xe�r�[@s�l�Ĕ&x"�w��0��k\ۙ>�Y��!vYB�8��� 2�\-0��x,�����n	��J6�κ�%/(�oU	�����?
)�WV@��. �{1	C�Y겯�����|�������Ҧ)��(���+���,�����s(�����| �*�Ǭ������Q�O�W��U�3���xUҽ�3�%�\1��)TZ���bP]�թs:;�`���b75ЕO�����+������J��`aΐ(5|�Dem5���q~�:FbGÇ�|�{�������U��~�@��M��M�T�c�
t:�K �\۹&�C���a�2�a��������vOVA������`�26�lN�ɷd�}�J��\8$����X�)��7����́\���y���jW?O��!O�D-E'xp:���b���g\{��o��-���	����={�9�����)����O��4|5�-�ٞ�n,q����xn���q�'sd-`�yYc�'�	��Wʮ�l���~�ک/�e�����x�$Ӱ�a�P�7���8;�����|��T�B����M���א&!w*�]�$C� �.�2��,]����
���%DL0��k�<zihA}�e�qL�q.{!��RYi��RFH��������xA�u%�d�t8	� ����=, ?�ي0��c�2?�@x.��35���s�Ϲ�hc^-Dd�;J�G��X~�:�GM.�o���-�p��L���|fs�����"�7����I�~;M��J׆@Ց�Z��7q����d�d9�}���>Z�����ˠ|8�ʅ�����W)�`@B���b��ɒ����M�k�&�OEw��S>� ^��/�OZ�Mz���l\4KI��:��Ċ]x~��lƢ�s�����;6���cz�񸓚�0���d!���:ݪ�� !��w��k��]n9=	'����fg�EIc
����Rs���������,"`L��@���[Wb��ޱ�6�i��t�*��Kz������4g#.��@fI���S�O�}烈�"�X��Q��Ѥ�*���b���5P��M����S`~�,XltCϡc%Q���E��'K�<Tj%p�ך��Lÿ�?i<>�>	�Y	�)��ؓ�!�Jy���D� ��b	��4d@�z_��C�w����FS"�nm:q^m�q��M��Z-�v3�"��<�פ�VE��k�0ܻg�²��d]�Ն��-�s�C��y8(��z�nm���8��|�NF�L:��R]�k1�n��<���㣮l�M�p�	`Ȧ�ge73�����ʿʓ�9e���<ֵ�E�@!��LN��5����.�W�w��m��	��](Y��
��:z���ɯ�Bt�0�%"�Jz��*d�M�]ݪu�)�Vt5��!�z}i�E�r��.� WF�� ��F��ʾ��@��>飅R�#�Q�@�q쟀��G�(Nn���L�fJ�1��L�p��)i��Ny�w��|y`U_[��@(���ƥ�Z�c��l�v�`��k!�j�ŕ����,�̳3v�T�� ���a�j�_O��������:�+ٰρ�3TO653Y�#ne���#���I����>�v�tA�ZP{�$OG��q���
��� ��u� �)�Kj�x|{���Vߕ�Yҫ�!��7nLyo]��QNg��(&S��m��K���O��
��H���; ?q�]R}��or�;�� �3	E=���N*��DO�d��)t�sB\�/�j���Q��u��H�=��Fpz@U��;Q���VS��z�Z�3, OZm��E����yE�M�d�0�w���	i�J���~�P�����i��}��+�j��S���:UZ��jю�]��21)E}}�㌮E�$��&yl�Z(���1G�O���Cߺ������Y�GB���I�E�2�� ൩Gz5����M�Vf�D�
�?�D���٩�ŠC����d�*0g$�  孋�fA���Iމ?p�LI^W4�ds��|n�&�V#oJH97���!����4S��[%jU���R(�u����PǄ��⪮��:e��]�ڧ%�����Sq�ԓ�I"ޥ���D��Eߜ��E�`&?�{]�4^�
����6L>j�ݽ�f��ϙ�a�yWۋ%*6c�H��d�(~,��K�LE�4�~RQ�Y*�SR��"��~
k��B-s �)ݬ�R��W� ����dS�"��A�$o�����j��>4�h�̨���K�]w)���$�H/T���5΀`#o7+�;�h�d�5�x8�x��EO�D&������(:�1O�>4|�w��q���xظ�~'Ek�A��nƄMc�,v�b��0�Y��G�h�Qf�L���� N)X�u��-�PaN�q�@���i�n���#�R����	d=��%Dܗ�~׶��#�y��A�a̵��;Py�߂�\��>���aD��^-��jo� m0H-��20�by��x�ۄwD��_(��H�0���D���w�.�o���*Z��c� ��E�ԅ�f��XfS��$0�5nFL<�+|�.^��3"��H��9L��$Y��b�4Z�F�'~��*Zկ��d�%y����_��+�%]4%��4�Jd�[�0�X#]��?����dƦRa�z"߳��ca=�C���U��TBvh4�A@�^K��4�
�(����x���Amfَ�rWd�q}��S�z	NݜS4�\�N >�T���~�q>P�8�=�Pc��;s��חO[�܁>�
x�S�5�)�J�����Lh:���S)Ӓ+�Z���%7tt0���	�	����;v-#�T�Jx�ѿ0��k�܊n�'}ߚ&��u�2�{_��3]���&ʩ��>���~����Y�K�!��ڼ��ev_k��*=I~���+������`Ν���=�z�R
pԁ$σ5-�o�=�a��qA@�l�Fg7'��<Yp3ָ\�j��0kS�p�Au%xǌ�=o�f^�ٮ�*���J�2wV�$ �߲?���|&�}J�x�j�)!&����03�`<�M��]�I�D�^~T��T�#�* �*�Ub3o|���q��*���),t��4���e4"�rEP�&�X��^J��k���x���.��SF��^��|���[���[ʭ�=�e�Q]�^]y7Ј��S����理e�D��vB(��l���`���О��*�E������6;P �x�߃#-݇�<U��2O��ƪ�#�O��	ݼ�(��D�L`�����g#X���gM�H���ӳ�?�FgA��iP��+m n�-��)�#�~+�0�Q�U_�_�><�_J����sU>}�#���ƶ떢��{�5��wur��^�:"��wdm�^�j�_�nB��Zi�>M����8]�3�y����_v�B�,��>I��5�����M? �@�5��F���l�k���a����l܋��F���#5���K4�7��y��t���M@CW7ʒƪ,���M��#5ƻU�+|�Ξg,���Oܢ_��Q>��d���1����NN�`��+c\��[r�C��5(. ����4+C�jP�b���Ƙ����
4�M^W������4k���B��Օ�B�v�$r���C�Ē��`���?�"��>�N�פ�p0��o�pCk�M3�T�m�{_]�Ϙ� ��YiW��|5�-�ӪC���eDE�{����R��k�ύu��vu\d�IZd�r^�x�Q��H5��eLK;ES7&��nQ�����)\E����̓eUJ��<�_M>=dt��͡m�>�i�YwG"�0�_�놾��.&^t���e��\ZvYxrF��2笲jֶ	 2�J�m�o}9���X�3k���}�6pyEZ7�,��j���g`"b����n�����0��+��F8m�OfZ(o���M��Œ���e�T{��Z�Ea*+�K�et^�F�/�l{J~��k�V��8u��wn\�)C���9.�`L���(�Ό�́���i��L}f�&�r�`�^��C�Z�n���A����{�Xt>g"�3����E�O�ɯ�;植��6�����eD��M!	����]L�Z���;V�+�m�����wU)�,��SW}0�'A��RRN��AF�V|x*�4�X�+�>t�}�\����h��!�v�qf�EK�AR��Y���^�I��v���Dp�4�(��)���V{!{�����䟢f�S�I��s6r~r�/7_S9ʗWIZ�N�K��9�~=���Y�a�`���7��|0V\Ў�^�1/���K�}! �͸�dt���-o�U
Θ�9J⯕�G{!g|�g�S�&^|��v��q� 8�9<�`(;��E�#p�>ة�׽���`&��]�N\�D�9-�f���W<�������蝠d["���a��=��:���s��`@��3'����\��B��i�v��摑��$ȝ\wo1��I�8e\p|�["���R4�<��µ��,b����E�6�,�h��T��j�[w5Q���ԾxQ*4b����-�A�7���
��9�;X����'F�T�9��W�@Lbź���'s{�ѫ�>�fԾl&�DJ>��]�4Jr��[ξ�p(�����?�"S�.y�a�֪��su��Cp;��<�1�c��е�D�i͜0���n�ʠ�Xzp!�~��������1p���
	5�$U��	p��u��M�R�qa
)��~�)0��7*T;�
���e��	���?|��s\:�K���K���{�F��|�Gb���۪:�f��9%K��'|�/E���:We�V��rPa]�(�;:n��XߚM���@w�7ݜd�\����B�eJʼ)ߝt���=�#�AB}5�7OU���/��ڬ=��CX����|�s:����������E����I���`'A�����P�����{��!^d��I���& ,����(\�H)-0̹-��%m�ʱ�1*f��<v�����e��������眣
/�[�j��d����A��W�F����b�s�M����u$CD�4T��d`�V�-�~�&��V�K�S,�]�3��Ixv���/�7�����¬g����;��R����/�w�c#0ؕ�dlv�M���&+��q��w[��gk)�xy溝(���EL��q�,b/^ywLI���e�6<�*�Z"��菾EOB�R{p4qC��W��q��j�c?��=�6�CoY���L���^�ُ�/�z�p ��f�үbG��f�J�'#�}ڎ\��$�)\)s�����4sm$eл�E�[�u�ɸ�)�2�b��{bw�W�VVE����y� ��է{�Ò�z2����A�2ü��dl.�o���:��\9��H�4�rjL}(#^�kc����f-O�a�<��h̊ �+���ʃ�S���[8���o�4Uzn�}�70վ(öɰ�����<��y r\�kVdeqe�(&~�	f<��5��7k���4ğ!&v�Ȱ��qK3��x�}�b��ׯ="�:��4�؈:Y����ˮ#���N�S��+�]�t��9�����-7M�����k�qɛ����2�q[��P%���<�:.�P5�?�!�*(����k��2e�H|b�SH��!$&]���M���䛒;��Nh�P�����4�#^+���{�x��S3a8LE��[]��i��?�Ȯ08'LC>U�&nW\�#d��բ0���DP�N�4������w��Lv�A򸙌���E4lO�j:*hC�ڜ�(@�NItH��(��)�RZ������i���t𒹊�g�y�V��w�=���	0��)��fRw�^ڪ���v���j��I���ԩd�c���,nFi}K���K�H�Y��i���w$�E�� B렮�1�5�N{�2#���p1�f�G�N#p���,�=&���ؚG���m<b����W5�O���n� ���?����n���J�_��>n��b�����kI�Ns"oyt\V5�Wy�6�ު��BOI-���F���	��"��S��xg�h�0+s�ly��3����y4�Q�[��˔���{��_�6�]��^_��4� %N�Ŷ�7���յ)k�G��N*3����S^��a�2�<����]���Q^�
ӞQ������/K+WN�c3Q Hֈ��+K Ǜ\��-����$���E��N�5�d+g7rNX�'�G�(������~�n��p��TĹ�qk�D�2"
ǘ��D� v�ܦ黲�̌|n�ut�]����4���#Z�N	�3���Wwb8�\)���~�ҏ�7��\�;�f�ٴ�ıL�ٱ�/��^"
��b����60Q�r`���1�q�ʇ�ٚ��Uc�ҟA��L8jVrW����Y�>�d ��"ڈ���0��
� �E}2o�w��6�t�O.G2)(�)�w����N�h Ҥ-k)���:�¬|���a
2���A��ė֓�f�&y+��W:1�� Hء��N	X�k��<!��SH�<k}d�ѾS' X�����)����A���L�C�i�:j���[X	�FAK�⪢>��ķs�w��W�ԥ����@��ec�j�r��B �l���2���W�N���1�.�����Xڒ��YӅA�~���U���'dL'[�Lk��ݸ!�E��A@�KhZ�U{t�mo�?ڀ�iO)�Ve$[���<� ls.]�s��-�1�'����J�$l��Ԁ�tXYa9�g"#m��T�m����6
7�M�WM�C'�l2V�B:
O���?uZ���l� �c,���ƳV�U�Xᵃ-<(��u�c��D�m�R��i�3��}�vGF�K�UȹY�g����5�)��FԆ�1�@�o��r�?a���⟋����c��}���m��p�d����v��u]��q�9�C�bۃ3�lG�{�&{�5����@֘Iyx��^�]~���9�V��J��+\�e�;X�@�^%�Tig����>䧚{'�skv T�I>�w���>�L(����d�Y�/I IA<�j��O�k���G�!)��g`��;ru�֝�=ĺ#w)�I�;�������py��Be�d*��8�ȓ,�Ӑ�_wH�1+� '�
	z�̀�|7�8��~�D��E�,a� ;���d�0�II��: ~m�Qj�|�7�����[�����Q]��U�D��>M�BrL�EiF>�2��xv��*|fI������	N�X<(�p~o��4˽�a�]���,^ �fąn��
U�>����9+wL&�
d���x���y��
��U�(����0�f��o}��'�r�$j,#��y��N�eQ���^�E<�+�����}ѩ e}RvX�Ҝ������&��n>9�=�LdI+e"�l������'g{��s���8b�}	\+�S�*��E'.�	}}��*l6`�{X�W��Ƞ'�ep�/��� -+�)���UQR���McA����:T���H.
�5O˥g�v_S�k��4^N�(��xx�؊�-	��|���^I�kA���K��˃PKt��[����h���e�r�*����Hj)�s	�8�r�+Д6��xIF*�<�p�B�-gF'T���}����iT����√W�]�	l��}x�v�����~��)	SF�������V�U����7I�q0-ez�T�8`7�I��wY�9�� ̞���IЪÅ7'g`��֜�v�*��I�3��m�O�!�Ӥ�a���V�j��3L��唛���G]��ߘ�o��'^�<H�k��|���R�0ʨ�����Z�g�t��}�a<ʸ>�>���W�2j�-+�s%��`�s[�&��XQ�����P��{8�.2V��^v]Ք��\>���i�H�AY��;)*�b<�\QK�����Cg�\~��4m(�Y<�"Q.�0߾[�7�x5x�؍�4�6�^��0#��M��N��g��G��j7@��DG]:�+�'�{�Iu��Y���3�����;c��j��9���G^ʔ=�R4���z�Q��l��7�B�����X7��K�K>���a:�J�I+yO��ݵ,�����嫊�:	��X+��a�*���+Ԛҩu׏� ����In��G!���>[���Îl�$=ɔ���,��h���M���gI$�;-�����V��P�E�?r$�v/"IT,�Cl��x-}���DÃE�^�Nm��=t*�އl1�i��=�s\�a�h��cPI7UO�=�Ѵ�ַ�x�Ճ��v�MPGe�p��.|Y���!J%��:*�蝷B��\\-�����Z"oh��b
.j���^�����6w�`����,ߧ_m,����Fk��%}�<i���1|��-��YSw=�fםO����3���O����(މ_�����V��#�*� ��@�8(L���xS|4���7�?b���D�&%
����8��p曲���{h]m��y�?�H��6���{r�)�cڌ����htՊYX���
���n����;M2 ĕ�[P?'%F:��Rp�)���q#��p޵5YK��72�2!�?��k#}?w�/R�mC�M���7<)�=��wD���x��&��˞����t�UE�}��]>��"jQ��Jy�����gJ����vLK�?m"ɨv���G$��Z� ��J����z�7yi�	�vń_.��h�e�]}:��}Ů��NTL��O�>"ꑰ���rr9dy8()$`�t�}�>w�&��T8�p.1R��g��݊S!�ށ��.�^��c"似L��XP�N
��N�I������\*P}�l�~h��x�`��W�ːs�:=g,X��ۨ~d�:�&���I��,�����_/�A��Q4ؿ��y�����!���ؗ'��5���t/
^�WN�b����������ni���5�ʊ��q��{�>��*nvfgg0ɳ��8��=�Z���\��&b�hW��roU�<�������0��3yji3Ւu𣅷t���-�%lw�ݚLʵÝ�IxWZ)l�	��
1H�^��C�.��n��//��p붝P���o"I�,��kG:�m^����Q��X�'\����0}Gk�7ë׌@��(��Y�R�lC��#4��r"�];����������BU��	F�h[����_p�~x]P�{�� =_���X��u�����y��dg �#�qnEأK���ژ;Q��p|���+|ǔ�,�S2e��m���g��T�S!fx����]��U5q~���
�!���Xl�����۫�c���ǳ+F�^|d\X�}��i�B8U#��Y�1M~B����ÕVd~(�f���(� ��[���@�xA����"���\K�Ϥ�`����t�O@�,���DOUJ���+��/�hSQ
V�@ ��uH��dPU.�~֫�(L��zL�#�;~�����#��F���:Ry�y��fY+��w�2X�}PX���W�Y�����{J�sA��<���`�k1Z�l�y����߲1���S���*���w;і��/�\f4��WVs�D;�bw �v���jo�q�}�c]Y����k��N���X��M�_���gJ���������NT�(��Y�1:?�.dVו���#�Z��>g�p3�f�K�vhvo"�.f��
�5������~�ai�{i�_��-mE+���W��j�CB�}�KV0c�{zU���O��tbi{��<|��>�9��֫�W�T㍨D���xS^c���Dp>����ޞ�[�R�PD6cpsΰL.���]���X�=��`g��W�Gm}9U亚W~P�[�6s������I�8�ڰ�MTBg���]�b��?���+
/Ͱ����XG=]=�L�`���ݓ�tX�0�^��'��R��ʶT��o�tJ�����o�M@�l�*��gC�dU�ź��/��Z]Y���L�tn�m�n��Ӱ�����a�=��w��� �&4�{';��No��G���f�:��5���J&����{o�(S/W.���߉�J+YR��&���$',E���R�e�q��?���Yh��h4��N�l�d�X_���nF�RŹ!��~���Z�.ޔ���T�~L-�+�4 �NϭF�,$�K5�A� ����z��e��~��������X9�ks��3
$�v��!�q��a�k�+��P
"���0�j��֩�H%y(��b+K;n�һn\ܽ��M��.x�S�u�B��S>�t�|u ���TH	�6�$��Ŗ*yGF��W��z�	g0I��7!\����,V�pXxP%Utު�W�+A�PX`ʉ���N	���9�>�ӣ�@�p���������l��� �����^�p�ul��_
�CF��sQ��	����M��B�`�Im�M�b���LKQ��cYkU��Wh_�ft,4%H�׏�
(��1օ��~��`�������yZ�'�C#�^��*#B�:����
jh�w��"4�c L�溊?�,M>bI�H��
�a�-r�~Dbr�����>Sf�|���i��8�M����Чy�)��ZH����\c[ߛ��P$�����ڧU��-wi��1>1^�7|j� �z�ƞb]͔5��<I���G�d��F���%�\u$׸��9�����R�ٳ��4la%^�5�`��ڿhG%�%�^�ut����]j�����|+ʠ��� ����YB��@����
�R�iR���R{ꗅ��ՏknbZICb6R�%Է��J��@�c\�]���С�h�$IO�éY<�0�{rCv�Ŕ��>����-�^r�k"ψ
u�W�H��7�%Qj�*�&].�2���m)	,�C�
�/�2�!C61�?����s�J]��'N���loR�aoc  ��wTV�U���$�����B'�W�5g�ś���,i`�z�G�me'�wl�$�5���]�*����rqD��ˏ��5^'�*l��-���!�f<$�l�G��_.]Kz��p�)M�����i �i�(GK����D�z�ȝb��EЪ���.#V��~v0)�|7�r.*�1!x�c�ω�j�f��u.��걪��䉷2W>�(��������%�W�����pb����C�����Q�U2�k��� �4�����~���6E����Niqw��t\P �c�8 v���a+�01*U���ަp��7t����ɓa���}�����	�����/�6�T1t[H �\�lU
�/Vf�Ð?3�i���6����pMϞ��}�t�@�,���|�K�ӎb�}A#z��|��q"���胗��$va�P���� �c{�+�sE�6�:��I{�I"��������^��ʇ�L�F���*U>��\шCa�P�{�:�����i C� �kQ&%.���OAL��RВ<�vO��Hsk���+�����r ��&h�U��C��a����[3�bH�81�q�/���\�FEc4I����/Fɚ�!���n�U�^��]J��c��zb9yS[����d�n߅t�=)Z�u�"��l$��D�kS��u��T/?<����E�%Z������?X���EG$����ik���ҩ4�F5��OZ��"�U�!!����A*6�X�L� T��I���H����w�*���v{�}!/̈X�+�q됿�!蓊��<��ͤM�І���Ј4.jK��W�u�u1orH�Ʈ�6���3L^I���SCgT	4(�(+ �>�O����m�H��j�w`��c�Z�OSP����EaoJ�[P+%-y(�D���
ѓ��).Q��vVh��[S;�
�j��Ĝ�*Ix�4�)�u
������>Hn��/�Z)�t��zK["���)c³��g�j��"���G�J�a���xo[�sztO x���M3\}�(���b�Z��׀��#OA;��2��;��Ҭf&s����!��\���v�����\nBɮ4*� -)�)F�E���E� �_Z��n�p�k��sݘ�/W���g�Rq�Bz�"+����v�[Z]r!�`:K�6_�UR�m�`
#�d���G��D�zZ'!�Ը��iFdq0��IIb��e��ɥ�s�]��K��*��Sg��� �<�U�NG{"���]��rD¡��K��.��?<Jr��I-G���Jh^G'\���y��³�m�9,���n���J��5������j{7���Lrڹ�2�7��ߋ[��aF�v��/ºb��ڧv6��ͯ"_���>H���@"�Ƌz�+X�(}�N��8����\I��D��[������ip���U��t�#�6m\"��2�$̩��4nr ]*!g.\�����V�0Z�Y�𦻢I�A�Y*�m/d��/+��<�W�Qk�Y��"����U��𗽾�"3d�`ٌ��;�nD!�}Dy^�é.��/D�)S�TƐ�F&�hRM� ���d� �Y�G���R����픥����^Xa�J6��Ɯ�9���@�F��Q��K�l׍`5������6�ͱ�T����)���jƠ�(��fzP{�4Lg���[��~l�M�,�SA�{��E�-
@����>�f�r= �� a�8V�	��SY��K����)1�����^Ջ��F����<� ����)T>5�Ǚ����I�J�K�p��(�{:D�zf�f�oǇ�yQ��c��d���+\����K��@F+��b朄�E�L y	3y`�؋�R�B8"v�bvD�O
A�"��s�����C��"]gU 3�C��)�v�q��X':�=�Z������9W\�A�������uD5j���Ip�+�h��9�0J��,θ�n���}6YM9�=hk�f�2�j��
׿���Y`�̑*���=�(.Նf�&&�*q�
km$C�(��t���FoT
yD�P��_]P6���1���2!X��U�GC/���CN��E`�~~��
�����?��JN�(��J�x?'�T����>���=�s���E<�Y+�C�8��o)���娱Zby�$���#C�@{�8�ע��Fk�v6\&�Ny�-(��.�T��B
r`��� X}�B�gm�Gެ�m��r�~�����\p�o�j��$������q�D�%����]>,�b��p��=��֮^č�R�L��=C����׽FFwn�=R4NM��Q���p臨���@P����8����1ڡ3�A�C���7��b��MBI���ps]|;$��a���<ȃ#�ۏ�%V�"���� �+�|�=U��g���V:�����m� �9������^Sp����
�,l��}�q��,�TVh ]0�R�V|����84߬�ů�_����=y��4c,��G�U1�Ģ�;s�'.�㤌�	�5|"�q�=�)�4�I]3d!��]���
�����H���D����ڻA_������N9k;�L�}m�$��+iZJ�މ(�^�Ϻ�Lk�8�׽*
י�ʔ3������z�đ�;c�s�y�Բ��Mp��/=�-�ަ߲$�*��	s����X���Q��42P�`��%\zG߇°�/��A��UD��+�1<�g��򭅻U�!g��S0��N3����X�|W�Eņ�`���3��v�؞[�52�"Ůz�c��W�zIL��j��iJ?�w/��:"]�=4�*�ϫ"�f�Hk-)���[YEP*����v�9Q/M��?���W�Rޱ�;�?�VG)m����zF�$:����s�֌�O��m�[��*�U��A�6}�E��l	u��Ϩ<��I<S�T�*_e����FR<bP�6d�W��)�EN��U�q� �7"�ǀ#����`��k����ﾍgz�Ogl�i;Y��f����5�X�S��pN� s�(V�o5i8������ ��y�2��_y|-%�A\0Hry�Fa�?�	���K�)6�_sM�c��'��b�	e���3q�&��ʾRp��)%jf"j����W9%�`�1��f���U����Hueow�֋�y(�3�(��9�,��x �)S��Ҁ�����UnazT"�oO��?t�ު#G������D-����y
?�m��}�A�G1�%�eP^�;�m3����J(y�P�ju��v& ]�C_B��j �#��m�eT-Csw�m,>",�<Lr?T(��i_#>Y%�<���T�M�L��]���p����)�.䵬��6y��GP%�HרM!ȹxI�χ���B�W��2N���]��Z�N3��y]t�5x uoXa�&fD/��M2�:*8� ���a5���6:�R�5�Kd��&����!��)��G=:�Zө.fd�!�Y�W1j4D��/]C��xo�j��a��\y%�J$Y7�T|�<�G��g�7[-�> ��iVޠ|���e�*�~B~K�{e���Թ�/u�A���(D����Hه�f�Fr�sa�ќ�2I�e>��cJ�U�7aw	˃�����I����]�Z�@�^�Vv���,�(�5�Gu;J�2E��a&��&�_o��wT�pT�#ќ�)�{���H~�+��RE#����J���uÈ|��j��$�{Z�6L�5O�Cg�U7$��Ϋ����Q����"%������[�n���R&PC�Lc����bs�#��c�7�;~�Xpc 4sI�	�]�����ˮ�a�XK�)Dk�;w����"@���Y�)�fMTv���M�mj�5�ì@��wMS���J�����o-�S�|
hu8K�$�����ǭ�:�K7����0��rsO���
2
7~�1��r�9I����+,Gë���+��A c�B�@�Z� ���2�v\oD�AԆ��C��u�c����S�����vk�I��	;^����*=}�����@�/�լ�[uC�|�b�����]�H�of����L����=ѯ ��O�2�(kk�M��;/&��s���O�- ���[��<�+4��*��Х�8U���~9L�]!����͖!a�1�@x�!������a_:r�^z��sT�g}� �����L�e��kM����M��UG�ۏ�B��Xݽ��;�
���2�˽����b�1�{��!Ɍ�i�Z��=wq�:_��U諆�h���@�~B�ī`Q!�� ڧ��4�& ���nUz7[�s�a�d+��NO*V@��A�:%Џ���+�*inS6�΂�KH\2�]�
@)�,�q-$Ce|=YBD!��jz��+Œ��Qo����2��L�$�\�R9q�p�;C�����I��Pu��b���AemE��d�lǥP;������A_�b��qɘj��&|�orkM�W��?�}+	�Uk����]��pq|�X�����_�/1 ��������Ï*Pe�a(Z�a�y�Îk~%�vaγŵy�;N'C��?j��b�8���e̗N�����dq�Wc��e�?��,�*�aX!��@�H��߭ZO@�\�a<��)��qh�ylݭ@m�(�k�-k��Q��O'3�}�Ya�Iq�����\��뎑�0�s��ru��۝�vQ���(4^y/]��;�O��Gq����{���(lI��kv�4���־�"�KB�U�V���0z�_	w��{VnT�'�~1l���$n�3�Ea2q������;_6�$<�3�<�j���#'~yk�o�u�3���t��;�-�7��+�%��/Ub�V�&�b/WV�QEs���3O�(?���	խS��#���YC�+OW|.N�aG~Y��ԟ/#!�0�]��� Ӝ�m���a��w�#�T����z�<�Xq�����pȺ�4���&Z���{/��@�k�-�}yp��:-�Q�7�m���� �՟�E��ր���$�G���S�a�;Q���T4�K)����A2;8D�/2�.�3��:I���Q;�ܶ����p�f��!����`�Ӿ��8fI�㡰 7nCY��0�&�G���vȵ�ClG�q�S���pS��|�s��?�iBa�1t���J�ݜ�����3���A�o�$�]ϗ���A��y��_41�;(V�&ZEZ��f� o�����hi:�$�W��m��RK1'|h���3(?*1���ʐ��hl� Ӷ��Ĉ�$���bʕgJb�P*�}O,�O�U����߽㯄S�r��Ht��{\hK|��t��))�U��.��M�VZ��X
�-l�]�_����4WGf��iA8zӝ��j�u�[_�4��<�����מ:̻u(�?!�׸�-i��t`�ψ1�[��>�}�¸�.�L�Ѥ=Y������
�f���	��w�� )���#Hyt�Z�@3>��a\���%I��s���Ί�\�E�ȇ�/O��߈�%d:U�Y_Pa5��pV�V�h�f�p�2%���~�
u�T#��ZY���%`�|tn
�����j��ͷH�m��.��X)��b�UQLQA�x� ��K]�|�8d���!{�7�L�ݪ��OQJpՂ$��A��l�deP�]�A}����u(;��2�oE[�����2,bҾ��x�=)G�[��B@WV��2X`	��C��s�yi�M��T& �8�m��b-�K7p�X�(rmf�PyE�cUL�T�R�g�\����iZ�E3f[�L:]�`?�<�Gq�����j��/�4�����������=.�[�0��T3U��)D%u��-�����u��R(���l�b
�#h���7lq�3�ذ�@�C�3�qPea�Z�h��͠vo�_�=Y���=�u��E9���N'v=���?�_� ;��B�)�Xօ�j��r,�i����cPgV���i���p�z�Z��E���dɊ�@����ۑy��\O�Ƀ��w�op�C\k�H6����7������J�������m�K(�(��;� �#�DA:v�x� oԶ�/�u)�顿&�~<��I�|	s�\e��(�á���Ew�`C>,��K�t%�`�M��#��1���N�˘T�����L��k"�-��P�N{M���nw�$�}Y�X�-�T��x�/���7���������T�h�z�5SH���QV���"!�S�%3et���c����!�pV�U�5��_4F)|�4���U���/G�gc�� ���^V�":y0�X�����ºN#���U\����2S>Ӆx��`gv~O�#=9s�ޯ��PJɫ)���0���%@����O���Qsa�;3��K��l��H�A��~d,F
Q(L�Ԍ���&_���y���B��:l� :aA���=�=1�<C^�� �8��_=�^α��0#m�-�y�y��ܘ�AY��|�v��i�@�����mc���%�m 
���!-W��!�˳B�g<�&!������Qi�O�� t�
W꣛�eO�����8�P�[#j6=7~c5�}�V�͊�Dd��]�T�R� C��.��*\.�m���Ԇۍ9,<�F	��0H��=݁�������p��Upw�혔�~�;^������N/��뎂"��C��M���W��B�ŷ:���<�OY�6��q2�G5K¹��U����S��o�$[�RN�
��&�=����]�^)�
:�8���m��A��TT2#��h2���i�@��WQ���O����}�+}WE����r������%�]���s�������;�������"k�i�� eh[ B��Kh�C*��S��a<�a��ڠ=��Y�������ʮU�U��=u�����+>����D��c�`���V�A�S�#�QM��Ԍ�ٷ�x$ c�T��0_vQ �Y��d������˩��*M�e9d�`H�\	"o'B7��E�\֠e���_j����s��aSwR����!����ȑq���l��ݪ�)y\��G���i�S�#�,Qg���s~0-��L3�6k|x&�,��E��v��y	��*
o�g4��c�Z���Nj�Õ��;�����Qq�<�T��G���h�"�a�dă����.&Q��GP�3��m&�@-��N�֗H8���>��g��< ,�nwǛ8o 7��r�Dq^�פ]o�Z�F�0],�p�45E�Z��i�O%%��	�0�;<���Vn1TҢcan=������G0⤲�����YyټϚ����@+��`C�%w��;�o���_)����8εy�6W>j#8�)7���G��?���Ȏ��j@:-�(��;;y/Ш���\�"����Il�dZ5lv�Mki$��D����0톅�q�"����qb�a)w#�K\=t���e6%���PTx�5AZ�L,sGGS�S�.U���Lm��������L����d,h�R����[aր�,y��[>Iz	ܽ�p��dF�(��Ъ ~���|"ǂ�[���B��ݫ!����٨pD�4����aY�Y����ǜOl6,�[�*G���^ȭύ�n����(���r4�4�Х�ln�nQ�h��AT�����on�N�@���"�"`�d�4m�D��fh?p�q���-1��%��x\��t2��~xh7�R^�Z��(�
"�_I1-8k�,D��)ܾ	��{	R��\��nm��qi��Ǒ�J[�����k��l���%tH{{��;:"���mhRϓ��il���k\��Ek��o��f��k��N�jȅ�j��ٸ� �{���~���Ӏ>���iI(�[������h��5T~Ss?�#�@#���s���0Z��{f���������.
����':a͖��g��pPE�˯pA��i�3�}[� ��е'I��Q#��`	���v�O�c���O�$W��d/��gJ�:�
j�hcjnڞ� �8��HI�@��S��Z�si-�pD�>gO�*�W�jII *	]J�-�R��'Ý�bP�q��ë�N��l��K��=�ޛ4�.2���*�����.+��y@"����R
����o��E�N�RI-�?��w�<~��	@�Z� ��Ӕ�����a��aa�9�\ߍ��=��
*i��@�����=f�L�	Y�t�R���c��^�$e��w��yVw�pw���z(Wښp�L�o��M�)���dŎk�h���`�b�c�|ulY��Bu�5	�����R����p��APV���������CD�ԓ��gM��.�,=%���0�V��V�,w��٘ZANy����*����f���[w������o9�������k��0>�/��}Mΰ���%S6E0��j+��G�#��c����	6wO_�	�䴘�TY���L�5�WHoB���|J��s�Ĺi����m(�-�V��A�4!�9��S'��͐�er>�=�A�C@|�����8�a��t��C�.K�f��#���w���kV�P̈́Q,:���q�Lq�Q���@����q%9���j�%�*�W�RYV�q�*�"�ǐ^O�z�	O��"�l�C�Ul�G.m�7ༀ��y���_��!�P�!w;������G�"_�˝e��h��+#��'���A<�n���4�(�j������heV.���[��
TR�A�q�k��U�C�Y�-A����
J}&`8Z��z�!�,.��6��{NM�j�/����p�{|tI��6.��r��Ef_�u�����#��?��h}0;܃dEV���<�L��ޱ_Æ�|LmJq�P��p�`#�IF�B�]d�,3��~�p��nb�*���h$Z����'�K����-$���[V[��s;����K��.N9)��<�ݯ9�BI}�W�����A�aE�����\�x ƕm`�ְ��Xb_F�/���O�R3���e�jH���g)�R��t���*�QH�-,@��h��ѝ�2+'A����G�%�����=9rcWDh�@i�څTJ����@�v��ί{�k�/P�;|�6Z��u�ը�b��c����ǡA��q=>a�ܹ�V͞&,�G�7b*�\�(��&Ħ
"ھ)��j;�){��D��,�ˏ�J�}�=�F�@S=/R���s��G�~��i|QV��|$z���%ï2ޭs%�e;�-�=�m��
��*VS>>Մ�p�
8	1�?��泃[c��<7V*>�?u77���ĝ�Fl���ݔo�z�9Rn�-���|#~���!U�G�3���ґ�I]����>Us�5� |�#!� �8fe�$?�e�y��6 �2K�/��3��O��U�)L���d(>6 �N�D��� k����a��̍���x�2���#�!*�d�F����X���ہ�`;�<��us�˴���U�����3��I0��|;��K�g�&Ifp`���a6�>E'Mx�x`s7aBXc$��V��wM��jC� �#����u*P�|�~�%+.@B&�֢K�=��:�Z�n@ ��y����5���o㣙i���*����.Z�_ y�*C=S��%e��6��5٘ot���]�8��1[~A܀O&7��H]	��6�W�1�4�A��_���el������-D�ڲ�S^r���j�{)2�|��G�;?,�E�Y21t�̇���W�Wg�&) v����>�ݥͭ	��zh������p~�V������v$K�\�]�G���?~>[�����u��� UAd2L���e�Ҥ�yo��ȡ�lز��;�d�����윲�TF$_}I���/�nDB%�n(��djҪ!���,��W����b����EV2�a[�\*�8�m��~.f��C7�S��0�-�����L%<���*Hy΍��05�ߐ\��:�n�`L]	OwqPr[n��ڵ�6�kfП
Ҵ���V+��lBuWkx�y�x��:x.�N)[�dĩ�@�JJEfe�Q=��*�uhi'7�x'K�Og.E��t�IM ���g�௴�.~L���+Dthןi���<��Ջ��1;P��'� �o�Y$�e�EI	h�)jB��زП��4��%;[[�\w�C�`2��B�w$|>$�������r�F��j�!t���P���~����ۦ����K���z��7�-��5�c���C���յ�E�W�z������rڐ���ǔŽ]}�ӾV�(�U#<�@S�G�1���P6�aP:�d�ټ6�[�d��l	=`��Ggz�?�U�<Y�t�@�d�����CGdv���!�����
E*#y7o�{;5c\��d��T�����0��d3z��q���&�#QÝ�+boօ����sa�m?P��j��}�U���� �R�SJ�c��x>߼~���
H���e~1��:i1R�($@P|���w�ʀi���&
»(<e�⬣��7��u�ֱ�9���Դ��(_���x��,��|�Є
��ݟ�Y��[�ճ4�Ma�&�~�W��G����ï�{�z!:q2<�(y���o�řLm9�\�:k���Iu�O�q7
��}2�VM�?&{n�:���#80��
���������/=*�эJ$iX�S�ݶRa���00��1�cT�-h�I�PhԨ�X]�pt:h��%��1;f�k� ��65-�'��F(�q�[9���0��C��d7ۯ�T�'yt!陫C������Č�X���].�� ��Crr�?��9��������U5w�9���l!ֵ��|��~(�KO�OMa����YF?w������jj��N	�lD��
L�Z�xP��2͗�ٷ�����[!�u��X��b��T'��S q�����ټ*� �p��4��S��Y*+�	ۏz�V���N ��£1�'}���ښK�[ �w�|7h�;'�8b��;�����e ��>��gS�.N�j�w0���E�|9���I�E|�3`�`]�)`>T���Bw����i|����灍?9��G�2�aL
�a.#+l
�W�����=��m�� o�0�6/�&��h�N�BC;_�.k' ��F�&iA�b��o��k92�b{�<#}]����s��Fyd�X���RU�N�ucf���E6L�l��u�9�
�i({�I?:n���a�~~+�j����#=4;C���D�H�k�d%q�'#�Rh8�v���4P]�"����#�5��j߷�ѕ��Q��������	?���Rx��L��;�B� `=��j˄h�M6��}��I�QB�r�-,G�u���2��G�L����''��� ��&��RC.�gj��FB����<~���5��e��Ƙ�����H����b��P���m��'�7ו>c4!�"~�ͣ�Y���Ρ��ts��S�ͽ�Lݳ"؉ft ���x��Hw�*��TM�5|7�c���q�ݴ�TGemth���T�IT�o⶝�<���ţ��j�.�&�("�)ԝu4z�p7~�6�4{1��]8����AtK��#�+�W04�9Y�EH�{K�+���d���&��-��*�<7�k��)�����+<S�%�R��,����z�¹1Sn�+A[��ߊ�\���2��؝{���Q��~���}[X�˿�i+]YaDu9ZP�D�vI�K��)��(�t�ZI��^�`��r����c�k&�W[�Ï�q�d|a�7X���/�3�������l����^��a�ޥ�ށ֊��9/L��G<�bob�*�\qxn�݂�XG�W��C�bh@|i#�?ȩ���Ј��m����� ��<�mz�PB��*ޅ>���G�Q��n!�ɲ8	�Z��#��:��Bl��Ά����S��	�4zr��6��b}��ա%��$C� ��w���L �Jy?Զ��Q�������L,r� ќ�Z�x�`��\�g�����4�m��J�d%0��/$˳�w7%=�DSSjYO+C3����#�~��{�O�B�W��u�E���A%kA�V#Ņ��n���z��{��|/�òli�ʏ^�{1Gڧ��9��!��>��Ks�@̬�Ȱ}U@*OG���Y渑}�ַ�S�NA�/I@0�+�zr85ߨ�{����w{^k������S�o���'��b�=�{B� d�t����`? r �h9X}_���,@p�ZįC-Ғ�����֙?�����|IT�p:)��j��+��{��3�5��ܰQ�!ΓF��ȁs�,o���q�+}*������bģ[8�ڣ��ňE����/�r@�='�#��2~�'(��+����doiiq��DHT�ܳ�g*��=�B��{�L���G��{�}0	q�h�Q��
���HΔ�7��yLfKX�*�S$��R�`��}��S��y�i�Lr�1��$�()�@$�[T{�@U�J�z3�^l](c|9
C��)J��ŭzy��+�)7#Ԛ����`��2���-W+	C�r�^r�gaE/���D�F�?�
b��IM#t�ng��ڤ3���u�-"��f��#4���U:t��:�j����3åT��AY��W�y�IC°=!Y
k�Sb���]�,���Qw�uWA[*�:�����|J����n�YPYE�g����͠�� �$����i���+���S�|�[��ni��>jX��_'���'r��v�/�-�K0�9Sz�s��܎�K�&=��x��*�X�E�J��q��5E{).jZ`sc->!Iv�}�M_n�`���[7]�ɾlGH�U�΋�-6QI!��֔6Y%���[�.�X���i";����s�-��f��4<�b��Q���!��`�|�Q޷�wm����G�n����)�̀��	i��Zm�H-�m_Z�*w[�f�^��$�0���N����u#[9X���w
'�vV@������)�-���(�g�i}
��Ǉ�?'sT4�Bﴑ��rqQ����ey�Aj%��f<�~�:�H�b�W��R	C���d�ۻ~2fm�TB����o/��c�tW����%6I΃����]��JH2i�u��֝0�����Y�T��W~,���MdûU�B��N�%|1�#����K�qT�������ؑ@��%-��;;һ1�G|�G����*B�!�h�$�{L9�Z��1(�Jbz��"`Rϡ	B�c���Cڶ v%�I�Ӌ8[��rZ�	\������{xQ�W;vό���N���E1���U�v�*k_v�Q��:Z6��L_F�m��ߟ=an2�K�͖("�{�����iW�J��an�'T<��Y:�kΟ��W[�hFh���n��w��Q�}uq7���h��1J��̻9��B�n�%4G��T/5.!��_���l��H�N(��v1��Sq��	�b!cz�Z�ZC ��9byw�e��.���e�@ev���fo�@�)���|����l{��"qr>��H���[���*��:_)�	)Mܩ���[��^�V9�\D}e��;���mlo_}�J��=֕�+�
{%ҵ�y�HF)O�8�/�wz~���@>@Η.ُ��C�:��&�(��?m���Zߺ�)HI��Qj�rR��U}�:��`�*>5�٭�B�%)�,ʺ���kx��EMX��1Pu����o\���C�ڛ�g�����}��ax�� ce�����'��{q?��Y~xҶ�X�̤#��C&�VHۺ����{����r^a)LŴ(�_�ۜ��z�w��7��\5���Vk/��n!n'yn.toe���xc=S %t�c�Xr��\F�).UV\�
��ݔ-�h�� gR�^�����Y��g�i�(�'7oƦb��6ʺ���5�4(���R���K�=�$-6�v��wv��W�b�Q�O����=>(fN>2Cs�Ù7R�Ѩ�ec�����=ci���W��O���/�)�qDT���N��:c��p�{?Vn��$6b�����o�Q_��` lbt>�)��k'12�`������۞@�[��`�/F��?��UЙ�V��n�L� ��t�n�R�Հ�ȼ~�0U� ���������E���(����˿W���7��A(��ۧ���\�_U�����<�"��k���v��E<:r��1�Px�(��\@j�+���뮷)�/ ^	g)$B��έ��N>](�|�9@��؇��M�e}7ch��8��r���:�>��O���Zv�t]�O��,�>ß�� ̠�a��;�_��<E������xK��08:���m��%�#B�lrn�s��c&[�v��k�ˢD�'��b{+&YBZ0+1����q�0�2��Y���*Q�|3���4a^X�˥9ז�ǓG���n��|Ѥ̐Z<|�l��:�911�B�rD/���U��N4�T�`߷2Xq����)��g�J��=6ˤZ����9x�<~�\Q��$�V�KJ�{O(��QȽ}WB��T�hԫ�����Y������Z���Dq��^���#��[�T�����<K'D\!׍,�J����c�����$=˗]^��Q��6)R_N���݊��3'��ͱ�Kv�:��n�FM������p��=H��f2W!�b��5o�e���3W��գ�"|������Z;���AJ$�!�������<��!�>�D%^��ۗy ��d
����{䣮�s`��l��@9�`VO�����ar��V ��_띶�~��m��o���x�_��}
�s�tmf�i�m���d�ճx+Ƿ��%����b8tԶ��K�A ���^��Tr�af��eNa�X(寬�6�<K��u���Xa�|��p,�	bn,>��D��v�f��
ȋj⻹;
������4Wb�Į�ʀ
h`eþb�*�M3�V�	�v�gQ�Ɩ��l��M�_��u�h(\}�b(IPigH_�����_6�,-�Oy}��Ad��a��r6ԕQ>�)�w��(�w)|�1t\B�������}�q*-��h���f0;� �����+?^�7�rLپ��dE�/�%���r��3ez��u�����;�toBgL����b�Gb������Im���(��[nr�/�l?�U�� �+�'��#�}X�LD.�R���|�$I[Bн�9������_n�y}�K7��\�m�%LxU-�ZRo"�Skb-�W�Δ�(��?^!��u�?��<"��On���PI��Y�5�r��<"f�t`:~q����(���p�MN"�l� �$`/��Zmv�Q<�Y�E ��G�i��EH��9�X�{a�|5���@��^�Tŀ>���'B?�1^[Iۺ{���<1Ve`��r]�0o]1\d(>c���>�1a.J�':�����>5�>��Qf�h��qA�EFG��A��[Nd�2�la�Z���d�3���I�����=��}$��򏍴�*����Z�9��uX$��8H��[s�EB�x���G4ow���~�R�����&\:i�3��#l6��4��:\nssF��3��;�n/���Bn�x�(�Y�Y�~�4�3�Aށ���� ��n�,?�çp�k�a
ZO.�CB��)И��O@��9.m[�<���@�o�gJtf@�=���.=�)5Fq������5��[$upZ�[}�qc#��m5F���M��Y�J��a}�$1xd}p��,�6`ɳ�����:1�~�A����>|Ԋp##!�-}����<tV%٥�{��Hry �m�5��ձ�0a���`j�>7.��,j�0S�W)vU��\-�R�r'�������3�Ug�c�+������I��S?~��F�h�!����=�t0�h�4�[�{�q�KO,�m7}L�ݕ�l��}��Bcq��-�;��Wo�����V�9+'��V�R��N��S ����n�e��H���50G��EE�t��s��P}����3|z�]���
bv� 2�N=��� ��!t{s���䗛E�-�7�y4��JE�-8��b;; [�y�Q�'�({`G�@��6����%;U�l���U�� ����6h�A�����A:�\���;�����S꼇5����ܒ4���L�6)�����P�xq�%�G� |9�x������x�W ǋ$�Mm��h�%/E�m=��j��ܺ�*��Q��xcI4�� z
��Y���f���s#/����`e<'lMPj~�ϕ�p���[/�V�w�[�ӓ���g7�w�g��'��L�⏜7��a�y��X��r67���
�����5��X���Y⸻v:�.��է���ϑB�4�E����e�P�BqZA{�N�}��8�m�#M��p�����={�]���`lW���>~���M�~^��wF�������U�gjK˕F����W/�z�\�Ow�ҷ��
y�)����l���p!�t4&\��sǂI��Zf�n�:�D�ɺ��￤��mм�-��%�.=�L��t���)����F^�wR���;���lBd��<�]3^�ߙt�{ [5���CV��	�����0�jլ�2]N=s��HN���=	zRqBTGE�@�v���~x����� ��j�}Uv��_4u;��6�Tx�<�pk�Q����jHH�����G���zIɌ3��+� ���$�����0���H! �-{.���I���z�'e��񺉖�Ɉ��M_*b
����&�YpW(�PK��#r>CK�\��?y��mYWJ.N��ǝ��s'7?w!gt+Bb�א��7�L�=h�=~�Lȝ>�g���-;�3��<�'*}��9X �W���G k�����}��������ʊ�����9�rr��B�z��3� y�حn��p�S�ӕ�b4��mK3�OSlI|�	�9�	V�����K�fUH�t���	��'���/�ܯm]��v���M��ʴ��;�+(0	ֶ�����?��td��Q�	9p�Efe�|�ɯ�xh}�7��U��I���U]_Q������!�`�B���=G��g�U�E�0����m���+k�eh�.lB�5~%�?X�豳M�«$1Ŋ߶ �j�1�������� Q�]�u`MJ�h���lc��^TX쮠�2f��e��)���4����O��|�HydϡR�"ܽ׀�o�_�qjzsh��6�����,��f�Xｮ�WՁ�t&-�+Bj��ym/&��{�OM��r���G�qP��<R=�
��4���D ��ׇ�#�������Zs����-C*{�1�`�x4���y�N��0U0�Z:ځi�	.��匴���l}-Z!���Y���I��IE�'�Zi�uº�4�H�Ϡ���Q ������`{Z߆� ��@��s�jKU�2��+X�:���R^��H����c*syu�l�%�sk�����著�vf��Q��L�`����g�S�-���'�y%�V6ESR������u4n�>��,����

~"�ߏu�O�� h��;`d���m&�y��
>��^��u�r�7,+�zB=�؍V��lvM�R�P��v�۱Hi/�*r�h���0���ۄ�b�&���u�ļ�Y| �il�
Wdi��x��:S�JIӾ�o��I��M?g��OzJ�e
�?���џ�q/\�\��g���k�9�4>�-^��p��r�z�_��,n�Yi�?@����ZΙ�j�F~����U��K��%�[�?w8Q��(����PhIS}���k$�v��e��0�O�8[ =�g4R��]r�;i�#^�]�L�e�{H^�XΠ��mIGe�4��[&�a(�mVQ�^Ab�b�
��[��3�*��^���!�P�-/h�W�,4�l��>���RA�"�+�&��F���pZ�l��Ll^Nw9�?b��鈁�>����B�$���dݡ�V-�O_�L 9;���0vI�H6㿏1���t�ΠN'�0~e?�vr�b!�#d�}�~�T���LY�?�]�a�򑴷'�1�)3 #��&=�XdFbT�T,/疵X���W^�RM9�q�oΛä�;@6u;wʸ/�V��)G����+�Y��rZ������s�g+�n 0Z��X�N����h�q�J� ��Au�A%�lֳ��.�_]:��ʱi�܁5R���R9�����ESޒ�����:u{"�H-ڲŷo�dG�)i͏2.)*.n�E?�I;S����&�z��ă�;��=;<�T����b�:�bvoR$KBx��R�S�	�ˢL�0�rr�?���0vl#�}�H������@�V�+��f��4��~��3���K�<�m?j�&E`��m��&��������{ 0�N�h��F�2 �'�{XC�U������Yn��?��o�@�uX���c��2�,��> ���Il��%"��Ю��/Àp
`*��������� 8�_n%A�4(s�,������y������e>����{�� *��v��'�x���Q�H�JW�Q�(Pt\���̓��C�U<���G�4�9)'����F�x��m穟((]tފ�:�k�����r#(��ڵ��
hn���EՂ������Υ�y R~>e�����:�����0J*�),���򛺞)�3�y[6�`Z���˧��UD=�E�qw�'�ؗj��fU�BD�����k��k�V�����T&:�u���I\x%��� �ư�A���(g�7��6�a.��������M�)+�y}t˚&��jºp�@�z_HS(dE��^?���6�a����)P�
��8��w,�G����&f	���M��vl�z�F9w>[��W��	��5|��)U��2�Iڏy�V;(
U`�˽|����_�� ƽzU�&9S�r&�
䘜�I��x&TNIg���b2,I-Qb� ��x>dzXȕ�"mK���i�S��ȳ�ew��L�y�E�#d���3
�ț����A��l�Jz/%_+,���_���`���jn�с�����'Ia=�iR��|QBY*�?��9q�88vs����0\�o#�G�,7Aϥ(�h�.����d��5V\�u���W����C{�̶<2�M����bL-|0�u>1޳ӱ���m�]�aѵK�C��{/���YPu�l�,/�0!N�vX���;��J��W3弟:�I&���e�o�9-KO�^��]�����9����3�8�A4EV4�">U��zԮ��1!�'7����K��Jp!�0�
&gh̖�?�9όg�u��1�i��̯��F�A�X�Ps��q��o�44k���F>��-�ؠ�/���*��*��@0�m:����M�B�2ϋk���"�
I��Z4�?99���U�x�º�O��ä$�jt��8�r@��P��ᕎڌ��\��۱ �Ign�o���Wg|vH���I��R�����A>�e�Fc̢j��� �.36��m�V,��(���1���r+��{�/g""�)E+�
�	W��tTUr�I�>E�QRM��_���Y�&Ps�<��	Jŏ� �"-�o8e�}pI�@[U�h��n���!�+^G���_߈���0�Tp�|�*�I���pK�B�z$��!�Zu进����`��7����DD�v�w�P�8�����3*!L��v�`�Q@%�@O0B�^AIas���wz��Y��H�AG"aF�GR�R��:�9����B�Y�����[��o�IMK]~@!qvО�>j��lz�}��77�a�����V����J	��iJ:1a�������y��:&P���i�?y=>�t�Ό>��
4f�W�UP�Ty����4�jl��T �1>�f��<f45xo�$7LlL�vɶ���A~}�;��u`����kPA��;�=�	=��E�)�3����;��̾<'�.��Lx��޼8�����w=Qx���e8�l���n�j�:�J6P�M���Ƿя�Ss�D�T�0y����B4��I,z��A��['��)���dN���:Ξ�?rᶵ�2��B5UX��j_������ti(#n}5es ���C���ڀ�݈(�	��;�jy�G/J]���AO�K[F&,��Q �X�5��V:Ⱥ^,R��ZR"�5`Í+l��S�AE�o���mSY�q=~MV\�A�����ǖ�B����~!�ق�s�	S��%��;�b@Zxt�s�^����Ma�&*�0�\w��L����,�$�- ��)�`18�guS��`��d9 ��'�5u�^7���d�Wc�q��\î36�)%x|Զ��@;���:������:��"�L~&#'*[܎��WOӥrL�V8������O��B��%Q�p�^���� �Kp�#헡�.p��V��������'Tк�8�i�)J��$��8L �+ep'���=���q�v�8�F�~{��~sg�W�,���nt֡h����a2(b�R��<`�sw�x�bw��� " �F�X���X�N��~�w�7�nBx@�=��۾Bu]	�:b ���2��r�A�~*L�R���a3H�-cw��8'"��D���ma'Mg�������0v��#��A�^2NI0<��pC5��]s�Q[�/���Wy��C�!�#C�u�mu�;_T1�F����T���-Fy�[�T��|�:q"��������m��u�]�y�:�Mi�qٝ�T�O�9��E.���Ļ�{ipo� �h��� nƣ�]���śpB�ѧl�aGA���{ ڠMc�Y�b؞�;3���U�����Y�}R޼̮��S�#s�|��/#(!�v�˻��������D�'�w�G�t��4DJl��&�t�h6�(�`ö�� -P�<Ǆ�WR��?V9��=��v�i�zj�%�Ȗ�	d����r;�~�  Q����M�2�}y
��������xA�q:^@�?
З���F9Z���ש}�I�M�W�}���˕��P@f�s0����}�M�^u�����]��A^��q��������^R\����_�َR��u�����FA�!LN{�Ok���Ͽ�h=�� ��|�Rq���]5�D,6��:IF�9!��s�W&���R�ɑ�8]� ���:oCv�tn&9�|��\8��i�����<�T��fZ�?�|؁�HP������B�)���\q/�s�q?�:]���c��P�$�Y�`c��s��{KE��:KޡPϪ=���X�k���f��"�D�V<@�0�\�=�=x\�sv���nzS+�P��ٹ���\(�UPEk�|Zn	C� �
~�"��n�vz��S�O�ep���|�=^���f9A�rǒ���Be�@��5��}�{M׋�d�ۋ'��{�W.��~ G�X���+Hl�;���x�<^���]8�|�k��טh�3h����u_��;N��3'��o�c�l�b#��ղ��L"-��Oa(�,%�55�����'�Q�O�7���ΈJԅ#q�r/1��?H����+�J���%1�xS���^+��yc�"{^�4z*��pI�G� ����
&}�l�EL���,^h��{ñaG"�d�b��}�چ�<OeԿ�$c�y��9S�Q�f���4���Y��j��ND��~�k,��ӴV��L�w���|��/e����t`��gd@�y���)Z��J�y�,�%$�8ϋDv-��T�#�?ǘϽ���c{_^LYP��������8-��P�=>�\�T�L�+:�$һ�������F����lVE/�:̀�	3���tj��DAR�-jo���i*���Mo�>���T%Qݤ�v������l�=�U#����,�ʓ�Y�	M^�|i����<�}^�t�����7�(غ��ܠ����rr�E�j!��/��6t��n,.���뻻]S�<���cW�N����l�/�6	n��R`���W#{+�/ /��g݈�^�m8���-J�ϓ�f��ҋ��>���"O��f��X����#���Os� �c
����t��y}U]`* ����.v=���7:�b"��=ǵ�
�
J~Af]5~`cB}J�7�$�)��/������Ș�r�bd���%"������`�.��%���'�o�	�+��h�Ǘi~迏�����+�n ��U6�]��&�׸�b�r,W��w�6ӧ��@9��&{X��J��{�: x C�쩍����@�$(�WW��!8�4#�����?(zqj�lt׃a�`�\�g�n��.�>�cd�h�������
֪T�k�:8؜�}7]:�<���1��L�V��n� �J;ۃd�jX���B�k1E�n��E� ��Z��)���VX�<�b#Q=�~i�S�0]�e'
 ��j��k@�:t���|䗂Ncg�����KDm'?�J�B�jE3���rF!���y$�|$�A��X��*ᑸ����'�Z�����밌}��6g����Q�D:ͧzN�����7�.z�"K@!�N�@C/�wk��j2�����{�>l��
y�v-��+%BZ|Q���O5��C�����V͗��;u�'n9����O@/j�^\o��$W��߷cO뢦<�1x��:QWz(bܘ�&߸ �M �,�a'+��NL�ty�a}��,���F�1)2���x����R�5��[��Hs�>0�GjG}O�C�;��gA.���eG~e����6�y���D6#N�o���N�j�A/�++.�z��=�7(��@���KkP&tN�L��\���K�ol�)(��r�U��7�u�Ohe��M24h�@Ή�s��FH;Y���>Ͱ#CB�t3W_�>��0�PE�'��wF�N��&H��è@ϰ]��?!U�8GW�m��W�|���RDP�&���k�I
=Y�;Z��,�� ���� ��y���$�7_�;�s$c�f�s�_��&9��!��a:��	�#�
K���=�qĻ�M2?�%�� OV)��C�P�TXs��,"%i�ݾy���ne�9�Z	u�}GO��	*EAq��^��Q�^��b��Um�DT�P�-��e4ނ�h܅$�9�����s0��U��V�qG��Ƽ4�62�|ci�2j�r�l,���'��	4��S�M��>�W�-(����g�Vy��=�l�"����J�!.���Q~rU�B�N�ʌ�ih����Z��NY��g-p�<�ѓ�o��g3T���u���"$j��I�gG�t���o��g#��V/�<�����X��+��s%��4壔Bu$�rй�~7P�ܷ6�Z�o��Vn�M���wz�r$u�5��g�~l8��Qy���S�
�2�D�S����X�5:T �|��%v�]?N�o����s���ݺ�md�t�|�U��?��>�7?4� |��3�t�~�?���\=�E�w_��w?��T)t���7
kWlc�$P�b�����2����}�������2�ig�	A@"�����z:�S��7%PYN=��j��Pս�'x��[m����o�P��b^0��L�؍���ՠ0+OO礓�MA^O�E��������SԱ�
�ɐ��.�w�=��&-��n����5*B�Geʯ5�7��"�z�+��ݶ��G,���m���mرd��(;�7��2��I��d�9�`m[��5�F�|��N:Ng�Ÿ$B#?���+�ҁ�w>�ѵ�D��O���#�R��26Y��� `-
T�t,\�+~ŀR>�U2��yI��������3��6����3V��ܧ���  B0~��bE&�~Hp��u��d�:�t�̋�΍��w!���c7����{����6�Q9yէ<+����}Z�i�o;���I�U{R�mʅȥs4��.����0H:���:�g�A��صs�2�k��0R�?g_i�mU�X�x''G��k�ѬQ_R�=��N�%bb6`��ȃlH��)����&�D\�@�p��y���l5�i������[��s쇦��?{m8Let�
�����D���'��4��1�r$zbwO��a' UO��3�򄙱J����o>d.J����Z�c�˗�{6yu~�9 N�E&ٟ��u|'�|y�)����A�R�(IABj�CRyҫ��m*��B<��6��.��.`<I�F5��}�h�o�����]�H��t�f���?�z���Q�z-��<D����
�!�@��R�������З�����g��E��Z�S}B%Qqͬ��<!�=4���B���\:���f `�
 H����{�H
�?��W4��Q2�Ɇ�]����z:�V���)�wv.c\ϭ�Ik���Z���EǀT΃W����	�%����4;�Q%HX����u����Ч%�ģX6rW��|���K����_�k�Y�������@iM��]���j������
�i���7{c�nW���+����)Ԣ-8��o��Y�d����2$Vj�^�;e��8-��A��_}�C�ǸQ�G��u�0>�ε-%�����#,��ll�`�i�F��gu�B��:�h|G��R�peQ��( �ip��n�]8�K��K��x'|��t�n{���	la���i�={-�ݏ���o
h�e������dYB0PN��Ǉ=�-3���n�Cq<��n��Ϩ3�Ǒ��q����C0��d�F��0��1�̓��+��pmS��,��Z�k�=MU!���a���?���is�p��\������*�V�9��H���THc��F�S��yH���#�8Ѫp[tQ�`%������$�K@R�V�Z��3����Sګ�.�i��42o�rk ��J(�0Y��9ȅ���*碫�G�:�\�E=��F��F}���THmH�j���6#�i��iTA�afh�,�TR����a�>*���������!�5�����+�p���1���3�̼�n޹�K3�S	@*�����OǷ���w2�k�.�������{��v���VP�,u"��=�5�8���@�~$snԇ�� �J�6�$󕒇0	������<��_�w �и��Hc�*y�j[3�qУU.� �����v9��<�[U�ǹ����J�D�exՖJ+�����ʡ[I���ͨ?Cxm�"H�VG�b�xv���[�瘇b)v���8�+у�e�e"���b��r����5y���	E�m�P5�%�C�����u�bU0����{�q�����^��o���Y�s�� �tE��g#g���B��9:|?��3��,h6��h���V2#���3�o�r�w�rRSs�IeCO@���G�/��ҵ0a�UV�:[?Y߼m�>� S5�wsa�npF*t?g�l-�R��z9����e�6�o(HhW��I(=*�1��^9������B�يpIM<�f�Չ�<i>�y��|7�_Q\tl���#T8�`�����ɽC$ׄC��6VMZ��!���ˉ��*T���W���Sg5k�H
8- !G1�:��/����3��(��kD���2���d�J� ����^J���9��5\*�a@	�T٢�����)��������}�F�� $�/JPԗ�Z??�.���KD�
Nr�ğ�E��I9���.���`j�N\�mM	��b^�G�_u�C�!]Q]����X_.��P愉�� ��RN7f̓�Z1�P��k����׭o���ð0)D��b��:��S!�~�䕿�W�~Zܠ"ϒ�l˙���4k����Fz�\"��8��)�C1z��!�ʇ�(�_ou���,��w���Ņ?�4_�9~툟��:���3���a�@2uN���gNL���2�h�oՈ�20 ��rY�d��M�@94u��OA�)���X��+NRk0Ȝ];�z���S����(��O�|�*�t^�TrFlZ�1+��ފp��W<^-�t����_���"��E�-�ȬY����O'%Å��"�:o�gw���~� �����K�^�Ćt1�S�s�ujm�`��ո4`�#�|��(]�2��%K��A���B���N�7&�X�wi�����-G���]À��7���8�C��"CA��~�l��-�b�e<C���`��%w�ьY��d	�,��߲-c��A��:z_]L+c<�Go��Ƚ"`V�S��5f�1�3�̏VM�v%j�O0�G�w]-`;��=�<:�PŜ�Y<@��A^���%�2�����r�&(XIP)���!�i{�ݏ<�$29* ��.J��<R��~h�8�T�L]*�r��(l}�]�CC��L.G�br&ƭ��	��o�ӄvf�����T��b��¦s�ŉ6� ��ײ����u�Z����}s����8�`dN�n�i�h_}IukN�f�5i��ʇ~Ce���u��Q پc��#�+�.;�s�ο?��j�uĂ��� �uL\]��6Q-���Y�bR��j���v�H똴Ҙ�*�[�P���J�o{S9�d���6����<wD(C�ܶL>�(�I`�������=���8�A\5�>�]�Æ �H/�K��`��ϵ+���0.��L�C�%jv�N��"�T�d����e��:h���Ku%@��N�3'�]7���
2�	�vrQ��^��غ�§�����w�O���9%�5A����9�A�] ��ݯt���8���w>*�+Q<Tk�*܅n@�lE3�0�ޓ�Vt�0Xֈ	�Z	�B�L���G�Aw��CQ����b�(d�~W�hTI��Y��#����h��G���د��/����m�}�$��A���OC�T�+3 Z�h\�×:@���E4XW~&s1��Z:�JA��7u�/�W�k� ����-�	b)d��%��KS��Ɉ�Ho�ŻLxS���6��^�z��A��9.���!��{���ٴ������dKRx'�Z��5fKʥ؏�~�k!�B,�rO`c�t���1"O���r��W��1)#�t�.�^�U�:ˢ���f�S]A~g#L�,�`��`�b^�<� �[u"����q�b�h���
�ns!pO���8�p��Iv>�ɶWSOm,�D�<U���{���f����P�S��dt�؀4E1��Nn��T��AcTM����j�m�-ja6g�i�M��^��!1^v.AC)���7k�#k�ɘ�~���/�;c��kw�Ͷ��:�̩��~��X��h���.N�!p]�S�����1����Δ�_��ɒ"~�=r!�c4� )�g72����C�>�z�}hg����P��nY�.*C��5S㚟DF��֢2Ot��tl�+�ˆ��ŅBD�$�E�'J�ҦR��OQ�ݎUZ��0���L*<$�E̗!�3y�6\��H�F�	��Q�[�VR�pϡ9o�\��R|\%)��.�?���X�c�Wv���%L�9J/����3L�m��x9s�jɈ�M�Hp�R� �a�-3B����x��N@9bH� �V�#�=�)EGS��i��Q�0p���e�R��Ԛ."*�'J��lN�OG�6G݀���q�tV����+њA�+EO�1��qΠ�����ӯ�t�{6���0|&p�rM�b�)v�B�Ӣ� N���{���a��EV�2āZZGS�p5.�z#1a+�w��&NA"ǥ΂]"V�z@��mC�͂{���_�V��~P?Z]����U��eV���9��_������'`���J��29��~B}}�-�k=OVt��Av��A�M��+�ܗ �2�݆���$c�ՋG�vԂ_ӨOv
�3�d�B�P���J�´'���٣��\�>�i�e��+���w���A��5�T?�'A1u�!v��?|����茧�R_�涔e��V1�"S��B��B���<y�3u�j�UՄ�(M>_ �TN�<T���@	�*@x���\��&)���§��SC�(.F�jGƋ���s�o6V�Pk�)�V��?_sN��ϸ�e���OG�^KA�p5��/�ޤ�Ԁ���PW	:ƴ0h������W8)��(��H �z�A�dE҈[z�gp���x؈��0�{͈�C��	�9 �3��g/�K�e�Z`(�;,�$�_$��2
�ZA�&ޤ���Iιk�����K�q���REۆX�2h�3�Y�ԓ�N��)�����l:��X�*��Ӂ�j�	�n�[u�l�#�v!�l�=����~��?�����k�2�JS��Ys�+�KDz&�w��ř5�b�'`2�(|L��l��Xe
]L��b�x���G�S� �����x���e�2��}���o����B��JbB\�ӑl�w�K9�Z���_�;���)���H��.�w�.�F*�����]�tq�c�|�\h��rF���A2��O��	
��C!j�7�4�A����l�j.O�����,Kn��ު#@Y �.�R��
'�4��+������h}�8���W��]tiV,�>7n�TL�������/�d3��s��l,C�u�{~�E�g�M	E��@T,N�u�R��(�5����S����/��7��#]��.2��C�$��W?��a!����l{��A���A��\��q�c�(�t7�[�ëo����q��F���bf$�ٙZz�JX"��n|"Idρpʆ�&ūA�_���-�Y*�ݠ�
W�Ďe4���>}���ж����*a�%?56i��c;Á"-/�H���`ۭ�Uȍ��$L+���O� �ݲ�w.6����-� '4�����rr�ytͤb�֎sw*�����z2M�RA���
w&�"S�H�TD��k� ������g�S������R�JR�z�V�U۵_X�ګ�a��DS	B����3�����"�sX��K���7ݐ^
!���Я�����_^4��n_��/�@����)�n(g���}�~- ���#İ:̿B��{���+�!K�<���L�ODVυ�>=e��x%����qFȠc��;���؄�Ֆ��EL���+Qs��c�ϓ��=�J�͓f�\������/x����О�W���H'!� U���?-9��X����j�Q�M�7�9��mɐч���&�m��*fM�$ZE�z�'��ة˅���S�W������RE�Qp���S�*Qn�x����X$��%yE�����^C�B�f����-ۍޣ|H��σ� gj���!Ь',�;�2͓%OD����.����b�c��o�GH��?O�CV�}��-��Dwdϑɫ�G�w�P���6��d%�伐���<[ܬ��rY�#�'&��/n�[{�Jk�I�4����L�d�1��v� ��ї]��	W{F�A�P��RD�$tD��@v��SI���0���f���6�A�^l����/���&�Fu�@ͿU@���W��Qg�; wF@.�GVǿ���]O��پ��/�vVr�d�Z+�r�Ļ��i(a!,[�d���2��$�x�4�р��k�j�/����Ƴ+tS������'�1�G�Y����m=���5 ��w~��W7���j��3~�8�}�C@�&�"k�z<��<�GΔ�,���= �� @���PFM�M��mR��|ԡ�I��l�[�Vݕ��џS�;a7�H,���wї��T[=H<f�=��c-vZ�N��@Y@Oٮ��%��@�~��EdI]	�Bb�#}6�^@xh�>Q�Q;褬��U�@y�����J���'�����wV
%�;�C��nB���{<��A�-��o�Q�#n*��u�B���eG;�j����yր,�q�y�%'.�`	95H��ૄ9�	6p�%}��,r~�)�B���]J{�B���/V1�!|����VIL�'�8RR����J�-"b�{j[Vy ��5j�1*ú,���0��)m��f.y�����Wa��^^��E�l�_DW�EHl�46t�2 q-'�FR�g9�d�
`�Ͱs��ȱ�~FX�r��G�4�$�^^M/#}�	�l�a�j���}���y��I��g�gT�y<��P��u�t�,�򺯚�G&]��O�0�R֩]��dR�v�)p�&F�N*�����Ǝ�*����R�-���ur�1VU��@��E�mb)yzz�\�抦L�mIn)�3*\%��e�+���z~9vF�2D�w�N� a����W%�$#2-��Jy�8�f�u�J���1���F��}	���0�B�;�m��q�
gh������ι
��~���X�~}t�����$�90�z��-�7�7��Ū�y�oeî�*I���K�߁ї�/u΃wG'�ޏn�3:�Q�_lB�Rw�w����
���+�%�
}��X }ٶ��K���#$E�b΂Ȩ�R��5!��"������ �g�M�gvΗ:}z9J.2�諡aƢ.���(�2�7��/fPM}qvB�g7	|O�Ѡ��n�_Y�2���V'����,u�:�l��O`�6qR����Y�!ê��Ôbΰ�S5�/f���������l���\��\;/Ǉ�2���
_:~��+\�ϫ.��G��^M����kzj0��G�A�t��˦����+����_Pt�!��<w#=��N"5#�������ꝉR������@���k` �G��c��蚯-H������O���)w���/�#�.�#qL�uA��k�ThB�R����E�,�	|�u)�z2V�oQ#N:�D�u���|;O#h�wä[��9/��m��Iio���5��=5*����,ӀW���J �vg69ݪQI�aPY4#rd@)�ג	�g����"%$n�����OŶ�6 4��g%ڝ��H�
5�:r��i6]L��$�~@�|�0�����j`���y.��wּy��C��@�G��Ǫ/sw�>�����d/��8�z�A@�	*b(x����5ސi<e�����۸��_m����t�<ɘ=����ђN���yGҲյV&?�7��u"�,�����VWFt�G	Q���3�;�i�W�u�(�
g���V�An�E��T�!W\viR`�Q9=��%�8������j�#>E�@�����d{��zq:�qꮐ�G��^�+d�R��]{c��`�&Kn��Gm"z�'���z8j�Ӆ�#�l#�컄fXw$m��-.YY�Cˡ�s�un�G�Ǣ�V��XrSii�h��qh-���PAN��-6�5}0��Ǫ��ᩭ�����v�)��W��Z�	�.�t�O��i�	̡ʍֲ!�Pmw�0@�D{�/T�S:JW<⎻Ot��=|�;������\T�䃝L�'���n�7���Y��5u;�t)Κ�ԅO�	#C����,s�o���z��_O"k�ŜI���s���."Jf�=�zW'`-Q����*e�͌��������TA"۞�R�l&��i"�7�n��lOJ���F���↢�D�G�dBہ�hwO���g	?Lx*�|G��x1�@0�aV�H�r�s��)��F��jtfc=T��i/��,��ޭ$O��ׇ�uV����+W����j�oi��{��˰��xx�L�_�d�T��
`�g]I��(�D�n}-eh��C��d�-Z��!�c�)��j=��x{��ɕ���B5kh�Q�pDp,��$8{3Hί�I�-"��Ӓ�ňÁw����/@A/a�G?���$�N���Np�}�&�:"*$D3]����]
6�tٚ��/"�7�l,a�zH�)�-����V�AW�+՗L�*��'���!��Vr���D�_��f�[�$b�;�9Ҟ������7w\=��U{[+��I�pw��#�F��'(��r�9C�:'��M�=��"���j3����8*�o\9�&n�s͚��l���b��@�Ǌ�b��;�\_������{Y����n&��ط���4�vzԔ�<Wu���HM-b�M	[�ހ4&t�n�|�u���vh%HM`#�_�»���$4Iҧ�V6��b�*�EaM�"�V
;�v�����<�XK�y%B�m-(��"�ۃ
�STo�P�4���Lz��4
/u8xZ'��rX�7�L¦��nj����z֠2�*����SCO���٩fA�����+ls�n�T�JoՉg�N���G�M�6j8��H��ݽs�w�����H�\�	�u��N�<�}z�k�^�k`�K�t����
�����r',Ѷ�>�G���n��&�L?e)�Ї�����k��4�i�
���˸s�l��Ԫo�O�e��X<})+"�V��e¸9J5i4�����*r�w�5���)�2�r��UG�3%-(��M�w2��8\s�s�U�^�@R -N�z��,�K}��z��q�ӓ��X�M%t١��?�����1�@�X��K}��no���<O��^hY��SD���:�v�!��C{�UGK���X.3�	���_�C�{�k�^ B�e	��Z5e�M��T��DL)�[4'������J ?�ȡX�M�a��e�x���X)z6g7���Tj�lyO�5�V�5�Q*�F�"���fə��4t�� ����p�l�6
������3=�{���s�
/�g"ӗ�q�u��.K�~�( >-�7�o6�$��z���c�_r��n����P�EE}�}3�ܑa]�N>{���K�F�~�+z ��+�9��t�6{b�$Y���u�vc�'��T�FI�z[YC���B�$ЕvBgzG�9�g�'\�t:DlQX���!oJ�s��A���j�4�������Hª�a�);����s5�{cž$����+`�;T��)M��J#�ܥ!�]g/���m��H.��I�KmLW��.��$$i��@1:��!�2�_�~��/�7��Yۙă��'Rl_�< Q�ێm(N8�w��x�Gv�q��8���ʹ�Bv�J��i���9g%�[�bs�ː���ԭ7���3�����R-�(߲^�'����m���ge�Gmj-�o����H��nߑPDůҴ]X���Vz;؆RM����]���+¡���kp�D��B��h�	L�b j��R�7$�g��"�%�R���=����N�7f?��8
�9c���v�f"`�]ф���ej�����7��CԵm�#������L<)�,�׹I�n�,,�eS��v��?�XG�h5�,�G6>��#�$���Vw�Ik`�(���u��U�G� �mj�e�Q�R2lX_��_�*��Bl"�B6�Z�� �^��[A���.�zϠ6�\�ӟ 
Hcg&���&��ץŲ2[e�{/5r�x�1������V"<�o���A���4p��N;��� �AIUX�[�}�	d�N�>k+�QF� ��9lH���v��ҏ��*�
�ǖ����ևv<�t��ֵ��W\� i5�<��"�<�&������E�q'��z�J�8�ͤw�[̜e��zӼ@*kߩo~AE�ou�/�s�(�P��㐀����̪ΩQ?�������o���eF
�؋�=����7��8μ�IU&�I�#m�+6PU��VX����r�</�Xg��{���]G\��Y���{����d����GeJ{�f�<I����$(6H:�0Eh���x�8�},���GU�[��-,�fa��%��� �y-+Y���$'"W�K�K���ȶ�l��Y�]맟*��Ǎ�.�t�5؃���u��B���PﯽaU��/����RG�v��~�$b}�$,��2s�����x	�vt��!�����
T'��7���9��?)64��.	Pӥ�M�87�-��8Z�#ش8��x��U�
]��y?�c�k�¡i@�Տ%�|L<�%��79��v6���ˢT����^�7�!;��ʘ�g[�h���B�^�8��NC�V͊��{WE� }mcP�?WG9�a�0���Aj�M�!�	5=�X�s;jkf�4�]�ʋ��G��U/�X$��#����/�V�i��b!����O�L+�$�?W�Yc�k�?
~����V�]S����]t8�3��̮���= �	�� �˵��q�K�W
&���N�<�ujN�_�Ǭ����}tcA}<�,R�sq��� i���v��M�0XW7��ܵ&��+�3RM��5~���JK�"RB�������|U�)\}���,c�J��@����c�v�/n2����r0j�
5t�X�f�'dg�3=!��35N۬"�	3�.EC��ha��&���gʳB�e��'Fx�� ���+ۿ�yHR�Ζy��%x�v~��;u���Sxh���|����_���R��6;�$,�K��:e�Pק���:M�<���_2��E����4ΧT���/���h�Ev�{��bH:"��(+YΟ�N��͙ X����_u�a�����5��a�B9���-��=ku��FI��$E�z�I����l���3.0�&��6�>0#n� W�,�,�a�=�f�V��P�):CZhh���âw�Z��-2�'�W�ZI�X���dݜא�}���GZ�4
!HA�ל�R8�O���Ҙ�]��ɞ����u��RJ|\��ʖ������0��D�Ʃ-#¼%,u0��WL�OAnzHo(��v$G�J}i�1�#���������5�@N=D��:Ѝ%�����5h�s�&�ЃnMIA�Cu	��$ձ�iI����e?�sO
�%�^��=&>jS-��3i��Ed��?��e. �B]�3�4�v����6�h�$�O9�9�j��A�sdH(�[93�명(RKe��a�<Ԉ]{ ^p��3Zbiy�1�#H�C��W_n��Xw��"xXA�j�F��S�@�[`i}T�9z�ˮU��J�Qs4���JR��������n�<UN'���W0*��&h��w�V�Qb�������B(��3�S�^��x��ϒ����q�[^2�0�����i�
�Z=4,d��r��^��i-/y�F*r�h&bH*Y��F֢w8M�r�M�`�.[��>�%8lk��"�E�Qǽ�����u�Mb�\ÄM�$�>��v:�i���Q�n��������8���a�HY��v�0���B_�Xle�XDm�� �W�Դ���8����ֱ��-"4��j�E j��C�b��%�?�.C����b/=<wȈ����!9�H�&��2��\@� �� � vI^7H���������!�Q��H�FeKY�~7Vz�iq��$.��U�6�J��k��� ;�ܚ����ȺM~*�5a�uI��-��$c�z�F/��9U�G�l�BWng�jEgP�8m��9���^�&��Z%ݪf�S/\	dh9�F_�w���1זNX�]O���E��7���:����0V4�d:J�u
�K�pK>WK m,ԯO�qs��V�b���WL�*�H<�\�Q��ݤ��!$��R���9*�^[�-ǫa�s�{6O����Ĉ�+e:�_����Mh��ɐ*���&԰/�W�Y`�br�`�-�����3��� J~��(N-	64�|SO�M!�g��F���[V��;c�Β�1�_��]�$2#-�!�h��o�cG��owD�픘W�d������R�����r�;�*T��Շ2�0�|\O��:��Q@�� Xq��g�a-&�f�k?�C�~9�Q�H�x�`���2�����mf�8���U�&n���6�i�\+�#�"�%ZP��sc� ����Q�Y��x��t��[Egv(��m��=k�9ۮ.��>�}��E��� _ٵ;N�Z6_1 :�&֮2�1��K�JlLz����*��IܩDY�gd�0/�z��"s�g �l΍��|yx.j!��!���7�)�dXƆO�ct���������SW�b�ɩk�b�r6&�dauo7rW��(��8��	%͞K�r��;b����$�)C�<h�i�!�m��r��|��5� �pX�O���٩�D*�������|�(�C�0��D>�D�����iSy�r�G�R��BrV���ʋ56�LY��3U����nf��Ք]bb�/;cj �������\*ZEVM��+�w<�;�B��-#R��p�5]����d��@u��>�o��>���Ov�G{r!�8E����������^'me����d�EV�~O�϶ճ�� ����O�������yjf�@� >��� i�-
�I�B��T���~7+����4~�C����s�ptr��n���%}"����X�E=��RB�C��[���y�ζ?m�4�P��=,�WubK�6�!�?z�%�L�Z_��2���&f6��Q�F�:�f��gV���c���ϫt*%-E��;�ROq�䊥ʲ�qv0ԛ�3"� �%(@��k�^".�Z���'}��[�#��UIɃY~W5�jK*,�p���#�'����[�&�z��=��wB{�6�͢�sκhc<�(n�|^3�B�\)-�#4�U�Q�=e��.�n���h�`�^��Oa��f@�:n����n6>@�>Q���� �K�<I�mk� �a�{�r�@�7�l�*+@��*/��,ހ��:4<k���>T�
^��|v��OvQ�K[R � �We��A>��ަ��9�G=F#P���H�[K
�-=�㤕� �9)��#d�����ͺ�SL��������"x�������NI.���죫�a����U�X��Ν1��������*I�J��ms��V?�`շ;:E,''kn3O���*�q��Iz����@��D��bTi�nɿT�1�^X=��/pΆC��"�I�L�b��!�����W?���P�1a�f��F'H��Ψc�C�4�e�;y��i�Տ�U�V
�J��J{�Nl����4g�-�	X�y��/e�V��G�-F!��=�	����\�.x���{��ѲW���Z$��z>}�&��,F}N�c�ya���i}>���[���eM8�
ղ/�'P���X�}
��2�����@T�
�M`��!V���Fa�%T]_�걞2@I�{qc��A#s"}O��g���
�e�)�w�B�|¸��"P����z�1�1Q���ď�E�:��<4�����ZE�$E�-���dp(r	Ov�ا���BڍS*�Ć�7������±8nt��s{G�?`��0�0���c��l��.���^��#t�=q�*c�a$�ˮ)b������<e-L[�7z>�#7�$��?�/qw�W S�����X���a��"d� ������5��eԔ�,�˜��ó�j������J�uzH�/5���y?a,�eh��+�.Wn�n.�`����������+Q�_�h_./�M�l5��3c�[�#��a-�Jz�٫�Q;�ԁ@�NE�W�//�	��@P�)�B���%D��T�3��E�)|�U^6kNS��Xt���4���zً'( �V��ާ�#�Ʉ�h$�r��W��j�K���U��D��w�*� �RʹAq2*C����I3��R2�`Y�8;�ɚ��dL��?=��J(j���6��g{U��LcL(����en���.>�*��8�+x�DQ�-~�nS��f���� ]*r�T	0��|iN�.4�s���4�m����^�5�ja��K>�4]-��"o�;<;�ID[���U�߽�I�o�^�A$tk�� zo��������������(\���]���I?x��������m����ЮQ�����:xO-�����!_H��a��կ���;3����"f����ix�WF���~��j���r���#'�EĀź����G
%�3�� iD,�������K����ݝº~���b#n�����U���dmF��P��]ɧ �4v��=*�~f{�Tټ|^��+�w�"�/�?�8�c]f�p}�5��Ub�����FV#�\��ni��m����WP���N����
�scf�P'#�_h�t�t##�O2ru�fW�vq���jZ�X8B"�0723^���UA0L&�	�c>i��$SC�R�H��Йo���@�s�N�5��~��(��b����Z��,���g�잱�lY����1���`
D��3��<ȁe�gm�7�+J&�?������ٸ�7ئm��OR�i2�k����d��Lհ<�тS?Ԛ?KtH�X��a�s���fR������V��S1� s��U�b�%���1p�Ȭ� �*�� �	y�Å���0�HD�r�����-���� ��2�I
�eK6�D�hr��R�V��=��^ E�?�.�q��^+i����-hb!-�|d�,����Ve���n�A�Q�\4"p
����z��-�`,x���J+en���t�D��X�����٭4�\����a�(�4������6�؞h�v��^q�o�"pP�֔9;��'���3Y:L��q�V��'fk��	�fnZ{��r���� pL�(��_�G����^~�y%gx���l�-3�l"�&��t���� q����u���Y���
ҭ9�-���(;Q��J�\��>�¸��tQX�R�.�O.�I7B' �
��[���e���D����hK�7ք�����-�;�YD�p�㻟����"Q
�hRN��E�����}YR�֫��5�������--�9�6��ک�k?^���U2Z�y�{	�����H�?Ce�v�3��-�}e�^��V�k��~>tZ��J첞~� *���7
1H�'y�s�j���dq�}���r�A��]�oy��)n��m:7�M��H�;jZ@Jc�n��v��뗸eue4I=�G�O�r�uD���������ݯ�e�������Q��`�~��Ȭi�gѕ���F�jo2����˕�B����8�:�#\��{���O�6�?��0&ڮ7�P�hEZV/��공���X���#ӏ3���&�����E5'N*{��ʍe�bUaj�$�x���Eu&�o�^�.��oڱ��gG�����^��|Vx��cM��I�L�2s�N*C}�U�"��F�\-N��d+A�Ip�,�t���`_��6�"�����c�S}��$��C�4�����3'�0����ŽX\��9ˤs�������[�^od9$�)�8��D����Q������w�P�"��I�j��rK����c��u�vc�n�c'k���Tl����zև��O���{�%������ I�#+�v��ו8fJ�y�Hɳ,?,�!nS���9���5��"�z�A#�ظ|��]u�z@?�2M(��h��Y@��U'z����X���H娻ٓI���c�.�fN�>��Sn�J.Ϫ�o\����Aw���QT�_�?�؊�j�{`���fTڠ��{��_�=�3m�J�Ɏ:�eO��� ��K�����,ԥsN�ޏ8��s�X��v�WY���vic�.H��2#��0w�LC�Fi��0J2�a_P}#8����	H��l#��^E��6_e@�l�Jcӛ�{��=��#P� a����Mo:����ueu�#�U�"�ٜ�?YaGQ�}ʎՀAS�����G�i������H�6�6<�J�~���3�P6�W1'�=G�o�N��x��?= ���~+r��"5�	�6[�vMgd�g���Y���7ӧ��Rb�ڧ�0k��n�
|Q�5��Q�����|�k����1�_d�"c�@��WN�I�v>i��(Yt
��P;To[��ߩL��^o�xo�{n,�5��kn:m ����Ǻ[���S��_�l�O.ѝ�����ٙ�Щ��#��u�HB9�;����o�gA��a#���ܝ9'L�
m�RE���D���D"�*.����16��-|Nc��Z���ڶ0��$[�I�㕾U,�u��=Br�x)^&"�WN��6?dT�yahx�IE���'`U�(t�|I�a�}"��sN�AEDP��>-��0>��p"B�e��H@Ǘi�O�hf����M�t�}�R��}���K��:�j��6{�f�����ʢ6|�埼�|���g�\@ʨ�ɪ*�����*A�����S�ۥ�'�����j'ȕ,s8��>m���c7��R�k�b�fԍ�q�c)��M��/}?��7
�<��Z�	k����Á�C�8�w:���Q�eY& M��?�䭠�pr�FD�6�N�i�Z��+����
�]I��5�-�/yT��L���3޸�Ҭu3�-��v��}`Z��士�NP�զ�H��z�:�Ot ��a�x�K�^]��0���K:��=�:T��$��L���D�`������k��C���܄L��q��#��	��<Q�86p�N�D?O�H|��x.&P{�/X�>�Q������}w	�6N�(=�ٸ��@��w��}Y;�j�����B7���sg-Mi�T�v6w	7Ŝ� �s���p��{%�mye�I5R�qS!b�)��|6P�(�c��:ع0DJ#�b�k�|b{��/��&&��f��\|btL�%�a>��^ѝ��;L/]�44t$b�J<���'�榑��Ci�7�c�0�"�Y����ttcH���n݆y!V�ZD�w��m�A2�K*U�B���v3sq�[(��w˛V򽃎sT#���<|�[�zF�j��!��|��Fc�������9�BG4R�9�kx�{d. π����IpA�n�
 ���Q�:z�ְ���c�B�<��cX���:�� Codo � ����kq��#+�1d~I�o�air�(�}`ۤgȇ�ٌ��^x��)	��\#v�u��PR��GQ�nN�H��u���A�<I�Tt$��3�;��}+Jja�͛���zs�d;׫Z�*:H2L��^F����t�kco�U/8���L߳\��u[��MKׅe��;$��r}��Q�N4��g|C�=�]b1`(�4��o�i-�=O�b��e&�Q��"��
�h�tA @v�1��R��Ī��щ̱�5a�FO��ynD�"�!L�;^re�R�0!.���8\�͢�?�zc#��f+0n��MTkU� !�'�P�MfP�V��F]1i`V̰���W�d�!	on�lU�Y_)R!2~�W�	�@`�Ku���%!���KnEý@#(�A����
b3���M
Y�8Ǡ��C8)�y��(1�X�r�����݈��)|��cȯ- &�4�Y�f'v�j1 )a��ξ�~q1,<"	9�~����砪���!�z�5F�Ҁ�׹��4�/�i�qվ��z�k��6���C-ހ&��G:�]:~nA��"�"��}�J���p\N͐�ɭx�M]ñ���tU���L�`�Ն��}2Ce��?�kĽ�&������ڄ���g��vp�Msu� ��EҗՇ;ۧH��S_�ߏ���F��rƘ�c䙌-��A��o�r�����ɆU��";*���G/�u�U�j�T��DՋ�j]-� �|��\���}Vq�ݎ)��4���G-�*���Q��@C|�@i��E�i��ѫǽ_�|�3H�^�oBz�*�-���S4�];K��	��K?F1�K�AhXZ0��~�J��G����|���8���V�Ȃ�,�
O$=<];����O�� ���t �0�
��C��]=���L�|U��J6���,sj͆&�ǖ�|��g���9��b*�X@�6!][R�����-���{�;6
�DE�5�L鸶G6�>D��&����u�ˌx`�X�s�F۞Cۄ���ꣶ{I�9Ȋ���pMw['��%�h�#O�3������nz��� �#�+T*�7w ��r_���<v����VC�E��
�x2m/ޗ{d402p�}�aI�:�o��=�^,� �<f�o1��<2܊
9�L�����{#�ӶBV�4�!z�W^�������h�=%��Z�00wrmL�uµiik�$-��]?"k��ӗ�@�DN`�˝"r��9ذ}i��N��)�dj��;�u�O6�-��߁�,|T"u�b�3�}+��9)����EـE�Z�Os>g�GX|�k=�M���c��loI��5�R;&O�[LG$T�(��پ���o�(���s�U:\��`��a<�'�"
���	;�	���e�Á�ed�����mv)�*�%�J�B�c.l�T�k:�� CR7p���������$�/u��2�ג��Pk���g�n}����x5��EҿԽ?�6FS�8���b�nP�$���,<`��	����ѯc0R�W�+�!�Y�:�Øi�n~`��C���L�F`�c��$��/v�
gѭ/��S�e��2�����Uz�Ng�߼����MX9���^�ET��M�'p�T;�Kq)��j��.���{jl�<-j�����$Rc�
��D����9 �0�����Z=�B�0-�p����FK���b��/͢M��S�#��0̯3ҿ&(�ϸDfTw>Cpe�R�̳(�#T]��H��Jhf�(��|)�r��4��h'��Y��e� ̲/�|^hg�W�`W,h��K�L�Kʀ��^�i!�TI>�Q�TQۇo��(�������m�Pk�sTVF{�K�M��W���ꐽ�K���,;�� ;�PS��p��dϰ�.�g�C.I�k/b�5�y8��n��<�������ʫ��l����l�]�V���Vt�V듏�H���9q�#cQ��;4e�P:fi=��!V+��˽y����խ�:^ё�տz��x�
�u��J�=D����m$��'�JSM�z+�a���ڂ��hҺ\��K흧�>N�	��*K��Q?�ـ#�u�Ǜ��8��+|A�����Z�2/^����)G��x-%Rz�S�2��*-\X&Qh����i�7���D�-�J70K�탆_�T��-������V��Q�U?�+�8�����l��g�1��/0��X���7��~�`sج��˫�t�d�0���w��Bb8,xw���
�~��q���v�G�C4�	�,!?I���T�u1aP^k��9k�j�ʀ��Q<�i��"�.?�7ϒ�<��<�?~ɻ:����;���d��jY�B~�b���6��Z�N����!��w�-w�#��6o�p�{�< K�T�YF�Uq*��l׌˂9l��������� '��*R��*bq��g�y�a�p�Id���p��!�)H��8 �nF�Q�wK�v�E��+i^}�!N�WG��� �Y����T�7��
�-�Q�8�S�<�$����%�,� ��KIx�v�ev�́��1D��u+ÎCo��]��&���������E�.���8j����*�1�nA
�cO�,4ut��~aүgt�L�3��%ty0ʝY�f-�}B�����,M��O��®Ҥ*�>v��s�8ӎ�Ή7�B�.@ ,P$�QF���.�k��V��-����,7�VKr���I��Ap;}<����- ( �����豋���a�(����i� zbK e�������mg�b�t�	���^�)����^uw,�O`_�M,dyz������+�$��}��5�_�VūW����І3�mds�DZ��nϱ�����5�@���d���*��H�Ũv���!����/�c �&�Is��q�$��2�fڀ�ؐ}g�q-E�����Y�b�d�y���=UL:�s`���E��L�l�yY�;κ��n^RWqs���Tt-�=�֪��]�C�t��2�lf�[�E�U��&�SkJ?��xk�Eh�g�'��Zb�5R�V�h<߉h<g7�WX{&�n�\�!�_�hFN/�@��!YW{�O	u����~�b"�`��5�z�Pj�܏![�(������ӴM1ܴ�q~F�!��;�~KJ��y;q=/@�c��P,�C�tj���c����ׅ��T3�T��OvG��D�Hm?'��x��C_��̴���7�d����01!�[�+�е7���ԅ�1&B�o�N�Ϭx���t�>G>�A��m�xdC�-~у
��H)�2�-g1��}�#�Z�և��w,��f�� \�CF�k�.j���?��ǩ0�c!B�F��(����l��l�n��ߋ���:c����m���AJ��7~��ا�g:ӼB6�}A.�q�=��+�]�t���뜭U8�����ɀ�����
�o��݄�9��l�l�a����O��b��8X�#EWo $\�����`��$	sb��a���!���π����nz��:��o?�.T�Tbv�v*��ŲM��f?�EO��ڍ�>�3=�:j�p�������� ����{�Ǐ�ue_�J"S���.E���(�!D��ԇ�!�Ν�U��19pǊ���BMEy�iFu�{�EL1�4)�[��7t�t�h�F��[��S���5W��Wu5��+�Ը&��S��a)�
U���*'��M�M��_I�h�{�a�!8��WzxT̡����F������˭���bnA]~G;ow�щ�]w��Oe�k�i�]�
aC���=�e\�k�/`��T���V����0QR��n��[g�O��0��V[�tA�X���p�7������8��Y{�!؂!��}d&͠��6UH�\)���p�mz�J� ��L�+E?Z\_t��YE�u�t,����M�Z���i�$v���eh��6����竊���ۣ��Q	��k�$Dl&c����	��B���{\Ƒ�$Z���p*G���_Y+q��
;���b�j6�n��NLD��A�Æ����uNa����l|��8�L����v����������Rt��ǅ1|-�������I�l��G9���̿�j�SD���K%uPx�mL�ds�.�>T|O��8B���Q�Ԩ���&i��VK�ٺ�� �.6�*F<��2��a�1�1�~�{Ѿݑ7� �x�d�D��ڦ�8�.^#�Vkq����9��w#������@g���U,
Ń�_�k��L��^0*5��Ҷ&���-�s����6g3���9��]�W'2�/</���1f�!{�n��C�#>2�}��npW��U:��ޯ�Q�@�%��&œK�Ƽ��Zg44��f���9�Y�0��ǚ���Zw�(yr�����w��~��[D�v�2�Bw�@�QMc��'	�E�������ڀ��jF����
�p�/0KoW �f�bIbp��Q�Cî4K,�o'CIy,���Aw���41� ��+����.{��%���$��K��_q�穗_����=��3[5��u%6�xQ@�N6um�m��K��-6?~����E�}z��0�QX�,�����MwѴ�f@%��L��%l�dޟS�:6����`��H��p5E�O�O����vN�4In�K6Hs+�mf(J�"�{��Z}�Z��
G����ɥ��薟�<�hu\ܻn�$	i��q����^�x"��-]���h�k|Q��{�{��pQ���}K6�> (���:�v�Q#��&�_<�sp䬻��M�J��;��0F���K���\�U k���]R��J�n_/G��t�C}V�W�M�B�p�!�����=�&ȗf�_S~!)�5:��n�7�2<�q����)�L�E&�?����Q�p�e��K�^�r˓T~�𞽛���f�7St��&���L�S?���/��!��=�Ocz�K-����_N�o4��w��� �����jE���/�:��B�zM�����!�o�Bw. ����4�c��l�E��
\��Z��x@��{QMu���|��g�^	lG��	��W���ۥ������
;�cLbc�S��΂`��A>99`�f�˲^�p��K�p!�?y������V�re?+J56���O�����GOo�9� �f+lN�#�$�0��3sP�S��n�kۓ1��^��� �!�x{�6�x-��qE�ďl�W�����1�tr�r�K8R���������G���&�S�8sꓒ3ӯk��<�L�z���}���d�^2*��K��[Yio�lW�.#/L;�슆����7�A�*8}�>���-뷫�}ZNּ��Q���J���F>�)�xh:���gN��`��g YVºZ��-��U��E��
��$;�yd�끹6�4���+�Y:~�02�^�Y�ZhWVq;�$o��U0!-�q�9�,����-��&�_/�*T�[�7#P4k�O����4�(Q����FYtd&��ܙm�B�bhR`�z��x�u�t�]0�Vn�.E�D9����%9X�`Νf���'�9e�J�h��)��XC׋�	�1BEU�ȇyk
6�Y��ɨ*��d;8�L�ib�s���dx�Џ��@N�5D�P�PyE�C1���B�dQ"A}@ ����	,��t��B�Q79WV~'����(��i#��_�u�B��U(Vs��z
��N�Z�q���օa�M%o��e>P�ǅ�t����]�wk�zV�rp�͆ ��]t�!&��"p�k"QG~�Le9��ŹGK~*М~U/�v1�� 	n�
£�@b��⾗�y�-poh%q�48���|�9>�S}�e�^+�|-2b-��A�e�,M�!""�:��6As(b�{�
\�D$I�ɮ�JU������il�%�����d��$l}�mS�8飅��M�)-���؊�}����Z�M�8r�_�6y[�ZZB��d
[���N�#
-X�|U��_�澗n�o�.�{�l;͘�ZU���2M?Ú��Oފ<fyU�F��,�����}���_���?̜-�笢/���i��z�ve��wu<� ǎV��y���MӘVOo h����X�s[���DI͋�;%�Q���Q�
o �e��y̓�� �]��ƿ�@k�j"�^���:�lW䯱�ѡѽ���*
����C�=̲�c��!������d�4/DPXI�xU�cm�����(ҁͩ����B �.����e^�2��a�G��tuV�M|���N�7�O�~yWuON%�����9Й~�N��i��1)�s)����PN^t-����&�g��ΡF���0?�L��p
4������0 �-��#��5�����#�N]�ZA	AQ������R6�O�Ћ��nq�P�H�"�`��O岈�Ñ�(�YHTnj�Ju9!\�7�{�j�cB�Hzrt9Zi�.��q���4�������W���I��R�BiG��򞬀F~���������%&��� �k��0@��<ag���3,��"Y��D�2��u�����a�Bo������XC*B:��ӏ�DH(�)U3�mUk�:3f\�cFT7�KA���@J_���ؚ���Ԇ��5���o�ME��%ܒS�_<8����vl>��䙋��77}���=��e_���o�W�}HIH*���-W�]lp�}��Ώ��wY�m�ɲ`�=�bM�q��[`8Z������L�d��Bv[���h0Ϙ����1�}Z�3��^q��r�"@JP:���W���K:'ɾ�ǣ�5�j�sިUR��5G�Y���.���]5���C�m)�s<@Wiը7�%_lk��=WC���'X��f�t��ߏj�N��f�e�!R/��&�ST�W�$S����w��܈r�q��6��c0n/N�7�M�,yzq<_+?�Db�'>���e`��b%�R2H#x;�b�f���e����O88��5'���K�+:��{�|�c�~�!��n?�K:U�Vri�d�!'n��H����q����,��Q2b��t-�����Q#�0m�%�ph=�p����D�.��ìXf��Ԇ�H�*�n��U^b桵�D�p��Ĩ^jEn	���7p����$�X���@s��L qJ@�.�������Ka�]��ʍ�*o������<���)��>줿}Q�? 5����%��ME���sA��� Fi��*m�j�D=�<�)�t��"9D�)���:��F�D��w.V�غa!J�)e��[��z���o�� �ð,�	:�'�t��+��hT뼥2���Wc�Ĝqu��r�;1�1��ݍO���&lg��e�,����v���hO�`��s>��k=��H�vM�7�� H��m[��k�r�Xb*�m��Fg 0�ܿF���3R�#{'v)�8C����Z�{r��G-�I�ȯm�zZ���tyGs�˦m�T��)+��I\W��ovg�Y�{:Y�� ��6x*�Ъ�a�qz�"���ꈤ\&�� *�m���sv�N�.�M�]���Q�ل#�8"������|�}���1�jz҂A3}��!���⑌��GM���:��k����e�ևOQ*��k��%��=��rByOn���#�D8���x���Ā5e���Aq0�f��5�Z����$�s�����ɍ�;�`I�ˣ��Օ������ώ��&��1�w˅�I�y���g�(�0�wNLߘ$*����R� $��9���[gߋ�F�62:M�HtET�
ø���M�G�]*\S�p]����C��^�]kl�c��J��ѐ�c�Vd���DQjU&��������3ܜ�YC�kQk�(Wj4~�%���k���y
<�h%�Q��/��ȹo
x�A�y��x�N��;��(�.H,��ޱc��)�[g٬ޝ<F(Ƒ>� �-�sSޓ���������e~�˹��f��;6�q혤 �k�_C�\��1Žz��-�;�5H�'����*�z����?�8Wff��<X�>]��
M�JΫ�{�3R�Փ.x){M8ٸ}B@&�1C�~o!�t��ʣ�7+N[1��u.��L�|��m�-/�.���d���*�l�_¿8�ç��@��g�HN���cL���ӹ����U�/�\�zP:�>r�;� -u�����p�=P���4��ʭ���eF�,;����|ѦwD�)�x2nsY*'��=nꙗ�7-��,/+΂�W�{ ���5��C����l���w�<K�Z�����m��L�3�( �����s�a��;�x&�#�]9�qmhx|�Ͳ�]Q tKu�����6^fj�� b��AП�8:YvUQL�3@W^���*U$�z_�PAע�┷B���P;�l�d��9��u�eܼe�I{���w�B��213�zX������p#$���wfSk1vV0�5�Zg�nv��ұ=�ε���_8S�������H�類���S�.XIO?���5����R+���n3�#H��� ��1�sY�p��I:-	0�J����P�,�?����� �خ�)9��HF?u�}'�te��e�{�|4r��`�k�F-[ tHW���A�!�)8�@�,�;C�xV۶:�ͱ������gl	����u� a���|J�'���貈r&8-��6��@"��c�a,�q�F�PP�r8��E�l�W�eSd�%�e��O��z�F��E]eYf~߼�J�l�Ř�]Z�IR4۝RM`��2ታ�P;>�U$y<�%����<������+n��zi�l0л�R:�掛QSjG���~*7��{ F�oښֽ<���h�ucZz8����yK��%�mP��e�awa�N�[�8�pT-�ϋ�=��v���~�I�H���+}pj{��z����X^ӉG�����DvG�M��7����O+t~ڼ�iIS�+  �2��n���je'g�۱���Z����TC]zf��n9o���	w�r~͍)ؑ�s��?i[��fӳ�lI�~��O3�H�����9 �?�Uj����mB4�
.Y7��#C�.e2E��Q3�X0ɫ�RW�0/���[<�v�'|^ҫi�*hD?$[�|��@��^�S��3��׻!@�k�W��gb'�NV�������9����2�Ss4�F+�	�[9���TV:	���s�<@����wj��SL���"5t�3.:32Ð��C� r,�t� 	I��D�o��K����UF^�0��ƀ�\L���=3�"��Q�{��<�w�sz�%CWEꖗd�]{!b{JK��>�go�'xT�I"��ɯ�d��2�#���ן�X�TY�Y�>+oЂ����{_y�:��}���z��o�� 6��)�p��h�9�N�Ln�� ��|-2�ؽ��4J�!b)��������z$���C�P�5���y�P-�W��\���2�G9wd�y40k��g���t��$q<veM{e<�N�(�	����$ ��p���;�󥰜Z��t3�Q�~g���?CD-mn#����)�.����ĭ���k�Ȱ��$靱=J�e*�����4;1���N6�	��Ih ��ߛ1��G����gR����3b0��T��`w�����d�CO<��E5n�l�h`�&lr{�/���$����ycSq��[�]���}�gΗ��y��5����¢!����i�T�_�g�	t��[}HtCk0�;�I��B�c��W</f�	F�L1�(J��+��$�*��Sl�:�\����%����l���AK^��?�y��\-�37��V�"ݱ,pQb�t�>�XlY��hTJ�7N<�-�d�3�poք�33Ԕ��O�R�ȹ��B�,^R�#
�^�%� -z6��c�GTX�]�r�cg�ȩ�R��B�7"��H�ceFт�{6N-��@Ν6��VG0_��b�DN���C����%b���uT���m�zp,Ɯ�v�D]1�����px�P�!  ���x6�FF�W�Y�V�x1W&�Q�	,"�2��;4�H��vP-�
E�߂F	[6�^�"f���_-��E_��{nX�ҥl��~ ](��ړ��jl\�.�ˀ�����D"�{�{
�ل���$�R�6�#�f�f�k'z�}�#.|������B�ʯ����$�v5ף\{!ؑ�Y��x瀮��^�Iϸ�C�!��q�q2P3�Wqǧ��[��H��a��#g	� ��C�`=X]�C�|ꔹAe�~zR:�E��߂׵8�����QP)����~0��h������k;��!�g�)�LTdi!�9R���.�s�"ϝ��2��ⲹ��l�O*���I����GΤ��.H�Yi6��hT��rq�IyӒ�t���I�03[Rj�o$�KG��K=�����P��w
 ��+J���� gy��+��P(�P�)M.J/F���}��qݤz��ξ26L����M���y[I�Mm� ��́��j:"�x��bl�$�-g�؁!��tl宲�`��=���V��m���cU?��[�N�����,}E5g��<L��F����.�O��$�ϒ�I�[������t�4"�K���i��!�J��%%R�f�8���/uB�H��nzD�� �@��������E:�;Ֆ���9�a���45��T��/aL�o��n
��!R�2�$��|I��c��	_���׳�g���7CJ��킆��?����K����Pgt���^���
VD���PZ�{<y}rr3�*5�,��T]�`�j�PوtR<6��"���q*5�y�*�TX�L�~z:�7��'����<�&����Ͽ��AQx�;#_�!D˖S�Ǿ��n:�nC+�\F�|���
&w���b��_���ɛ���7xq���������v��Ή_�:i�+���T!Q]�b�{�k���@�3"��*y��S��7~��~�oU�M�K�����A���`w�Dn:��I�l�^������V��#��ʇEǨ��	�$�^����<���i���`���q}����nZ_�ƹn�/]��0N��.(l��Cp�]0W���
6le5(Qn�ݛD���ꦮ�W���@e�f$:3�[4��\�ԅ�Q��EG�߇f���Y�� �~�K3)Yi����;�@J �����H�2��SdA
�o����sZ\�@c��|V����d+���(H�p^�a$[GLl�"����%����gը��=�x���}�$�����*�_tRJ�T�TU��[���F����y�)�wO���wx�<��{TF	r��N�v�A�[�Z����栗�8r
'��Ȝb�Cy�f�z��l&�2�V'!����ݕU�f��\�����g)�����׶�ڄsb��k ���6��+vW{ώ$lh�F2'�l�+}�h���8�6�����H)�CU*@1�;;S��%>�� f�}j�?zy�`i���C<&+�R�}���D���	��\�q3N=*v%��:˶�ʊ3�:���P�n.'Qڊl-����f��$m�?	�'L�Y�x�f2�B�+�nb��L6ʁi�T �;�򴃲�+�%�$4��X([b��Ŷ��E��k���|J�m#y�Ֆ�/xh �K.��u����Ш�q�D7��谿�zN��ү>
��\���]O��4��)Y��J��>_d��t��"���-ٷ����G�571�#>#�}W�P��b����iԺ���)�Ob鬈�������4��C�Q��"
�=�6�E�����"`�-����Sjz�K��g.�XR�A�]��oY���=�H�E��y))
�W�1l�iƸȟ��<c�~�����{6�gٌ0P/Q�G��su_��Z�&kǹ^��d���-tV����ɼZ+����>���l��g���ʨ��k�1b@�c��U�k,�MV���K�x �hd���L�^r����~p�����Z��s���������R�����}|5��Sb�f���\�W6��q�"5���xAK)>��Fm�W�eG��8�E�wb
Õ"�+ë/�>�e�W�({���Ԥ����������`�_%���i�i>�(o�3��u&�]h��]��M�<��W�Wbz��m$����~� ��-z����9�\��X�\N�>�IK�r�XcM,d���/2��&
Μ��D(��n�O�V�_�,�^3�"�_ �_s#B�b��Y�b�o?Y0�R��ިf3��X��5�E�g8�$�r���M�E$
��=�r�#�;�Aw�Qo��_�}mC!�ߜ\L�W��v`TH���eS��)(H�w�jq[o�X~��r9�0B�L��X%�̌�v��T��>���-`��ڻ���b�
.��@���O,���ф�ZB��"��#)�Y�����z�y1rw���8�&l��� 9:��$l,�R@f�a݀9��[`B�A��~�h�z��&� y sOi�-��;o�K;�!s��>�Ȅ���C%�{/�^�q%��o	��ȗ��S��r��>`�v`T@�5��M�5}<�+�j���C���a0D��j��O۔�Ӏ5�t;i�Ԕ��c_ˑ��U������n�b��P2:'�z�S�O5v.H�@""!���G	e��)g����Y��0O�K�7��0�.��cK_�v(ڜ���n���`��<��:�'8~tzI4_��c��ѯ����xR�������ف��yձ���:�1T��
ۣu�t;­�)��M��2�0����L��%�ٿy3��:�M��3&��:��P��Dqj�諢S3�U�{�!D��<�E.��T�BY!�'���V�R�(�+5��pQ�a�����M��#n8l�'��t^/�EZZ��+F��2���]}ba���#pC��\N��pm�t�t8��?6G���W,�jD:��#�(0|mk�!�G�x����L�g��ZB��G'mݩ6��?&���*���ܟ�;�l����C���O�n�o��w��ȋ���7zd�_d���9�c����v�At��+����0������G�/J��c|�٨IG?~�~��w*
mۄ�ÜxA�v6O3����/���f[C��K{��~ɛ��'T��"��A����TP�[iXҦ�����+y�#$�.�Թ	?���9��)���\xC�1G0�Bt<7K	����/6t�8*�ԚS��6�CZ4q�DE�"rs�i�����B�FPo;C��W"=!���dA�M����gG��@�(sW�����#{[%ד;9jP�e����Tbi�D��(L���y%�8݃��f0w��^�K����j��U��,��Y}�^�0���֑9����G!@��n<��Ȁ�����#�{�������jn����8�ɺ;�6N�g�r2¦1N�kQ�����@=d-<gJ�W�m���0��)@J�;�����L̶@��͏�C8A�C##��Lk~�l�[�7в��� s�1Rk |�gmm��ܢ���+;~C�2�[��o�&x_-Q��� �M�$.$�"�+�����=B��@2mfr�ߟYt�;7q��{�	���	@�
c��r��A�v���¸��0��*�qf1�x�}�n� ����t)F��"?��ɚ��*��|2�q|��:h� �XKR�k��O_K��8� +���Y1b4�V�v���+�/|n�	nJm^��׶Mį!2r��Mn�V��<i���2����pV(�U~��:���rR6o�~���Oy6Ԧ5���Ck�y���[�^��[�����N)���"7��K4(o��1Mw�j�'�]�\_���2�d�V%d��8'��Q�[M��-	���& ���=�9�bf ���2p����*��Dw�kY�{$�kЦ/�h��k�&B%�E��W�h����t�bW2����;?��;c��S�ˇy��� $!�WAJEb����R5ܘ6��	�N ����ڠ���{���R0�L�DtsuA�H[z�C�!���o!�אQHx��n>�()Pj�9UV���똏��7ߺԠW����§�K�p�4���k��L���笃���g7J[��<OE��W�dm>����?�Xr��<R�8k��֎����	/#~�٩�}��i�(�$�;:���U�}��u��$ѯ{���-�X�N�mFT{FA-�����6����f?i1
1<#*����B�I�kY����/Jm��>]3��v�� >���?��o�{����+���<�ݘh�De���б5 뛠S�������N��5��HL�BԐɸ"ђf	�9�lV���y�eҫ�9�ރb�a�6�����2@�Շ��)��*P��V� �A>�y�곢Geq%�C.�jdҊv��b0���J�θ�`w�Ȑ�P*O�l�0�_o��O�T��=�eP"Sm7A9��*�y�����Du��y��br�AR��&[_0fx�+b�x��	����۸�P���+cl#n������K�qq�?m7h���r��"u�>Ħ�!���~�n7�썞?ۗ�?I qS�y�����p��k�^F�������B�NIJp;-o�P��C��k�ܷ&�
�-��O�bcș��ۦM�Q�Z��v] ��b��U�����m��X��Y�)���S�#&�R7̸��D�mϗX�o�5r$�����y�m&�ج89Xz$��<�J�*��	�'W�a�$u�>1����D�R
��rA+�M��r�Vn��Ft\�)�0��,�8��V�Z�=��8 ���m�saM���lG���N�xo9��S�I��5>�]�f�p֕�)-	IUJh�>��c+��Ko�p��
��L� ��=&-Ο��Z��OhK�`rݛԬP�~L��\����-*N/��������)�]���H����9B�����Ҩ�t����p���U���x��g� �=+�
�;Bn�
�~������%mrIA4̬�
u�	e��ऑ��iU8y'�E�$�x������m���bґ�[qH3�8�"׍v��Ǒ�-"���H�d��$%��Ҥ��'���y�H2���[�g��C��)��e�c$`"��f��7OV�^���-���l"ui**T'O[����mC\d�~,��d�Ls�"S`<�6�`7X>&��	PUΰ0O��Z�r� ��Qp���C?L���	��o�
�L��'_�����TQ;ӿ՛je��ΊTr)}q�*�� � ͺ:�UJ�*��؉����4����J��s$�;2�f�W���a�x�C]�
<�N\F���i����-��f��p~8�z���s�ؖ�t(u�t��w�tü�^��F�kG:F^3��j2�F��Y��+Vp'��b��
Ms��`r�+1�L7&?��?���"��g/����+����<^k*����<�6�7�9����U���`��O|b'�J�wK�}���K���&[t�� _k�M����Z7.�6ؑ쵖���/�Ւ�B�Q��c�.K��u����X&o��13{m;�����7�)�
E�M�0�"ǀd�߆z�wY�y�G͕��d+@�:��+)�x��4H��X�<8M��l0����,�7z:<i��9��\}�h:cڧ���s)���cV��[��Ǩ9yт�� O�[vy��U<��b�"bp�	k�X��/�����U*�(� �&y��	
�LqMIAb�Ƴ2����I��ڼ}3����^�*e��h�u���X�Wp�{��݌r.���
~��͈��T�#fs�)�qF�Ѓ���ͮ <8aj��	SuX&�;]������0��|=��xھ������ O�>��M��/��կ)9�4�'X�[Oq!ϊWmB����e�����_���,h*'«��(��J��\���Ĕ�TY���k�FR²�1�:oWC�{���s�Se_��ax���j�1M1��W:��%��@��ё��FlІs�w�
�3
Y�h�S&U�@"Dhʾ�+��B_����`:|���`��H2ƽlԿ}�yS{��p�I��xlj��g�����x� _Z[�����30~5��#�+!�{?3�N�[5�Γ�5xs<�0Z���!��R�%��Ac·P�. ����%K�`Q�3�S���6p�U3�p(�F_��I�y�?fC��<F(��,'�׏����	T�eX)�ڷC����(�կBCu�S�ͧ��2�t�6�Z{��߮��npNF�a�j��["=�����A��x��_2�Ȥ#r���M�0\n��>����:	��y�>Q�Z"�O�\��xZu��'�q��I��85���w9��g�%�5.�H�d^b�s�:��G����f+M|E�r��ޡy峟��W(��)ݝw��Ԡf!���vrP��L挙�h:F���8u��H*j-����ӊA4��\�Ek�}��xY(2�����0��y���J5��G5s�R�rA�*�7�r��ߗ�,��yY�,�5�`�q�� ع���Į� ���(��h�V*��1�N���T!�艑D9�]$'�-y�����v���K��彙׊�O��geM�|.#G�7~W&do���y�~�j����Fo�k+ -��[V�R�,�&z��A�4�yɔ��mA�'�D�P������o�eu�9����a�j�#^U� GK����]��҂�H����~���ՓZ�OSmbg�	ܝ���v��c�*}J��ﯠ̸����`J q��vϚ�-F��Q��l����Cz�?ɾ���}��GH���a��^>b!��ou_-<��d�Չ����ZP��Ȗ����c:�^���H����Gi��b~�Z;��]7�ˀ��C;,KPW#_|iqD����r��ev���P�t����(v�;�]:�e��2�x�{rU�AŁBb�&@H`UKd�ד�8��!3 ��u%*�f�/���n�4~�װ���!���� �-1T�st����˫b�TN��_ye���,���ь�;�Χ��-hy_�?�\̷3,�b2��P�����N�k��.N��Wm�:�>)�i,.������H�{4�h�]���s��y�h��]��3c8���˕_w�E.�>���� k��3�?:؞2gD������gz(dc7��ٱ*�n�������/�	CG���#l1E�����ݝ��jv�r�u�d����2�j%�5�I�x�dD`��da���d��nw+VjdV��gRW�@&�:�B4��r/���9����Y�˼�"\i;<l���]��j�r1�'~a��S�>ٳ��耱|	�O�3�Іm�YK�y:�J�t�ݍ����i]eU����wa�*l����l�d��@V�Q{��5�:�Zb��(�ҽiRe	��9oy�D�t�@��Y	j9�S��1S�j�S�)ZuL����*�|�5�a��	ߣ��}��`6FSP���q=3HbN0��S�7~9ʢ�$J�9@���HؚY��:h͝������4�XF��f t���2i�"?$��_�6��ҟ˜)}�`��l�l�XA�k
ᮎ��:���=�w��s�p����
���@��=����ц.���P@K��Z�PE0�Qc{�/�=�I��E��B��h���"8>�گ݅�S<��P�_���[,ջ[{���s��E���0��v[���%S��(��'��8zl��6��Gf��H���H�5gQ��Y��No4�Emu��
C6c��VJ�+5�di��T�m�#����	���e-R=�`�!t�|Ct�t�l�����3�Y�K|D��p���	�h�^*"�]I^t�5k��}�Y�%�6/[/� a�UDCF;@a��>��Ք�����&���'��	�M�t%"���{k[�,��|�bٰ߲4!�G�ɫk-FxY��K^r�يl��1��#����}4�8�㲚@�C6��I�uI%����>�[��������1�e�ㇾ���:�Q��x�̱q�GT<|���(�YMאCg�������ZJ�D�=�����&�"&P��7qek��я:@뻜�A�Ɵ��$��s���u�qP�ʱ��zyMW@5� �� ��	�Ͱ剋n�ɷҧ`�����W��(���w(5�1�j�%Vw�'��M��*jm#�`V��ӧ#�pLd&,w�g�	~����d��c��)���Cn���Dh��\t��������z�ѫ��\����zoF=�נ�qcy⼰��B�����U0[w���$4���~؉���A��;ʸ)d���S�l��� O�)۵�ｷ2�q�̍�p� �KD�u��π�@�4�=����B�T�[e��]�[���6�PpH�D`����+�N�޺�q���Q��۶I��_}n����l�ǻ���XP��΍m����D��T�N41���ؾ�҄�H�{:P R��4��cҚ �ۑ/4�/7����������hu�͂��8Pfooc7�y,�n�0 ���6r��LN ���b�6�~Kl��*[���՘�{�&��z�y�g���B��ĿX���|)���՛�p��w�ͺ/Ym�����`j�`����P�9��)H	�����&t��ҘP��%��'Q=����p�N�� fx�L:� ��:d[(J"k=����L��9ӅІd�����ܓz����~P�f3/�'OC�� ���K�_�u��V���@m��_^�Q��'�/��ԛ���*#K�LǢ����l�N�+���1�cc���bL�	�
'��L&xt��T��Dd��Ҟ6��ʐ�p�@St���8�)Δ�}���e��Y�t�aC�M��jj���䎐���,�qC��lࡹ4�g�Eb���*�%_���SȎ-�����W�Q���c&	�v����i��Tm���e�����1�8H�������v��Lע���ɩ�#�����O��ĊZ�jAŤ��n�P���?�hc�?U�d.M�����y�˥�	���NZ����*E�:�О��Ϸ�&����`|��u� _��F*�g�h�R%Cl� #b(2�S.�Q�*\�P[qŻq�=����;d"������p#t
#�s�gFZh��V�5JZ��������,�Y�:������W$�D��w���.���ӿ9��'O:��S�*hY�(�D#�
9FOc�����<�FC{�Ư�D'6u��Mŀ'�v�t*���������_U�*�����!�s.����|7"�a^��q�1[���N`��L�Oy8������%6J�p��k6Z��O��ryBu���H�/��3�J���7�T~� j������*�Ι#$%B$��f:�X��]U���U��ui5�Y�5�Ǒ�*_�ճ췩	u{���ݿ�k#�: o�ݔp�z*e��h��a�C��M� ��:1K��!�ﵒU��u�0sV̘�1������c��N�Z!:�:)X���4��T�Z�65N��eG��0IR���Aw}�
J��4M4`O�H��K�!��Ptw[%L#�{:b;��ɒ?	D����'���vҪ_��-�����m��xw��͟T�%��.��4�|V}�%�Cd�*+��M���?Tt�����3>��	���Z���J߯E�/��ݴV!c����]�'悈��L�zF��g�uF�X��[
�&�ȭ@4Z�]+)�.����M》���vfB[���$?���U��%��Ȇ5P5A
n}oo��~Pݖ@�]Y\M�ʣ\Φ-����.M�9�g�~B%�zq'��f+��P�h���sI��~6r�s|�gmJE�݌7j��42�N��Z���ߟ2N����lQ�6�lL��K\�M���K��8�	\��g3�i=f?怷��o��C�A]���X 
B� ����|T���W57X!�vi�P��Q��ʆ���r9<�"�%��OMK`*o,r-�@gB���*Gb�?�+;��<<��B]���Z������S{	^P�����eUٷ)���Br�@^(W�ב��q0��=�HU���ᏻ������64x3�c�4V�
���`ld�X�x�yC�w���>�`�EQrm�Z�ȐR9�R��AŰ�^�3t�M�ҒGC�qM�P+М���M#����C�\�8��$��ķ�u���b��	����wT:��y2�T��s�ri(��T������p���Bjza�ǉB��zaKC�9_K�.b}��1���L�Ɏ�o�Xj>4K���E�a��S���HA�/Y��F�C��NG�������P5���%��]T.sw
���:X:�!yt��G��"uhYZ?bSi���i,�h��WK#��3���P�m$���i� ��LT�/�Pٹ����8TJ�׶qƎ/���}��hՊ��g���������
�P�6�o0��?�[���E(�KK���=IL���-�Eʙ�G S�ƽ��L���1͹pk���J<�A�է�X���� Ɩ�GJ�����SD�1HR�kq'm���5�Ұl��-+xs�bދe+z}�@�M����%�.ꠣ  ��4]�iW�N��<�x�!�V+��O3�2%1�,T̹�(�(�R��}d����,�~��H4��V���$A�R�*�)������U+(��S���>4�X�4÷�%ǐVg|Vkn�r���7����X���Cj��f�О�}�Ŗ�T
@���y^�r_8r���)��Y\�����1}8ry%s��nk`��,��o�mGLa�����w�̹�ccsA�9{�2��sH\�G�z���h٠��!�����"6�4�"@W�-7�5������ ��R�ff���LN����dx��x���WE����+��l�Py��P������=˫ �,��uv�fY�xf'�����g�|ؼ'�V�X G��0i}�t�9Ps���mS�p	x�x��<)���j�}~<�Q�f�Z�k|F���If,�����i�3�j섞2+1��p���2���q��x
�сB�����<��EQ��{��&���dx RX`R��&�<-T�g�J@̬�Ցk U�{s��C:�<^���;�N�8�	����ڄ�O4�[�c����N�Rü��4�FU�/B�w|��c�_�1��.����D-.��;��D}
"&�'�Uy�R�O�l@��]���r=1V�u�1�Kמ��`��Ț�[_b���A�ǔW����	1 �fgj�O[�G&.�R
-�:�XCftE���a%W��@vø#/���z�G�1�
�Q�����3�|Խs��?�^I*� 	9�֜W�zV�@�ٖ��Pº۴��DZ�q4J�ܷ���M�:D++`ۨZbuZ# ���F�DT8}��>��E��Pʡ�JK�Л�&������n"��t�K�e6������b%Q+�3�c,�h�����G�?��F�kp�|Rc�$�C �Hb�$�8�j+=��[�����"�"���(���W��/K��l"�=q��}.N0g�c �YqB˛^T�&�#��Z�ܭ�DU$`_	�P-dv/��c'J��	I�j�E��7U	�&oS���'RHy7�Y�jz���E�����'�l���~��3��}��*��М�dor�(ퟪ��Ukc�"�֖�
�T��;��B�μ^6D������~��"�w�Svq.�9��xW�5���!�T`],����1{t#MsV5��$�̭��_��� D��@�K��3�.xm����̲�߇�BL0n��:	�R�X�ASO l:4d���y��x���t����Gt1����#,�P�^]���b@TC-�L��#��;L����ҕ�p���5?i��AG���1����k�NEX�i�I��>v�n:��K �?����Zuk��E�4�*!0A���@j��[J�7�8�pNY��E��s"��Qyߵq��i+�����ܷ-�	e�d^4��&���ɓ˚<��}
�k����2,��	`�X�`�M5�3�:����r��3���>f3wcTK��Y/��z����?��X�NY����UZ��/�����&�G7-�|[Yi=5}��Bf�4E�ު���U�%�+��_�Q��B]i�@�l^3�f=�4��'�ds
�v��湏g���2��ؙ���'U��	�u�^��}�z�0Q=@B���j���`n�]�J���U�2���hë�x0�/ɀ̔'&��8��+�uH�NG�ˍ��0�
qȨ������<�ڤe8PB����Y�����^�--3�K��?Z���@��&��O2f8���i9Ҕ���%���\��Q�Ǆ@C��'�]�O��;'�urT+��)/,�BX�ؔY�����B���
3�Y��L^��,m����wӉ��WĒgp5���ye^�z|Ң�<�H�m�)��c���%�������?�;�ZP=!t��!���,S�u��"=��^<Ի�R)cx<N�Ɉ���x^�ѓIm��/쯭>�$��4@Mc�A���w.���BOa��OnM�R<ԄH�[��E*|�-��)�b̛�2K��9N}q�Ip���e�6�_��c�+��%�X��4sDBH�I��t�,�b�߂�������&��cY���a�)W��`}�U�I����A;u�Ŗf���~�������s8�"y}��b�r�4#q�1a���� �U!�Ÿ#�^.m�uU��t} � Z���+��S��}�i�{�k��B���_����񱙒��sK d�e{��'�V8qh��?��}���V��#� �|c������N�@���Z�*������^�bF;ү�o�]��K�ﱬy�X��E�v
�eh?��ѫ�,��g&Dv����Ѡ�_3{V��|fR�6U1`6��Nk�Us�Љ���U�!���"�_4A<�W��[a}Xsr����aM���Ti��͊d�{����i���I@�)Z���d�:Y�]ONW�rr]Qn�Z�	��	�x��=����X�Gɽ��F�o��`$�\���s�@#�ƨ�����{QM5L���b6�(�¾��k=��_Tz��l v�DiϸHO�Q��*[3tI����ܪ��ݚ�J�}�Mڟ=V�.&#��c��uw������L�w 15^��o>���%.�0gm����Xh1k�Ht>�pB#7"P]�T��^è=u"��Y�X�=@�&J}�E�=�n�:����d�� 喌�*�W�4�-򴛒������{2���X��8�:����W��2�S���Γ?���DUE4<K������q#�Sv-����r+�&�(�_YC;M���Y'�sm�}z�EJѓq(V��&z0݅���Va��S����YO$���i�4��\��ܵ�>]�0��$�ԑY~s���r�t�c-Aʭ�:AIm��d�S�5^�`�۳��{ć���	��4�(�����m�}ڨ!e����e��5~�Q��XY"\$�%��]����Mn���5|�@@\����y��8#.]M(�8��;E2���ioR�b2���/����B�r>�m�0-�Wʈ`z�m?��'uM���AŽ@�`^0��-�/��G�(|��Ϝː�&���2F=>��Wk{��x�>�����B|�e�����_�sÂ��+�_Ǿt=�q=:���1� ԍKt��!F�S� �u<6���?4����p���@� ��
Gt��H�h�S4��;i�b/ؼ��\iu�t��{+��C���_G
��@}|������|��+��b;��-2��y�Et��HEM������,���M8d%~r+�z���{�v'�n��}]yt��8���d��Z�4�q�V��j�W�S��Z��!+��j](�7 m�Iٺ��Sp��le4�2up+C����ć��#2�ح4"��6���Ŕ�WtQQ@Y��R�-ر%�gh����k?J^P��SoxTsCM	ˣ�(
LW��Sd2���=�����U?o��q�e3��l��Ea�����Z�JՁ��n�S(q3;��9��t9/|n3�mx��J�B�O�������ȱ�KD(���F%Y5���L��';\�x�l��E��j��"��.;RW^C�7�%��Mk�Y�A~���g��PS iE�k�v�oN�X����i!����گ�l��SD�;5e}X뀷��3�m�U.	7�Q7�|���^����4��sy�t��f��s�%м�)ɉm����X�`���������ۆhq�����,O��;^JW"�ʀ���>v���x�(Ja'G\nlg�~GmH��{�b$t�jX>\̿����!nxR\�(�$����J��#S뢓?�xJZ�X|�?�h�bgF�\/�
~�z4�[���^jl:� @.�-������Ttgo�О�t��h�*��ڍ�$]��hꂛ�z��T��lA��w�c(�w ��=����AW��(�A�9��u��}�UU�����M����W�7�}:�R�y�ɆJ\m���P�m�B=�9t�`����B}>`�.�8�
��2.$-�T?�Z"��w�0|�f��?PiNTa�?��o�5�p.PZ��\�	�rKtl?b�gPB��1�_���{�k�
���a���W�[�;�#ȇ[	#n�ƾ�|1pXbj��%��2p��Q�]$nٺ���8����f�X���z6�'C�"�nh��r���J���)����t�\�f����+8�����ᒪ��/���5����處La�z�vydnY����'� ��↤�+6-�,b.��0I2h����ʚ&E����K�ͽ#Y�����/����.&%��X��6	�����ēf�<��������qh��Ӗk<�x/.���.!�~@]s26-�a���ÎتT@9g�͚������L_Vy�=j�t5�t�������`���� �,FomR�rp!�`��8]�i�+x����\cYM��p-��\��Wh�!���%k�?D�y�.cu�&�l�Wuʯ}q�}M�R�ǜ{���I_�����7�qA����װ��+h-jRq\�Z��:6"�qMᗖ�āy[4N?���N�N�������XQ�<5�߸�z�12M��`�"�F?�fQ�u&M�#��.�O��������Ռ�';@$�&�"y+y&T���CT�A#��b'̏~�o�k��
ձ�����K�M!�����?RNr�vWJHPq�9�u�8��){��=�j��gU���*����~���'���(�ё���~��GN|~,("��y�7>}���[M"�v=�����m��'<*���ډN'��-g��ћ�ށ�KʭRCSf1|�(E�[=��du�a��Ns��=�ukk�ju��j���5��0��z�5ƣ��Km�i�8�-�mV:x�M�ж��?wn�J��Mk������u�y���aK��D!�茿�D�ط�mh
�'M���\$Vi:�&�����#����gR��<��=��;�L�o���A*P]h�g���m�"��р��+֎Yaơ�cv�ƪ��\18j=��i�%RV��zB6��8������&����k�&�~�xV(y�\> �Vv@]����Eg�2��_�>��$����nk��zj�3t����u.���g���TԶA���ȞR!@�l=i	C��ERt��p{ܵ�3��$z����$~�fp�e$�AZ�vS.��!U��30�����懈�:���Dm$��kV��5�Jfy5D�\D��L���=a������U�M�`�lo0����W^	�|(m,��ٸ��V��W��Pl$��OV?u�~�)Q�DfhKb���~�F��X
�����Dן&��C�9���L�Ke3N6Bz�����rS������ }�����V����2RfC�C-� P������ZS��F��M�4�=`�* ��]�>J��,q>����K�.o��~�F��b�@l��[/�e���+��,j?�,
o��XO���HS���.@�<B�=ꀉ��&ʫ��o�5�S
Fo kǪ�;����|�5ẍ.^bЉ-,5�p�T&[��L����'AAӪ݂?�u���-"��a��6�L��8��N�8��&iд|�Q�-\��wl��)>C�~�"N��|V��F?�үB7�\? �������j+4�yi�%'��`4�Π��l0v�6��R���5�&��Rd�O��uA
��̙%=|�B0��6�-�ઙ ����{��d%��(HMA(�-����� ��Ū��Y�>��=a�E���:_p_t��Up <]��߸�+�1��.��H�����*��G����F�HxZ�͙y�6Qf��(b����y����.�&XDX��ٛ��&�]�f�u�+n�.[~1G��d�~��W<�z6�	m��Ï���I�h�R���r|
?��h�ff�TfGD�Cu#�Џ8�����N�K�	��+��	:�h��r~g��1�JH뗴����"ߋ�$�k��H��(�C����E��Bئ�1�
9�.�$���D��9+K�M��}��,����|�)�g�e��o��~C��Sùs]o%���w�Gg"H�l\��_��Y�����"�̱�&zX��X��<�勖���-n�IXf��V}��qHM�`F�|dW�r����O%˫��+�����_��������NG4�,�xN�2�F3�ޕ�<��*K�@��ɐ�	g�A˵l�Î�v����
�h��$J���� �s��ϻc� G`S]��g�K�C���`2������Õ��X�x���\�V�Q�
�d�Y(��
�����a�1��=��y�?�ba��.�3<��l���$��������\���O/��G����D��%�MI����xpstC�l�P��z-ȍl���F;,�3�$��T?��0�`j���ص]����AT�SYx0� �	l��/�����T�Z��T4�b��=wd���ٝ�PИ|PK ��+Ҷm ���̚���4k�H�К���7�����:g��l{<:p�����q�J�Q��p~ݠ5��cGmyԃ]}��~�V|4��F1-��)���V��u��rݫԛF��HvcW�y�D c��`��^Jc� 
���HI4���˲�ۅ�������(H(��ǉ��P�3����K��~�M��J�a{� kTEH��LX����`}y��M 0��.�?����=��9R�~`[{����v�q��K����k5��E%�"S	�~��$�{�&%��]źZ)%l�VT	���DAAZ*:�pt��aSf���߰nS��ͬj��勷��w$�"~#����b�="�
?�(@��4�nFJ;A�G����/�TS@8�jr�R��oWG���b4�j�ko��{^�?��+������#�Wd".���gj\����
�[(������݀f.��cdF��z~8�5nM�\:�%��a����8S"aOf��-��Ѽ]OѤ���D�Du0�p���U�4�!��RPU��ր��F(��������y�Y�:�^��P$I��y%�s�T��V"%���3
�%���H�KDE�{��*�ryL�(e�gXv��ej�0T�1�X2f���3^DڨK� /⇍v��x\�H��?n8������ăsk���p��j&�ل����Sf9-�����2���+so���QN�n6s?��5%������=T�O
���qP���n�|�W%�ąŇi*F���ž����V�Ar �=�� N5��yVb��!ݭ���:�������rW׽	�U�^Vt�1I�P�q۵�3�_�_���R�y�bA��Í�Z�0�I,�Ek̨}~\d:�*��l��_tT�6�Z-v'��1:�o��H���=o]�� �W�#��2�,?��y]wa�;,��-u��!!�F��[+���*WM��l;�)0Kk��8���iKҬ��9�`�N) n��Aݪi؈��bU�M�K�a��j���i��-�ˊ݌,,���D�7|u���uÛ�ԴH��Vi+Vm�işWWU�]>/B(��>T�x<H����y9���?�A��bUJ&�� �������Ǆ��,KZ-��Z�?;�%�S|�o�&i���R���EO2�?Ԕ`���ծp&�_22+�ƽr����8�ۄ�m_��dH��B09��ZB�C�ߋ`�K��U[���QH-��`�Q�O�}_x��E����e���r�m��c�[�~ܬpxh��&���9��/4��W,��Fje��C*j5��M(�9��砧҈�ޘo���0t�� ��� ��G�o ��8�b�\�T	�|ʜ�r�,?�N�M�V������b�Vs���ә/'�]��� /���&lh�^5x,XzC�z��N�L��X�G��5�]��Z�%�ckΡ��PEDm��Ж��Ķ~��_�$�2��L��ͥ�����0��]�&g�o��#��g��8��������g*15+E)��ٳl�17��]��Ik�|ŋ��2��C^���8�D_Aup�^vс�X���A�5CzT�`0��#?{@�k*4,�|�w")i�0o����g��6Y���#[ځ�D�F�s\�M�AX��&��Q�,�`M�n���%���7Jc���d/`��jF�0�P	:�1�v�oj��XG�]��%�ߜob]
�k%�ܱa�]	Bg���u;2�8~Z`����o���
c`SO�e��ÛW������t5d���ZK��+w�qqE��t
D;�*h��?�
��4I���1�8�4��:a��5�:�eՓIZG�t�
�8W�#e.f��]�I�<�hr�aPW��
-�� �>���VL�`������-�C�>�j1N��2�,�w���MSu�����gGҞ���~����s������-H��ù&u��L�1�Ots��j�=S�4���%�O�M +�褬5�J3Z=%�MC��M�.�*��]��-��쒝}�4��e������y���5To��8�/�C3��^YٶԜĐ*����9��G�(o�J_�����#�cEY;��@.v���/}!a�/qnp(�ڌtH�@S��t�e�*��,5`nI��z4D��c���;}P��}k�!��fk�'���zC�:>�~V�����N͹giZ�!���H�k_�O�o��D|����a���J�U��Q�OYl�	���}ѓ�v�e~�a͋�����yb������r���D0�1r�i!�cU�$-�q��w�U�e�)R����T��$��PRlB<�<�ځ�M�:!��/l����X����R����S����Ś	�̮�i�p�ѵ�Z뒽�9�xl�o^�1�?���^���[��(�+�wF���� R��)���N,Y��#�'NG���x�7��ڌVA����j���`R�ˁ������۹	��z�#�T&(+�|:��0;��
 Z����<��/ȭ��Z0vL���EQ�;�%\�6�WI ��������ze�9�*�i,�>'�K�A>��¥�U�dSK
�\+r�*�w�(J����4�m�]��qxm[�h�G:�m_�,�N�)b�2�컬$�C$�����$(��0c��0׏�;$�\\�0�5
�e�R�xbJ���ƻLAЁ��[�'�I�����*LZ�SHŖ{ٴ�m����^�2>W��~�����Cƨ��?�AZ�yW�Z9��ơ���p�����C'S�e�V���d���f5Z���������GP��4��s�8l�-uޕ��\�2"O��"�h(|ظ�nDU�^Bp��.GV�^]�ih@Ӣ���f��2!��7��F�Ip��<�]Rr�i?����a��}�1�!������p6j*����+�	���k���W���qh�(�fN����g�B�: �;�n���vط�%&�ƌ�tp~t{��Y�eQR���y�AU�YA��#�2�ܶ��D}B<�FV�X	X�[С�^TJM�PTI"�ᕵ��^���� �|r.TKn�rd�C��ɔK�4�'Z����d�'�����tR�h��`�R�-�o"�g�$������ ���[ڭ��� �Q_��YB��2�@a�47p��H��h@_<��4�HO�	N�9�T��0^̜u�q���d�G��70��?�ѓ?�lO���ʝb�bm�����KaC���ൃo�A�r���[�|H���"3�U�I;���[j`{Y1X��� ��-�*��c��ͧ�{�.�-*�֖�
�h����@�J���d�՞Cm�nv?;��zJ�����ދ'(�%6���?�yܟ���?�r�?ܫ�m�W�}�w�I�ޣt�UW�g_�N"+���D��_�=?=8���dtC�[԰u��ޫt�bgS4Y_ݓ'�8�Kt�׎P��(�7��T��Ӝk�@��X�_�A�A�*u�a��{����5t$&yL��\�ұ�؍+b���?��hQ������~`P헥�Sy� �p۷~��.�'���l)��ښS��&C�7�I�0��\L٭� /:�l��E��c��|D�P���pFV��+�#�ʁ}�qd�<�Zw"l5�UM�e.����n���P��
�"t��_+�o��K?^�'w$�3�f�e�,�'
:ē6�*l�N��~:s/�e�$�%d�x�f�b�Bt���~\�#x���Yq�5���9^&����,_";ì�he�7K)���
��75j�b���W��̘T�j�Y@��vJW���an��8�w���:���4�����'̍C�s#�����h���q5�yf�Q�ꋩ���V@C�ێ�M�
��UiAxp$<��7��Ι3���R�|�pH_�8�@��C�b��� `%�j�XJ��� ������趸��8	�����z�4ܘ`a��^��{�����k�[����Z�)���SZr��:��q'=4��1N�o�n>L$Z{�?tꯂ=�Ά�՟5��K*�ShZBWm9�~~�-NGr���9>/3E�nzY跡���h��'��1�+�@e̽z��|�s"��#I.���H���.F�6���3�dN��\�u�Z/�t^�ƹ>%b��v����2�4�'���Ԏ�� 6B��=����6�KT)'�O��&Y��糖2RG��3�N�B��'�/��H8&ِP���_��X���Z-�~��<p%pRځ���H	kZ�>J;��S_������{aԎ�QMC��&�*g�F����_aP�k�v�I��_df��1��L����Y��r��/�_���f�[g�%��v��;�\+�2����ɜ���*���sMp����k0�ak��o�%S�%��3!��B+׏`u�� N���_K$m��:�8�{�=��.�3@~>��z~R�}	�PcV�䐺��=z.�E�i�y�F��7���q������5z����tF*��W=Z�t��+24�L�Y�0Y�I>�3���T��7A��Ԉ�Pi�wx�M�0�}$7KA46�\p~S�Y?3��\'��adG�58�ޓ5ي�����Gw���i���ߑk��\Զ+/���l5wbi�O��"P��L�oUy�q2���TP�?_���t	�@a��D94�M�]�vyo{f�	X�b�ו�/�f�N&&���>
����WQ�YK��-�;/���#�VA�vl�w�E���GXrQPJcx9�w__u�����Lx�Vx�C_z����2|����O����~��HIF/@8N�"|���c���.�/h@k9K�����ǁ��_VL�~`����y%ݪg�M���Gط�m�<�_(�J��V	�+/��!UU��=���d\O`fCF��?�Y�
-�H;Iw�6�Em�ޖw�ә��4�[)�����ܔ��	��g��b�����k6bذ�����o�b����m�b����2{i��M�t@`;t��A�F�Z�a��:�J�)?�����u�uSE��8}R�*Ռ���dW������c����y���u#1�`BZـ��b`�|#e�X'9&rl����u-���	NI3q��ΪYm�gbJ��%xs-�8��n�d`�'���1�Q�Ϳ��"�7t8Q{�)�<3.���������s@�pK�,Ƿذ}a��=r���=:)����>}��p_��FZ�r69(7����J������A���������;^^u�<(��;`�^NA#�	��+�X�&��,;P���5����ls��x�Eq���'���T�b$���ZO^�\w\��5=�W'?��O �]钡&X�\>�+4=8'�_�n�%�h��|u�"�k]�K��|,���^3Ҏ���@S�F���ͧ�-�-v�2I��M��_��8tT�5��u�A���?��M�EgL���5��2�!���4����"JR����T5H������~�9�ճs �1�]E��J�]�ț���Ê��z>��<��Չf����C��i�[��5�?�z��8U �m+1�h�n��2���C�s�i��XݖTn�Ƚ�ܫk��=�T:��O���o�hC��a)��,^0��A�kDN�ͧ�y�ϝA��S	�j(�
!nW
k
i>!Ka���Cv���v-��_=�|����B�O'F�O�I������~"�5&���d��#8D[�^�ZAQ9�9Ux�s�Iv��'��}�_ �k�!�j�s*O�γ�R��am쮳�?�%J��Z�慓��V�dsx�q�}��͸�UhҶ#x���3�$}P��ݞ��y�!Vv� �k%i2�����-�D�����P��F�5�� ��5"��e\�����}�Q9�wl9H]�84`����i=.ޯ��.�9�����u����۝;x��H�Wq�7��+����J��|&,N,e�u;���O��X�+�$��.�5�V3�i���jS-��� ����F�ZB	�V� ̠�e��W�__��
w��Yi���6�W0�U�.�J�X��ћ�l�-$��+%l��|���7�$1���;���E�%���ɺȮdi��	�j�����p�@�
Y׷G�)���]�O �pP��2���t�)���VaT��l�<��}j���Ə��ҿ�9]�ȤN�����6��_#J�!e|؁�N]� �}��#ty��������x��h�4vA٘Z��ja����g�K{�E�Iu6�^&�e��.dc�B�ɘ���na��w�	E�-�'���{.�m�4��O=Zެ��2�R��!+2��~�-@�Zd��	�8��p�Ef�:�a���r�4�5�6�IB%[m�sN��R8��N�k�rg���J�"�!�8
�������oU�322��V�:�Q-\�ۯs��`a�+�q���oa��O1P�KՄ�LK~�_�\��6C''����JP���*Ѝ�_�gQÒ~C��&��fX���$B��([�x5;��&������$ᙏ-�׈���Ҧ~P^>�����(g�d'}���+�o�N������)]�h5Gy"��a��=�$��xe�	��j�G�ʥN�\�N��:���8;�dfy���	0st�gw�O�E�K��	Ӎ��ʷ�����G�NbtƢH�`m/s��?Uqٔ�V��b��9��1��.�6��I�μ4ȂA1����Oh̽.�oMǘ�ose2�X�{���w�/z�=SCv�S��ExA�N�� Y�J&���s��5����n�|�Ѝ�~��1Dٴ�����h�M}Y�S�,�cŎ	�����lK1�m��	�R��A�:�'�`��#x�sAz�U�����'B���2��H@~Q1m}꡴5Pޥ�`�{�@�� 6��"\�=4��+��|.݈���h�ے� w��	�{���4w:b?n� Os�h5S���;^�q5�&�
o�'ǰ��<ݯ	����M�������D3�Ϋ�����5b5�D�;�춺�����{=k-QX�'�����3���{��-�\6��6���a�éJ~q�2��;t[��6fՀ����O���Nqs��.yi��ܧ��
���t:�A��R����(@gX�/�JRd�@�-�TUR��6��Q�E� L_¾{�4���ρ��x��ݙI0�Խp�C�����0Ϊl��4U��׮i"�D� ^ŋ`2Lk� v��Fi8�wM23U��
aπ�9����TВֱ{�̈́�z{�u�A����.G1��|��{ܮP��ؙ�+E�v_o*�(w����L�o��_;���h%�=�S!�@LZ���5<�:$�?���Q��/c���}�"���=�su�'Qk=�w:�����\�m�k[ԥ�.���0v̌N@��7C�Pw��d��3��,s!��/��Vn�Ϛjr��~��h�`��� __�βd��(6���[�"g��K��������1�GF�d�^�%++�J1��>Ѫ��gf�M�����!,�lDjh�8�����"��]Q�o��T��3�(WH�r�@�L�9�L��tc4��7m���u���ݪ7��3B+t�sW��R�ر�ri6^S�o��i'���y&��
��~�Č/J�p|�+|G�)8.�S��F�K:�Ϫёg4(��Kǽ��P�4�����%��[!R�Kz\����x��<�ۃ6?ɧ����M��c�	�����E�&2 �c�-%4G�AI'�*�L��R.V�f��kyrp@Î�&Xl�2����� h��e��� ���,\B��z`٧jb��!<�Y"�"L�����_{�+���/���2EZM�X=������\8�
�%J+�`)Gʛ��Mɚ�K�
`ү��]�k	�֎�&0Y�����H9��R�d�T�#�?��'>$���2���Q�����P.7j6Y�h�Ⱥժ ҠBL)P�n��&��$�0�+k6=s$��><՞�6��(G��Ӷ��V���Z|���-Y�AE�v�"](	h���@{�9qp�Ѭ|�Z�H����K�`���-we�p|�]̓�5���L��{�Ў�|6h��{��B�D!9���:޿���j���6I�&�9i���X�%��-WDəC��>r89P�����������xm[��w^J��|�PT�)�ȵ^����JIص;O6���`ga�촢�8�Y��'v�Xi)n�p�y�=����J�L��K���)���Yl�a���:����C24�9~�+�[Mb���-m��$@�ޠӕ��J��@�0��@�9SX��=�쎅j�������)Q$�)�2}O�q�=�.C��P��]��h�aE�d�B���	g����s�N�t�XҢ��5,����I&w�I7o���� v��%�m�6��2�X��8�6ctz��)���=�p[HRrہ�ip���xr����Lɍ���ҽ�۵�V��)�+�*��j�m
0���zƋj-����wrt�@��%gn�$������y݁�E��N#;�ng���pof/���@��'e' ^�(�7Č��댟�˻�ʝ�����ɸ�T`�
j����JN��&��^�+�t�GM��yV*����GB��b"��H�YD��D/�H�K�]T�"�EO���D
D;ٲyA�5�)uPZ�)��������5�����73�х���X��'lk:G�ϖS��s�g�\�{��4�ijm��ɖ�v4cZ�Zh���o�?+C!U\�(�^-*\�T`�o2��|�.\u� �'��0��#�7�?�t�w��bNd���NIq���LE��BPF�5��,F����0l���?+�q~2�O��M�-��oX�A*��:��W�������� �}Y�W��a�&���J�V��&gϡh�;�j'�ɒ7�����{Gz�>o,'� ����K$��N1���]8%b�P&}���t�i��~�mW/��R�x��Rq8`�I��]�,��V-f�0Yh(������Nϭ̿�1w�xEu�Lg��T����9�"��zZ�w#��Vu:uG����x�tN /����V�F�_�댾��as���9�\��c��]�S�i����6F9G�H$��\:і��&U�_x�S���W�H�u/'��-z-/��ӵ��:<�d �=���������v�J3V6���m7ip�]�����{��܏
�{�_�y�q�
P�5��2F��l68�ў*������*��SH���"@=���f��"���x�[=���gmV�<9��'dj��na`��J�wg���&Q|O4��h��CK��F�b(��=��|t�jfX�o\S�fZ��[(e*����ͮ؍�{� ?ڏ��g�����y+�P�gS���ާG�����G�2��h�V��I��J�}���)�\�����4���+����M�\8�2��1YY(*R
v��SskZ���f��&��ZŃ�i���\��^�cnbBg����2�'��Q��פ6k���D7e5c9�n�L�D��w+[;�C�n�-���·0���wh�S��I@ADj�ڡ̎.qB�=iz΍#������ՒZb~�#�R}C���f�A�ܝ��B����2��s��~XI]���n6W�r�Eʿ:�a�r�8����j�Q�ӣ�T6�q/�}�����@2-���d��#;�ql��oL²�\B�B��+��T��v���wg���� ��pd��Y)��.8e�?��~�m"�^����iR1�+ʠ|�d[b�����g� t�0�����
�	���~�v��\�Д<s�r�(r�{8uFO���ظ�	W1�~w����ȥ?E�NI��Ef����䳾�i4�[�VV��)�#r��K���Q����Q��ǯ�!'1���-��t��0��'N�q\J Q^m\������.�|8{g�!8��>nZX�]=�L�[%��{Z�Dƾ4=߅�哉���~n��>t��.�X�t���ݡ���'�,o�ç*NM�s\�`#]t�A/��%�,�XrL�i��U�B
IW<7Z=�����M��XuO��+Z4�[Y؍�f�^*D�b}7 ��@�L�VA�п)�I_ja�F1܄�6|>�*�/Ѕ[�6S�z=�kx�Yx�g��p��Ff����2>ޕ�L�p2�~n��d0����[G��٩�� �"�(nL��R�(x�XX(�dL̈́U���lA�:�(G��7x��
��}����SX++z�%�
lS�^;�z%�Āضmߖ��|+D͠L���q�*�i�i�����+��{-�٘,e��7ġ�\��\/�t?�[ߙKUk�`��X��%n쏘xQ�K�7pW��Z.��j,^M������q L���!����mW����`%00N����=^��~X%�rO�=�S�`5ҋ�~�aD^%�i�
���="bh�o�����z4����;�9�b53/�.5��ʟ�e������$^XފRz?�uk�n�e�����o����FiM���_�)�;��� 9^Dz�����(����n��,aЋ*^��P�#w�ֽ+Δ��'��e��q�すQ�����3g�1��Ƶp^�mC@u�")�$a�h���8Ε�\�c�4�\��g8���T�o>��X���ۇ�W�����m��e�k7�Z����^\�������,��֡��Y+ڳ�.7!�S@m�V���Ǿ�<�ϲ�XX�����bY'�����&q���8:��Z�4�]�~j�寝z0�.8h���5�4�R�ѧ�m�2�
�*�]}�����V"��C���tG|!Ef��d��C������J:��@F^O�������ٌ9M�{�%]rf__�x�E�!EQa�D'��-S���'���\�6M�ڮ��� cx}v����ޔ˗FG�@�h�p�3&�<� nl���o�B����S4�����(O'���Xn��L���J���{����<e�I ʶ�7�����q�
��F[���{������mK�O�'� ���#�E�7����˺( �O<rǍ��2	f����Hl���r��n3��n��5ާ��{�{F��{AfI��t�R���?-��}c��pm�(Icp�JK���b�@u*z����W8�k�~ɹ��������#��)3O4�����s���1�%���w�&GZ2���#�+�v?�V�/}I�����疬?���䏖�3�ħ��Z`����G{9(Hb�_����9B9�;D��gV���0�	��d�:L%�A�',c��j��}ga�>[�ذ���Q��n�ʲZv_�f���^'�5t�q�vza�lc�VN
��mt��ٜI�)���B���)宆�P?�!��l����S;F=�~�`uy��zN����j7�j��w��j2fO��6�RH�&�=��ۋ`�?������qk��	�ڑS�&7�(@�l-�'fy>�����r+�����Hs��o}�r��8]���"�~��#�IqPz �۵tډM��8&���3�mC,����kW��Z�X�Ū&)Ý��@��bm=W<mZ�� �Շ�.(����4u&����I��8�)�6T�۬�$Z�C�y��3� �p,�J�=�	�6�G+G4�C/�=��Ld²��y���I��7<���3�5�M�PFUs����R����U6bj'��%,���<�� �d�`����պ�+:95���C�IN4�U�0'�6R�I"���g������D�[� �	���s�M�P�dk���
v��QYEʅ)\��Y��fG�r���,ѥ�Ą(�p:Q�d�s�������9$��(߹����k��V)b�2�Ie�h����.��@��+���ѴM(�͙��G�[�q���Ͷ�Ս�V��X��*��*�m�Euys|�o��ٓ����_EK��m;�e���0�um�'Q�␫쾁q�o+&'�:�"4ZN��'V-*�Up��Z����zHLqS�^�~�,#d��RZ}E���$�
�I�$u���1�ZdW(� ����^�g\��;}��
d�.;)b��cv��[?��y��m�Eq�Pb�W�f\A����$�i���uaqA+�U�1y�[U'��e�$º�Q���������^z��U8���M��6����hf�@��˰"i�K����([L����F���W��M]�g�CLV���Ѥ�f1۶�Z�{��Z���S����~i)���^^_�I��=�:����JϚ�	 ]D+(�Ag&2��*q�&u��L���5a���`h�nA��l��,�1��*u+��0ui5 &��k��9�Y����B���ʩ�1��\^� �ϔOYH��ᚏ��t]<���z���"V��)��)���|���"�g��ı�z->ޥ�W�z�{v�u�qv�@������an��?�|;����m �7g�~'tE��;�ַ�[#?�ɢ��s�Ҟ=*�U����j/i�$;C_����z�"��D�����-���1EEP��?r��k����ý�ņ%��DB����#ǫ�S3��a���>��S�p�!��1�^��`vD*:�i��1%c�q��k�P���� 6�_�C��+�X��_�:Lq�be������	hZ����&�r�(�=ZV��g^mn;((�a|4B��Ƀe�N�������I��*���CU�[M�f�����k��<Y�x��
��nR| ��j�t����M� c2�|;\�f��%����4:Ue���Ao՚I%��AJ�L�2V[���#(��+h	U��52��_
/���{[:{���]�`�\h���FyW��E�ˏ�k�Zd7�	�L��۔�'$�r?l������!�x �FV��yĎ+ �&68���,H'~�zX�3�f�����j����>�I� WS�!��C%�;�*
������"2K�塖�M_��D%��L	 �e~�\� @3��=����^(UM�XX���2�>�d]����+�*�����Q��pl��-�dw�fc�e`[��o�g��Q�huTi!�"
J��H�hnM���c�R�������z	#��ݘ�P\�7	��y�v{�VP��S��!tiÎ�D#�w��_�ˀ�U��Dv�I�4R�О���ߕ��3q����}��T��;��|ȮR}�U�>-Oy�$�VW<!�_�E���O9FHd�'�Tq�5t9[�s�>#�l����I��d|��*�����S,ߒը�F�Xu&�j��m�(�_@��_��vѼL����Uו���Ғ���mK�q�@LZ�
���R���.H�.��]��d��&r�ս�Z�����M��U~E�K�|_­����2yp��-��v;x���q�F;���5�� F��|���O���Q��RY�7��� �AN��t�]�F���a?�0��uk��[�㼇*6�i�Q8��X�T}�"�����#q]8����58sMV�8[y���lZon\�L}鍯��i�7��G�&X�az.Ն� �K��!��Q�bAn�D������\j������A�����j�*�y^dru1E*���7 RyU��߾�k�S_�Jd�:������ˇ�)�ut����1�T�����+�zo��u�/o�b'�krДI�5\�����G��m
��К�?	J��ay�׎�]YAox���1p�/c\�V6u��	�	O/���U��Nc��m�����ʢ����;n#ՎP?�x]%����!��!|��|Rk�.�;���4d]k�9�g���j�JωS�.�ޅ��K���:�M�ˣ�6�H��"F��d
�K����v�1��P�xg�z�V3������7�K�R!NXo5�n���"��6����T����A彧Z���GEp����;�ح�w#�)雱9+������%V�_j�;��,�흭��$�j�� �|���De�\p��e��J�F�A�6�n����C; �N��J�/`~���.4����c]�X\  ���7�'}&�ۥ@x��;������  -����4
z!���7
p���N�|V�Y�7b)͜�o�f�=���T�A�U�#��T�h0fQ$8�b��Ac�jdć��j<H�_]L)�փ�b': ���k��<Q�5���y�����DB�Y��Ǻo�Y� e���=k����`ޯ�Z�]g�^���P��T���,tM��Sp��e��Q�f�|>��F�\bw;�Ȅ��[����i���z�՟����	o�".�֖C�!�9O$N���0q�g�^����8d��D�4�o����1�r�R?�� ��1S�H�v���κ������W">�9�|c��x�5�	8��ꂎ���v�(�7+-��5���|��Vzd�I�g�;g��S�k$w�Ԗ�,���m�:C�4�	h�!x�܈;�ۑ=�����Kҩ��" oRE��H���X�
�>MD#1�I:X�(}xs
)/>�V�^�@H=�>4�f�ϔZ��<��]_|����m ����S�N�V�`L�XQ��fj�c�J���+�/T9��Q3K0@�n��PZ���nW���y0��^D)^P���ط
eT+��kp�D�+�	|F^3s'&���w��[x� Z���]��y���G�l�Fa�E ^���_^`z�(���o��=�Ͷ�\N,�r��Q�+t�r@ �r<��	�rܯ��X `z8T���{�T�e#�i��Qm͢�K�(�p�9�� ?�2i��@<~�k���O����RN�{��*7{r��Q�1i.,��*	�I~���1Y�>��<����?V ����1�ܿ�c\��p�F5��r��1�N0�F(�����߫ݥ9(RӶ1֛4��V[���`z�y赣�c�T�����Q;�H0_��	��������L��&fVP�n��|��vs3}nü'�sX�n6�/�x�C������F�α�PE����z���P�J��WJ� 	ZC�2�;Դ���؂���L��L�]���V���-Yb~|-�]T�q,�]���4߃
N��n��T�P-k���gF��%�<�oJ9kHėZ�f�͊���8����y���mf0^8�\�T2)���Q�{&=����\"s���}\A/� �C���B���k�h�����Z�����RgqU;�K`q�Z@���av��19����\(Kȑ1/t��GQ���і��{��6�`�vWZ	0
$0}�Ϩ�}c�?�G����1h�PtAM-%\sE��of;^��FΧ=�݊/�}.9Q�y�6-4���������qZL��R8Z?�����Nn�p�}6h|��,lB���m�u��j	�I�&���=�k*�5�[���J�yU�Cj��p�J��À���uJ��� B����JJ�忹�n�|�����nj=�|�l�7^�v���𑵺5_έ�#'bT
� ���	\:�]M&����b	uw�V�����cD4�=����^h":�_s�'�:�itlA{]���c��^�C\�}�-:'M���p�cH��|��%��iqI��e��R	���ה�=Vǁ�#��/_��znwTg	b�f��mZZ,�S������/%�,[�5����=�/���V�55}� �y_4�ɦE��T&�Ө��7�r��i�Q&�@k�CIQ��ـvP�k���v��KP�`���G�d���5K����U�#����ՠ����o�Bv,S�a�)�#�U�am%��/���<��%q�4a��ɻ�5�LRI0�����W8`��cv9�)[�x�k��g�Bsd�jC��'�5c��%��VTtC��w�jB-�%C^jr��a׽_l۫�(��Zj�
1�@W-]�d�J\�VpzZ�,�k@�hRȜi��v���K�k�Q�5�[�8��(qL���8S����:�2���ǽM���f�G7�J|�� ��o5Q��y���IVh�%Qp���+�璠|!�ķ��	��0�ߴ�DK��LD�,˔��(T��\d��tf%�����Y�4׍�'�~����N��_0�G��u��QW8V�X�W��q$�e���3�1�2�X��i����8q�����Qd�}�]�d�5R�A�bZ�wv����X�\�K�D���kz�ҍ<�Щ�HZ�v�R����~[9��E���
��M���*;QL,N|�\�タ���I\�06�����E���/��]KTVfs��kQ��	ӵ��w��-��J�b���՜�ik�M�}�?͓'n����b.�2��~*��]VUo=��sb@	ˤ��1��k����&X 0%:�Lw�gIs�>���!�4���7\^�Q��n�x��b��]v�s�~:�#�.��w[�\�<l�p�3vT�f+��A��o�C�ۃa�aDGͨ^�^1Fl��9���Ѽ�D_*���t\��t�
xh�I�֕g�_ZK��i2pLe�3}�ePVHű���+����3�V�`��-��32��hp��X1Z28��h��w�;�1�uN�IN�<�|t�F$Av����. �[��e3}���[JT6U����,
�]���|�_ T��X��)q�"z(~�#Կ�4�X{�e.���P���`n��g��|���Uҏ��&3�ZV�<���篗�$!����I�D��9�nC�Ʒ�;�P��`ܴv�a�O�t5W�n'�UeOa;��C�)�I�w����EOd@�4������}aLP{���Α�L)+%A�s/�O=�(��t�Yݺ\�0�k!;4�"�$�����D���XsJW�;4+�f8y�7��f�yW��%�)����#���:;x��&n������`�c�8g
�]�P�Y�T�Ic�}YĻ���L��VDUݞ�D�$e����S�')�\p+GP�*\ Q�`�=7J���/r �R^��������b�J�ܽs<7ȭ���	j�!���j��K5.�����8pI��P��!�!M�1�p�8��ov�j/�p b��H�xҹk��R>T�}��6��vv`��+��&�*O�կ��edM��
=?��ܺ����Z�E����[�B
�YA'Q
SF�u�0���F�qY]����]�9���>UYz�e��J��_>��:���rpWs�G"�=�5�O~l5��;�L����6&�+�YA�ۓC��+��LF����+qs�>��[#���68)�IĦ�0�\)O�ӓ
�N1>mH%����<���W������[7���6�ȸ&w
D�[�$..�ؒ��%K�D�������7�}����tչ��H���!��g��D0`�Y���8���A�J���TX�W�Zr�t��1r�%>��E�f���X�s40��:���:>�2�k%1�g.q�+�$���uSH Yl�� b2r��s9�DIk�oXγ��M��9)
��z��²��<٬n`��XÄWE���ʯ>T_X�k_CHg;��1��Vq�H����k�b�8�gؿ�C�v	EfR�N��D�u�~3�_�Z�lJ���j&P���p3/���ڮ��UN(�a��1��н��&5B�)�sF	�擝2���N���G����y4��&p����<~�@��8��W��̂�>�x~:aEC�i`�4���'t�ZI�D��rb%<k��U1(�e�B�$a�ö��H�U�0�����pY1��e>LU�{y�l����bm$�'��8J7�ȵVI���e6�pNQ��'�^�+>�r��o�O�nLғ5���n"M�'���LU�^7Zՠ����Z�"��d��F^q�9�u'�g��mn�������X�)�ƭ_�F ��.HeSH�D�'�w�h�/򩵻h]���!���}׀�L��a����V�1-o�5�����?�0	��0(� ?�$�6� /��5��\�d�JS�B�G��.D���$dDtw�'�}FTJ�zeof�/k�t¶���>9��^D
����z2.^A�혔��8�kWϐ�V�Hp�I���k��]�<���]'�9S�O����%��@��kBS7��:�wEFO'&SQO�	�
$X�vV.}���^���s�Y��1`����`����,�W�W+�E�ر��C<�+9.�� ��jy]���񸻉�ʰ�A�z�q��;k�d�H��Y��`@o�QMu�溩ѕ|+l�k��c��>|�o�ُ� .ه~X�����?��d��Ic��'�ñ�k��ޅ��*�05s���@F�Lߩƨ{?���0����$�G&E��)��-��\�?��1Ǔ���3)�[)B-�J6?�]s!&�t5���8�؏k���#5�k���5 $4���Bx��p-mV�`��G�.+�?�mcO˲љ��G��U�����D�����*��bT��Aݰ�a"��H ����W�2B�8Cd�.�hd�e�LФ�n?��_ܛP��w?�ޱ��oO8��GJb��l�!�|D��}�3٘�l�B��֓�%�����D�Ʀ��&3W��F�W6�SX��{�����JO���j���V�b�g�r�di줏�u�!��@l�%AX��2�_�'�|���S���:�t!uvU1��o�B4���y$J���f���x���ٙ�\���[&��ݟ�K�V���#����.9䣞��G�����0F�D�yt4Z�S|?������}b�t�y�7��R�~��$�Up���x8�-���.�L����\����v�+7�p_�S�l�\/!P�v�S��7f����Wi�B{�_��tх��T8��V[H�R2��s�	p���P�b����i�OI�z_72Ţ��ܒ9��XZ����ؚ)���iC��6�	;j�,��k�D��̒(�V�r�#w����8)]�PШ��#�,ր�V|J���v�5�-p���>rM�IY��b��J%��>�u�%�s��}%��zX����B7+0wN��Y��es�r��E�d9��� ��J�	�G�Lݬ>l�ߤ�`4:Bys���DE����۝᪲/;�U�eL���V!>O�������Vu/����T�ä5֐yz�̇nvu�6��������^��H�DV�f�VF�A�����n��G�ݙ/�*�pW��W�Y�T]!Z�aku�vM�H;M4L7j���_� ���� ?�BV�`B��)�C�lSS\��O�¿�c����i��<eHt����+���7>G�xE4^Ir�5�!��q)]q�^v;	YB����m]�.6�\�G[`Tr��-!�n�ErU���1~��eSߒMM[OKeR ֦x<������6A��09�`�#�w�z��2�-�2қY�� ��E]Y��:�I$d�n�sO�%`'���o�H��A���� �dx������O��b,��B��ёB�9)1�!N+�Z��K	�vᗲ%���}#:b	<��,Ê�q�oo̯7�q4\m��c@"��u��/?���H;Ⱥw��㖳(��q?��9�Հ��a������z��$�5�\ej������#���A�):��uRj����|����{��z�W�/���1*�p]r���%��Q<�Ɂ9~��Znu�S�\�u����x�|#�ZI_.=n�}�AL�t��
�[p����m c��s�/��7	R~�8S`��R�{pcE*..$������ve��ח�@=3�p���AՌz)��O����ªe W��WM1O�p�����g߃����CX;sP'1Wp��]|��؏��}>�q��pz��Ʋ2�_���V�B���/���㕎]��v�	���u����R�U"��_AJ�CJB��h��%H���e��`�p]sN4�� �,�{����)/8�ҥIi5�H.H�H���w=�Y�R����(����C�_l�B��֚�~�/o��T(�M��/�mþ?��f��$>�:�z���n��t]���]�e�z>�"�c�\�K�<��{4b=�Kc�0r.
��as�����RD�ԍOﯹK�ޔ�����/>~4QZa*C�k�����l[�Ӝm�� ���^u���Q.M������m��|��57&idK�%V9�t.�
���C�ue�xȖڤ�S�����n�|��}���0C���d�ӻ���^൲��k��<�c!z�rs��ju�3�J�"�݄������R��iCh���Ly��ls
R�*�Eqxa��K߼U��E	��=�3M�=t��jF::s{���1�i���S�<w\�|��/DW�I )h�7X��`�,p$ݟ1��ŧ2��`1��1�7�L�c�`zs��{U�H�h���=~���t4��W4�!�۹��m����h�՝�������2l�)��x�k����}`��� �i�h�r��g1���4Qc4���ϵ葺���q��v�c,�������6B
Z^�d�R��d���Tt�.�t
W8s��[�G<�F��+�b���c����ֳ�F��WSLM��/4��Н��XX�.{�����?����������xg�Wt����=�ŢD���F�$��)�M��W�ڼjm��/OI��i�H��9W=�f[Z��1�5�ug{� ��v*��;���4����@�M\L�Q�	����17:�I�~m���I�F�Z�����<�5�t@�)|�c��wR|�r��O��?�޺���$��'�5l�a37O�0\	ae�i����kË���p3 �¯:���u6�gY�
	�]o8����wE,eb�2�+�J+����1y�����ӀЬ��p���x������`�*�����E�^G&����!Wd���������3�Qw�e�z{��_�i��Ӡ�����=�M.�� ��B��T'u��.jp:}�^��`u[fz���T��-�VTw6С�T���q���2I�K��X?��F����D!�\(0a���K㩴P�������aё%�zM�2\�Y'�	c��#�`TyB\��h��0�u�➜��{��OH��Y�/�܎u���E��(:�L:?ҽo��S�Ы�1Ja�5�
_0J��_�2�wٝ�>,���<��H���m��G����ߑ^V�d������#P*^�_x��U֛�6�Cԟ�7�~��}�%$�Ԗ�9=�^[.��PK��?o֜yT�0�M���)��<l8(����$	�w�?�C�)t��!����X�%#���`�4���6o�K�σ���_�lz�@�r@��i.�z���m�9��sŚ	�����N���3�oIő��<搻2�_`>*��%���(�Et��iK�V�S��lP
�U�R�P�5��W�������C�	�,jشK�8̥Tos�����J���
��B+7N�u=T��J�^�� &��1�~��������d=�^n� ��Q�R�y��[��4����'WWIق:B��t�i0er�3R?)�z���U����c�@�T�L}(�:ڂ�P�;3مM�y+/���V���xz���8�\PV�\;�G`jb�T\�a|���C�(2׷ qO���`�`�6w�ߦb��x����q��p"��Y����6���� B�u�Bw�Eq�wf���H��ɵ'"%� pF�us(�yllD��i�]��Mf��Tq��܊�bL@�]	�˿*.>��zU1~�+�/꧘7�@��˫�����c	�E�ofю/�B|�Q\'�����=����>���^��oq���?�$K7$��jp����	;���V������!�=�\r��T������:<��
>m�.�ܰ�Y�-�fų�	}D�������x��и��5��l�����AkJ��x	w]���k�\�׫�Z�7|Z,ߡU����6V`���
����AԦй��5n��@]%��M��x��=��ЁJ�[ ���i�0b����%�ѽ���M��7�\��Z�8S2�I�`Q��qgX�ra��.<�uH9���{�����5-<x����E��U�a�\�d�0,�@PV��䴃�k$qkA2to�A(���Z4Q��#쯔�Xz��Ӧ�����3��p� ~md�E��J
%�լ�ɉ��%��d��(0��*�+6���Y9���*���td9�l�+� ����j�P��F�tΡot&��بv,�0�d�a�����eR(�m�4���ĤJ�@`]!�C�}�V@l�ux5'�m].�!�@m�LO\��$�--�?�a�f�3�d|��U��`���і�M�����C�����>�F����Zc�����7��7Y�+[Vk����;6L/��b���K�ډS�y:.S��-u��7���	P4���/�y#h	�QT�Bu�u;&��n���L�z���xxP���(�*�0�� ���3�G�R��lBW UJ���
z#~�]��(�\Yl���{t*`���O�x�Dµ��9�`��,x��7�o�2(��2�K%T`y�*�%r�"����#};�6����L[��Mդ1]��ʎdӆ��k������'@*A�(&A�\۳sm�Z�蜂�|ևE�kyTM�� ��$]>A�ޜ�\
Ss1�����k�I�mjNUw�<8�fj���Z���d�*�8Æ<Cm��3&��� 5���T��3�LK]��`��WH��A�����G�(6[���'l� �rſ�1�LuA&����Q��R���n��>9!��B'�7��3���C�w�����E�.���S3tmV��U�b�̇�x���l2��qB��S'��>&��ojЏ;�W7�o��:�=�VR���ue�"�
���`a�`T��o�\��x�P̑7ܨ��"L���N.�S�B�lBf�H�m=(f	T�_�2���~�#"�/�'�ɏ���.��u���
E��.�]��yQ=_��yv��47;�$_��d��ٙ�1�^��+�|��8C�ʩ��s4���J����x��������> ��GdP�$z':K��!�a�B�`��KW�x�i2� hJ���-�Zxtx*�1��!~����(��<vGi�L���B{Ÿ�l��d	���)0�Z@%�$#NQ�22/B�����]��8+�s~�*
��vQ�p9)�x��YL��w��8� F��}��XjvT�7dXWH%)����#�ĺ����8��8|�/��iE���#<�Y���4�)��#3 ]P���{[T|�a6i��M5qϟ����~~_0���n·qb�P����N�؅
.j塴�e��jd�|*��(}t�D�%�g�F��]H�E�N������.�2p�n��l)(�5���d�����p;f�be��Y'>aX%q�`߰��X�.�L	I��rƈwx_�2��M��u%��}*�/�8�ʽBi�!iE��cӴ���Eз�1�������ub�xS����Ċ�9�kL�V��X+��UѧB�Px�"��z�C(@�+.���9�yU@l��S,���#�7 ����c�X�ޑ�J�͸C��Q�7�S}4�d�(���oט�e
)V���h�$~�* B\x�iP�ZWBu/�Y�J����O��M{Q���Cp���K��%3����4C��(�D���T�y��i��=^8p��F��bًNj�7���1��_�Q4��{�ާz�MEt��`���� ��!���;�����E��� ��z������l�쭸V�#Hm�Gq�Ɗ4+Ҕ=��イc���1�uٍ���ɘ-��90��An�b���_ƛ��0d7v;��f�VM"�E�2�,e�X�l{Aߵ���j�sC>/�HmI���������^�Bc��Gr����elD����A���K���u�E��~X���A_%ƈ:9��gQ����D�-�R�_�s"�0��un4c�M�q�D�����>W�1�Z��=E!xBKwA'D�i����B�=Du	_�ؽQBc����σ��g�J������	>���ŧʲ�'��(w��u?����O�O?����hd�����ZX�Y�,��!j�s������9��į�M��E�?�g��JzZ_��,_���`���������O�Ǒs��=�6x�� �|�2�fmk��<�5�(�z����'�o�칿�T��>�P��8g�0��m��Պ���o�:{�Q�=n�](�|s���r�4�,�N?9�������R�M.� p��1�x�S���� �\Ȣ�HL��Ɍ�q�.�)~�Ď��=�PW{]"O�:/�G�U]���de!]r�Ts�M7u��2#���2�R�����N��g�����H���%��޺�G���y�4���i �eK��wo�;ر��S��1�_��J�������!۴yZ^� GމN����J�� ^�<�7�d�&��."lX!�֊{��'���~w!J۷�3<:�+Sue����%�~ ;��j!�Rb��� �}��p���z�h�(%X�ж��Y���g�����)��9A��c �̥&br��a,���܆X�"g  ل�\Pʕz�sj�`)?�������%��dᵜ��pV�ث�:#Xk���~�L_�yHm͖�Dn�R�8�S�bV������0+�4�ɲ,MX�u�?J����ۼ�� B3N 3��VJ���y}o���&���>�Fb� �.^@�@���T��k%(E����$���X���B�-��e���ފ�k�p2�h����A���v5�%�9�3�:`PC� �N����h����� 6$m�E*m �J�f|�.�m��N��-c�<Q��y�W$�X��B�2���~@�����6H�v����~�A���k�)�AAN=#�"�b��'���G����R���0J3�E�R_aĂ���^`�?�M�~����םr�0�e���R�%��&ӯJw56���dL��� F-��a>cF_I����$u8�ں�!���<�U�fP��e�B��ƾ��&R@��b���t�h���u�?�u��8���n�+OH�$V�R$p.S�4��L�	y �ž�U�'h�,m���M�`��^�[�{�I�E��k�!�e�M����s�.l��xbxڒ�5��A�,c
�u^���y��c�Զ�:K���2ڰ6O+<I�5
R���{�I���&�ȣ��� ��uN� /6)"V�S� �ό��!5��	9��bJ�N��1��,��w�)���e�z߂y��j��o���c!e��Q�Ǹ+
t�»�\p������p�i\�Z]^�ǡ� ��x��
�B͗'RR��I�4�.)����YOcg��
+m�pn~;>b�'�ט�<�v�/�`����2?O|w�u-�m�TO��a�:�)�S�<�,���eԣ�oE�z������M�L�u�2��x�ȑ[R ���1����L�4x��3�Cx.�a�UscV��+�^�8�\�H)KkA�f-z±�&�X�a�&�l��aj=���)Z�)�\h�F���8��ybx͛��~Jgj9oK���+��2P/�s��&�u~�3|�☱�yK���b�>�|yt6d�$����L;�.79�ծ�?��[��f4QU '���a��0'*��0[�8�mojaP�QY�X�K��w ����1~t~׺�1�piQ�z�Y��u�1�:ӽ�Ǥ�Z����v�,�e���o�)�%Â[���KcyB��
&i�S����g)15�-��e��w;|t����m�x�� ���A
.A���4P�BP�egTMC�"����N4ވ14]�	���.[,�c�5z����,E��@��L�5��B�!�t�����y�����_��PgL���6�����W�Δ]$Rc����A�e���������*5�l��ѣ��U����k��+H�B[K�z�iҰ&X}W$�q��ȐRWӠ��C��)H*y��G1��E��b�>��dv��ܱƩ�9f[ߚ��ɮ
:�畤�n��O�:�$` },�W@(��b"4� �us�TCgǮF�ݧ���tlE���������"F�S���Gy��(��:wċM������B��qEn��+�)�궶�pXrܶ�;O	��|/j;.�w��' |����FLł��p6+�tn�B�V�К�-N�B�ј����_n�;b��\L�&��Or��'�LU#ٸ1��M��Ui����~�BT��?�9�|��d��q�|�e�E$���Z���@���c��ȳ΁O�K+K/��4MF���8��A/��]1k7e�����i�F@���٪�d�APh^������$P8��Bj���a��^�q*��G�⻰ �aa��2�Lb��㣲���� �jhay�o!-ew�7�=��P���ɌWgf�CvY�C�=%���-� ��lP��S��=R��K"��0�\,!p3E�U�l�^p��}�|���	�Tu�}�Wʟ)�#o{�V*�j-]�U��42������E��v3����x5��nԩ\����q	��h+�/|~��j!N�OOڄl���>�\A��z���XIN���
3Nǫ��)P�6ĵ/K
��N�� �d���f�V��,�F���5\�+A�y�?�D�yjv_+,}��?��J�v,@���4�d/� ss�ڦ�N�DI*��]B�F��4[U�5��Q�L��S����]S^���o
��H@Үڥ�M3Dֿ�+ =�%��Ǫ�C�KM�f��~?�U�ľo�g��{��H-)~Y+��0�,T�U��?/3��=8�?ϣI��^����ui�����?��Ln�Ic���\H��Ҋ���hA�K됺%�>��~�@��:��� {�:��/K��jB�y:7y���']���z����o�-ƾ\��"?����#9Y���'��i��\�p0��SX���a�E,a�*q�o�c2g p��&Ȭ�λ����Wc]z�ʄ�F	N�	#<�=�����x�g�x��ř�������y�@O�t�cq�8��ļ�;j�?Aj U��jى�c�o��ۇ	�����XY�pTؑ������!���ӛL�HnziT���a��s���'xp�0IK�Yp�+PO5(�9x�����S�!
>�](Y����	R�A�s ��E��X��m,}���C�4b��%��m1埌IJ�塋��	��_�zɒ%���$����1k �lP{JC%vk���<xR{RP���|U�_�7����D���q�F�6j����C'��_[dAπO���O�L��^���߇�fs4�1��b�eRG^�']�����h��$�HkK�1�bR��	z.
��Tҡ�X��Ly*Oʣ�_����Gx\y���O�}��D��xO�,Q��\ǹL	[0{6���ګ�ě���a��EL����i!w`\�i�ckCT?4J�O��֮O�e�����⏣�Ƽ.r�h}�.�T�[���]N��o����Cr��h'ˠ��i)�F��XobKKk��ֿ@XC̩x5qI���N�MM�^{��V�G����p�}���1A�J���ȋ��:�vm}x.Q���$ͯ��wS�J� "h�Ӭ�]mf;Dzmڤf�� K���Ԅ-�����C��!��ּG!&m�a�5��8�F���s[�U'�7�(�<�N���C�_��Ymh���xɥ�l�tJ!����_oEW�����rnk=�K�H�B-�����n?�!�k�Tw����i�����󍉤V�;z�hi|���jTm�ȓ�|����:4�P̖�D���(:-9*���[�R�J���l�b�v��P_���?�I��!Niq��5f*�玾~͉|eu.cKCL����ߍ�?<6�'t��V|Eeu��bW�Mۣ�0)�T�A��>���D9D�) �II���⅓�#�Yh�À@�����~�&)G�Rӌ�u�!]�i�0�>܀���˃�Y������bH�È�9�mV���Si��Z�[ٛ�o�(9�W�b"ZL�CL��%j���
$M4�tbРΌt2e�Q�O�}%d�63fh!%��F2}�~�e|��r�qE�Z]55�vgi`��lox�<�:�תd}� �M�j^��X��&C�r��z�ޖ��K&�g�nn����Xˑ��G��i��BJ��{}������<<_�����p+H�w������
5B�!l�Z��b��"�WSb^�����H�l�v��^�9��>M�=��8ɼ�>��X����U���;�I��|���)�������Ȓ��/�7�+Ƹ�k���ϝX�'�i%GHD7�y��4v%��sF�?I��@�R����<@�֦;�,ƱK�ڝ֕+�nf&YuKX��6��?+ q��'�� �\75L�f`��H�$�GyK�a �Q�~�̫�<�-�~�}iŤ��\��;�,m���%m���t�Б���b���N8���(K�M[+Om�:��h�$=
�@?�% �f��*�XFX!J�a�9�)S$�#��t)^=x���w$��=4�*^��y��jq/��
�����\���u�7ͻ�N>P���+F��Q��@)�{[^ Y�5��t�P�"(��8�qmE��GD5�QHb�g5G򽡤�Ui.�S3��^eΚ�b]r�-�Gx��5Is�6�]
�௭�ߣ�z.��b?���53��ڍkﯶ@bb��(ЮW��2P��M�N�����[��1�����N�g�#�\ �u��������M�,^�.� c�ng�8i_���� VI4���H��r���+MC���V'��u\���a���k��+F��_�S/P���J�:@@�yBǞLfvz����VS�m�H����C^S����m�2��3h�ܬ[ᕟ7����%�ΰ� ���%�وa��:��`�XGӭQQ]  �	��[�v���Ui1�,#��4�LM9X���找o��U��1�]�b��6�)�	�"�3|W���3:�A��5�,#�k�4Sz�=Y��n~�0óB&����1�	���٧�g�g#N@^I�v�:0���A��H�W�"H���y�{���?�?/�Awm Ņ@�1���u������������~q�Ե�Fy�V�� �ct��5�ܖս�+K!eC��/}6�7u��e���i��jGb�w%� ���RY*+c�
�RŅ�<�~b�_�C�?9��ּ|�7�7tǽ���tK0 2�A���/j8؟c�_�~��Oq��9�}���爢˜@��Im��v�DY�\���q��Bv#� ��H�[�$,�g��VsaQ��0L��Q���.��yW}@����b��!=�+������_��ᨶ��	�eA4����I�"�<o��ӲB�)6�����|�B��)�@��$Tiz�
v��:-ͼ\�yL����7�T�y�%��B0�L��\f�d\�C��1]�~�D_c%��3+;�.�)�w�=؍oM&e��h;v�!9j����Jh�;�}B��/��N�p��0}rV���/�P~q��ـ�̦?�
���!`<>K�`�D͂k:T����{�I�Z^�1�D�m�9'�v�������5���+�D���/�����Н���( H��C�`}ݍ)�=7�y����Q�1�6��6��i|.	43v�;iX�?A�����8�y�9'�^�u*����*��Ƽ��r����.g��!�!l���
��!N�����V*�qK�'�w!�^Dū��l����(�yF�	��ZO@�j
ǽ�b� ���e�<��o�b: Se��B��V��h��,RDέ�A�y���5�I{�a��T�!��Ź5��P�D�+��Sj�2�N;��F���}�pk2&� ~(sʮ��|�^��V���/�	��Fo�B����R�]>ý���kOQ1�|���[�<��։w�Z��Y�p��x�É����b�����	�Ox�r��V��˅dI[�ߓk����t��p�w=F���y�y�-�`AV��ۍ�-�lO�3��h�!�P@޻�E&zk�7�:���nS��N��-��K_o�1�=ڈ���5U3h�T$Zax	y�f%�&E�B�"(�I".lG�v�sV����r.K8EX/g0~���׈K=M���<�/#\t˿��1t{e���w�k8̍4�
ȑ��+���N��)`��u^�@O}z>������#�~���uU^��_Nr:��h���>>��f��~v�)�n	6C���,B��R��f4{O�z�ͥi�=�Ub}��ֶ�l[ࡢU�k
�^�Z�3���CeH�WO}MV*u��4��o��=�쉂���=y�	ZQ�}I�6�j� ��Z6	�.8G:�+	�E�ݧ	�SgD�P#n�+�Z0_XWg�+`E�A_<��Z	xPE� ��=5cnZ��2<���نt.�ΔQ
�{��ă��e��c�{ܶ�G���
�k���F<�H� z~%I9��%S7�Պ<7�	�m��!��̭A%!Ѫٰ	A��nѥ�1�F/[bo,>��V��ըcY+I&)%�}�a�_C���W�2ժ��U񰏣b���!���]��s��H�p�9�;O�T�o�+5����㽍.15��_�bO��(����j�T3�&����ND�Y�M�@\'��<R����
C9k�aW�h/I���Ka�W=�U��{s���(�n&4��T��%�Q�L�k=V���B�Kp>��^�i�M�T���J�Q5|F�1�û×��!��-�sZNh�?��2?���b|ؙ��ӈdE½�Re��e�%�����"V���6�_y�f:�6Z��
�O ٲ/T���_9:#;n��k��U�rM�{��$2a��aN ����v�+K�Qe�q:j��[�'�@��?i���n�)�땮��jHԇ&�x�rqNe+��!{m�7���>�8a�f�
�����L��|�����I�j�AE�3��w�O�(]�ȷ��1ӱ�uF첛�n���hL�B���`����7�4>�As����9��t��EYL\�8��(�w�����t�L'� �5"��4Kvo��x�U�C���PW*�����P�[�,C��!]��{54����$v�#�@c�B>�1H|��|hlLz
H�9�%3o�zb�P����>�QCXn#Oe9�;�����AUc�n�N��U�fH$�l� ���i�ʺ��@��l/g�yI���b��ֹ:gq%-���gC�6t8�j|em�9BvծF���94�_��^�N+n84����VG}$���ɣ;(JkKQRRD69,IBQO��W(�@4�<��i���nj�!�|�.����F���ˣ����4�G��P���rS�>I-����j}��M�m.p��nL���M�;_������_���G��Ż���^ߥ`2˹�������A��'b��\�ZH�+d�AY��M��ND�a���t�T�
�YOL�����C*���e�w +�C\�[H��I�X�rw�/���5,�������eP�S#���4lō�a�&Б�ֱK=�ΉhU$5�OA:� E���X4y��M�
�M�a�0�wp�i�'g��>Z�'�q�g��'�
�GVŮ������� BiÿM���0���Jf���'��涞���#*�i�<���51 �B�"�Y�;�����~�XV3���h�BRUj�.?�x�Q�_��X7�������mc\�F��Yd`��i��y�3��*0 U~sT�Ӡ��b~�:���ʆ�ĺ�	0�p���Ǽ� c��V���ą��~��u%���F�{/#��9,{9A���˄��r��G�G5欹�	��#�7�5OH�@#^=ب�ep$��w�����o���p�V�-�J��7 ���<�QI�������׶�ԫ!�:w|� 5��G۴�Ҵ!z���^9S�X6�*��li�(�gr�^����ߵ"��h	�N'���2Y�6���yoS�q6:J=�'��1Cc-�	xr#01Z%@�񙕝��VR�������A��!���z9Jm��ă�D��G������T��w��i�Jj�լ�$j%� 8�f�ڇ�~�E�}������!d�2E��(	֮��=A���K������1���O�?���,3�S	�t[s{'�X�վ�D�X�F�歳�N\J%0%$t���Vv����3�U�I��_�M�]����j��<Pg��uCC��~���|5.jN��>���.���>�ݸ4g5L��w��rN̨�ث��^iG��p����#�s�A[H�`�8�un��>��q�/�`l9��e�0fy�jtjۃ���K����+���RzVGE�c{.�7xU)���q�9�֛����9�x�0��(y
M���O�����̈��� ��Z���&���I�޸rY@���%�l�2d��&����4U��F`� Bi�j	�Һ�n�̠�1P�6�>��:1W�
Ml�Ke8��<_k���cw����R�A��N�����Ȭp)�ֵ�c`W�=�VU�� �f����O�wt�ǂ
�q��Rq
c0�%����c;"*%�u��H���m�@��H��܋����F�>���L�bs����4L�󰭊���Zc\]�g���;F�1P� �r��<ugzLo��X/��v�_W���p�]7������K��P�V�Z+��=����;ÆP#�Σa�4�@܀��i�6u�_8�@A�q���o����f5��e��YEu�q��E*yc�?]��W!�PI�"�x4�C�"��FUwk������k�#g��T= ��V6hp�G����C,G����f�4�낍&�6��Z�$�Y�)��Dxu;O�Xb�u��gֺn�͇��c����Ѧ��Bn1�Fٍ�5��b�ܤT����swm��8I����
�g^}q.���w��>��:������n^��自!Dy���N	�D��Rd�#^��}�G%��1��G�&�XD�ի��9�PUU&xؙl��v�޵~ػ���N�6�����98��t�y����W����N�e�fE��'� ���|RԆ��;g��D��)v\>�l��I��Ղx��`��t�}�h>����9������ݴ(�(b^��%�p�	{C
�N��I_��3A�b�!� ���<��¶=Ўu��x��� �Vk���er�[0����Sj.|��;�� ���3�kt�l��(��)F�E��vQ�4�p/���i� �Pa׌g���ө�<ׁ{���� -��;�N�Y�)X��QlO���iƩ;�B47:Ԉ���3���S�%h_�af�WLZׯȢ�*���X$hcGX�E0�q��I�C���ՀmP��F$j����"��\W�l��ׯ7���hx�O&��&4!>������Y0+��O�b���E1��琘���|3�$�)o� ��r��rnv�f9�f��xY���3�<�ZYumt���t�kW:[�~(7��4�f��NI���N�R��d۹y#/���ݩ;��3_�~�iظ[���0K�{��0�'��
o��1����3��'h�ɍ��y���	���_����T��o>7f2	���'�o�l�R�A>��121��*Ḅ ������Q]��I��������?:Il��㷐6sU�u�{��1��+���3e:l#*��bG�z�t�Z��U.�M�o_��Y�s�T_��1L�8l.��&����Q
�桳��H��1�rcN	Doo�U�@{o#�;��(y��zM�0$9=��J�~���x�3'���=l��L���r6�I��$�M�+V�Z ԕ.�/ub ����_���ą3��Mq��!��~ބf�8����ꂴ!�m�m�[.�F����(�zj���M;��L�U!���=
Ѫ·<��}Ƶ�9`8�z?K�l�Q���+�<�P,���SZg����$/BK�];,S��'��?!`���ILMx��������C�gTΦ���K�\:o�%(�`�t�T�5U�;wU�z*]��K�/h���Z`O=x��h���o��\p�"����8����.��x�39��w���0"�'�2yB��C�b�:,��aOP��פAU��B�h��ѕ*�����c�FM�w�z�̞��y���DW?���<�[�X�� �B3�{5�˶��Ž�8-�b�{}k�X7{*�M�C�t�_����d�6���
D?��<�BX��TCp��w����� ��R��9��2�A�`}��KU��i��s"���%b�Zv&��е���iY_���T�1��-�BN��݅��t��}o�?U��^#H!"�؄��ӕFB�Q�I7�ܧ���,>Es���L��7���~F�)���n�����$���Q��C�\u�,�ɖ�:�if���u,BdyΒ%&�a��dI��F��c�.�0�(#�;{�tZ��Z�@�,��&��ょ�H�:r�8���D-��O � 6��"�:��U<���������54.~k|ax�Ȕ��Y09^j&��ƒ:>�y�1^�}�Z�g�?�����m�s���{�us�a�ñ������G��'M��3'��r<?���>,#�kxB�^Ћ�(��߷��{H�о�o�M��>���u���p��� �p�Q�"�-��|	�J�.!*���2�+�X�F�-N�>qvw�5��G�׎�dO�VF0�����ĵ�q�ʬ�,�x浀�&/�~�q{nZ�K�팗#��{�?s("�c$�J�*�~�I��ߟ����͏�;�I�w�ے
M� �Y�	آ�U>p�BC�3GԢ��vkIa�4n!�F��|��Z1!s[io�jE��!�S�|"��g�n��-�����$�/���2�D�R���;F���Z4����&��_9�Z�!$�T�}�$�g�b�`�ϭbnJ� �)nʛvYG��iR�r��{E,"c��K	{�~E>+/��%,{ج�q!|`��֟��s	+�d5�q\~}/�w8셊�D�#փ��
���a�_F����Z��1m2*&[�I�b�& �F��$BLO^�^j�ǿ�eV<(�֯,E��f���r�t����W�][���$�`��V���0(�F�D=m�����y>��Ѿၱ�� 8���v�I�H$��1v�C��'�V�	O��ǀhL�J�_�Ԫ�7z�y��Fr����ت�}�a[a�6�K�9bG��3���֊)P��!������As�D����Q�['�(�'��"�j��x&|Gïᯣ)t���	��G`��^XK��dy�����b���ER��CBF��4�㑣� f�V/��� �5J���`�G�a_�C�c�#ť��oeF�n�(����I�>���oJLi���6w�����q�ܝ��s"\�η�Xe�I:'�;��6�r�Be���UC39_�1l[w���!�؏D�;U�'ݼxv����bjT�D5������+���f/�&-��ލߛ�S;5�B��RZ���T�9)��2qZ6��
 �s�~WO�%��Y�K�F�D�/�u��E*� �_���\&��_l�<��pɖ�*��b.�#k|lLKe�#�~~(�3�o�o_�It�|�O8�(o9sTv��[�K��N!�L6|�kH�3��Z�o-c�$I��c�C����.�|���IL�����q@�����K>⸢�Fu�*+��������h����������,��K@e!j�j]���J4�A�寽��a���~"QA���4�diY韰����8y�0Y�0,�L��@�oZ�۔�6s.L^�^>���0Wű���r�^*F�����D�Jt}�����_o;݌Sa�jK�������0�(p�ͱ~5#y�L�1���+�׈`��ʔ�9,dR<D�p���	���$��~�G�����ދY�mM�w�b��'Z�v��*ī �l@#�	2M��L-���ҿu��{ī�6����:-Dc���qWk%\�F�ԸP�x�>�wQ?���uY����y���>�l�ɳo��:�����+K�y��%�r���8�Qx�0�m�1��J[�'�"uq[E?RƋz�&H��a��1{�o&��8�ɳu�Cx�p���?�J����id����gxf�/�����&ѝ�U�M��(7�Y�XJ��;]�����6���%+�#��zUv� ���/�Q�=4Z �Cu'�1�@r��j�b ���d��}v-��&N�+!�L���w['�r�|a,�S����F��L$
�In)9	8�1v�3f8�L�:���1��v��Hмiz7���_���OTOFRBpW<;ä�r��U*����=K](�Oϟ�v�Ƣ#�$����4)j�ف�� F��������·����:w6��A8s�s��-?`���� ��t�	0�`�Q�n�9�0&��s;[��׊�r�M�?RYI�'S��3϶Bk��h��Q�����3O��e�����a��O`۞#��n/�W��Z���U��d��,f�0�0_��
e��	;^�R�RD�B`��Uj!�X�0>�&}��P�x��G���]G!v�h1I?�V���lv\sT$���.���XA����q���H-�������?_�
}P�Q>�p(�|��-�b��߽�n�jh+� �ƤR_�c����� �����y�-����5� �h��A� �$ڱ�U���,��{�,��PX	��3��q8tB�@�}���䑩���!�E-D���]S�O�W�B|��2�+�s~���?��w��;Nj���C��A߱'5�t�`�����vx���ZTS�v�H';;�q�$AE�<~N?i֯�\s�]�6��Y�կ9g/=�:���]}��)��a�b��(���{\_2�������RB:7!*|�1��QR�����k=)�.�͎d��b������B}�(�t1r/�Z]яq���jy�mj�M���1H��\�}�"HYma�}��%��Z��`��G�i��"Bk�3�9L�y��~$�p���,oBˁ�'�Ö�q���7���:�,�鲭�ϼ�U�|��D�R��-q(xg�*�z+՞4t��/@&���8e�������r���c��%G��V@�!U�F�;0�`�:�+A����{�Qd��Vvfٮ��ڰ�蚭��ެ6G�HaW�W�֡YA�U�e�l��~���oX��p��H�~�ϸq�Q�!5�	��G�*,׀%����k�f6 n�F��63���3d��|^��c�hǥx�PJ����v�x[&t^l�- pP�ll/$�0N�<�ۂ� /Տ�y�25"T#�v�����Ǜ�2h�8��[m�L�"z�J,�O��x�P�'N�04v��@W3*�r��$C�Toh�b�~s�}����^�S�1���@� �A �x�5hĭ�o��iND�zwF�q҆�=g���11+EG��E�D�"���
w�ʐ9�ړ@{� ��e.�+>�uT�D�Xب�˞�E�a�%�����Io��W���rq/}l�iO��*��_J��������7үEG�DH�Ѹ.�E����oB��lh[#��Q��nv�J6�sy:���U_/�3�$s����1��E/6I�+�ѭ�Q�5R=�R���{���Ξ���,U��H+	�e{����M����#�1_̻�kHzrz*�i��$�2a��W�_����=�=��,��3�"���y�k(w���h�Tjq� �#�hl�F�mvjSPoE�;��5!Q��<k	'�q8�  Vk��z�^u��E��Y����+����<���^��&c�@}�S%-f�WH�<tMA{=$$�/MW�p`���׾�#3S�����x�Z�H�]��u\�k&�~Bh|^����ʲڜ���,�3�2�	c�^�&�E�j���^��7�`N�C��|bb��&���b�d�a]+Ly�����J�$h9R��?$L���������.	[����1	� �!̲�2�`�z����B��+:����Ƽ�}�� ��!��?��{_y���}�ޓ�#0�GOw\� �����4RKf+-�}��4�_N��v&�I��2޸»��?�$���X�k��ƺ�)`���jTi-v:�ܱ$�}�x�Q�˟&�o")X��Ӧ$����BA�$�9ͫu4Z ڕ�܅�
l7üڧ_�k��@J�Hx�L�ۛP���I�%��N�Ս��g:5����<g�]�̊0��)�8��oS����~�+��������+I�{���*}\��h���g���5�:�(B�{3��/�S��: I]�������>uݾXw�s�`�_��#�	�h���r�
�-�j�;\����|?���!�/�B���'&i<�{у�=N��%���S=��F�.dGo���K@�5qe��	�i�~��f�srA>�"�1�5X�1�wH�&qL�@��,�����7s����@��d&�G
��B��B���hO��A2����^i���Rζͮl�d����= ���k�Y���[
���T��y��aݯ"f��'jܾ�8�ihj?���.7��D�6x���u��8�$вr�{89[K��t�U���Eo
��C�L������3)	uG3��4_��?�Wv6�tv���.ܭE=����#�͛��t/�v����P!�9N��	�����N�ȍ������~e5�:������]h�(j{���=6l�gc\s1X�U	�Q�-�H';"\b<f��!����u'��{/W/y��Y: ��E���d~��)�}� �)�<�������#\��iVE�~��ѻi�i9�(�і�TB��P�Ɔ?�̠l[r��|��m��"�a��1P5G�w6ѿ����L�CX�'�	��S;�z���w3�{	¾�pW&gU��$���։.vJm���+�gB�/(�b�jV�kG�BSk����b��q`�����Vqx��v�� 6���)�huwr�`y�3���ou����}d�!;��"�޻~�w��A�����B&��[K���=\�4�85�.(�d��s�ܷ��_Z?\C�OL��HM�>ìi��Q�`B�sG ���'� x�i����n"Ḍ-�IW��қ#��5bgd�[��+�0�ZuY4��}��R�wؾ^V�$1��� ��Θ�h��s���N�bg
Q��t4O�� ����"�l^�O�*CoaOy�j�Fú�_&�f�ϥ�kH��9�Ewwd8�z�zD�5W���z��}wZmL��db	�~;W�T��r�L ��Ӕ'��l�����ڹ혇d�]����$use�B��������$
�]�*o�Cc6���������4Q�DC�lcX8?��E�� &�t�d����� �.R3'M�7�}��"�w��l��fщ����|�vA=��R��{�$*h?f��(����w�bt�i4_���(��̻���dHC�a�������3?�B���\E�.X�w�|�4hk֓�b& H�������eP�Y��2�s�~gi��\s��ۗ�]�9v{�2������X��a�%f���9i��2�2��z	�ؠ���d�Q�s¬��<�����Y��_�� ��޶�{CS��>��ް��r�s=�̽�7�X���Y�,��օ«b�O��3�s��G���-~G���#/�D���^_�	�s�f}�GWk�kK��1
�%�1%S<�����Sdz���1ۅP��r=3��ᙖ�[��}�#��r8���_wZLw G>5v�)�ojFb2=69 Dһ6K���F�\�z��,c.��5��(�l'�1 ���6��YH;�1��b��j��LR�t�/^�{
 �z'����Z���:�lI��Ķ��2+� QRRv���d� �qH�[-^�Os��:ǃ���l�ȋ^��H�`'^cb���~��L�Mؕ��S: �-E�4sIN}v�.2��ё�[w��^M�5j�T�p����U��l|�hVm���������Ռy��Zo�&�<�,;-��3G`D@�,�����Mf?����	xՆ��t÷X������,�z��6����c-������/``�F�b.�Y���P���/^N��~C�uOux;�r9���5| C�͈��F��n���3_Sb�\L)�v
z�Z�_Nb�N<���m7���G[�A^��U%����x�wF��e���Y@sL�÷寔hXk������І����ޟ�Ry�T��#�
9K؀� p�"�-���\X��#�ӯK�пg����C�G�)E�9��5��a���y��X����3��=mI��K�2B�Ӈ�d���?	[ҋ�c#ݿ� �T!Z-�R5>��b"���	Є f ����̈7&VZeF�`F�g^�ؽ'�\������&ْ��-��\������% F3w�U��(3ɳ�j;&��T2;9[2�����/K+'��ȓ)04�������$Fd
BOj��E�2+��t(w/p P���H���)Ehu1�9���>��D����̯��uڕ�[�PH'"ӓ_���^����� �Ցը��{?64�b��ر"c��B�jPI�+m���Mm�W�8bS��z��,g�P0��uh�	����E�ws���.~����>��^OSrp��2��5N5`�:�'k��
(3Mxo�Օ^�?��6lm��.k?mR6������Z�y���% �_�d�㑯@SV7���<���.\��	�=D�숲z��E��!{tF=� E-��[�^.���_2;ş�{m�� ���-�~X�fǸ�Gt�z��Np���ʘa�U������픕x����H8MA�q�3����v�x�2G:�t�����\�A�HZ� ܁���|��9�9�  1B j&��3�������+�d��R��&�Ҏ�e�).A@z�����#7sޢ˓��AӖ��Z9���-����ϣh
I����:T���>�h�9���+U�� /�@�蟖�bŸx�<�P}m�h3���d|�Wq����Nu�x��9��m�c����8�4���`jZ�G���Nl�׫�R�S+�7,�wT�=<��l�8gO��V�����Z�Ɣ�N-���AVT��{�iח���}8�`Ct��߳�h��.UΑR֚�b�8��:��>eU��}��Q���A�I�%.ƹ��w��	��2E3@,��	�@d�#l��~l(�[�⏗
4��RT<�}�g��}U	��+�0@Ur?��S<u(�qS�"�׋��y=��#O�)����e=A�	��(@Bd�!q4�D�����
�8^j !��_*�,J�G�H%@����%���#��� ��������1� �T���5�>�8�t.�X�D�-���cx�;VRФU��ŭ_;����aT��9�$�=WFhi5<�+ʤ��u��;We���1�Aݝ�}�R�l|����&r�4�&���.ܕ��X��Z˫.tv΁7.�rz:���D���"˷�D��'�^�ލ��O��=c�=��LD�Y�-�q�W�=!����}�1�jO��lsEU~���)W���D5>�y�>���������Ry$�����R�g~���QA�í��ܴ-2	db�ù���HW��#.� ����?=/�*�ϸ��u_Q��4�J�����-�(�VM�I��D0��@
���^Ű��AF٦D&�F��V�ߞ8l�媓Ε]��d➒�)�e�M��'!<�4I$fz��[��0�,.�v✗�p%�[�<0n��gj@���3=�V����j6&��0�s)�G����<�A`7y0��4��Q�ƸW���,����|Ӄ7e+B+���[�X���,;$�̴�D[���_=p}���1�3^!f��=�:+�_�E��뛂�+`��$�W���ac���0�������ӟ�����Q!��{y�h��M�;uC�H}`nM��6o'�Pi��v�^���>�ƞ�ˋ5_k���dEAaVs�q�*~�ŕ0v�o�\5�J�M�,��˷$�,�w�)�/����W:-G+\D��Kj:����-�.�Qs��a�[�0#�"�Kz���z��.�}���D�^W �:�Oe	�f�zxZ������[`��BT��G_# ����$�����C;�����n�n�3�8�!�ۣ-��И(����n���f�2���n�g���4�QDK+���eM`���44�i�G�lS�9a7�+�*�D����$$�`	����s�-"��W"=�db��7`9����t��!����TF �deR�m�a0t_]=B��{'��,�3r;�8�yt������J6�[p����d�oW�����>s!���(�'��y�AQ��:��>�
%HL�A�|)��M���D歩�Z[�$��n�g$Y�o���c�ʐi�p���?q2���� �Yc��K���C��V���E�BzQw����e��������c̨S��l�"�3]RCP����
���"#�+�>y��nM>R�u]LJ5�=��$�b�Ǯ�W������$��G����:J��W�	�"�$Do�@}l��N�k�����>��a�Vz˩�oX�#��h��2�nNo�)Ia�3��i�Z7/�,�(��.ٺ�t8�D6�~�T�Ǐ��(�g[^ĥ�l�P�4���5F��U��M#����m�
��A�f�ga==}�'��U�ψM2OJ���-����U
�dJ,�~c��}����f�U-�}F�aI���{�6��u��k�ea�	��J��ow�!��kܺz0|􎶴�IH���u��%��N֯�q� ����s�v}oc�<��p���7�I��Z��@'L��~�Q�+��Q`��|����k�9i~ސ�s{2��e�,�)��t�٤�y���1���d�# +���}��g�� [��Y�C2�=�<���v���/x�-4�ۮB��)�T�ߣ�yO[7���xڗ.��������'4�@�bc�	��rh�t�*�%�	N�zз��}�uaGP2�z!�Ϲ�[ꆥ���P�?
�Wx^��ޟ��	ޏ&��N��KT�Ӽ\!t5��%Rz����R��8x�-p>0�x�Ӧ(����՗·��r�7J�&C���h����<!�#Q�1�Ё����v��,�p1�*�g�������n�H�m�Hh��-X��+�K�i�Pk���~0�6?�.ƋVjꄢR<�|1I���Ɉ��`ފ�O ԰�`�����\j��5<���h$���j�T�4�-J��� �~n�����u'�C9$��Zd�U�ʂ����#��E^�����M�W�h���?��ޖ$i��xGo�i�N���F	��M&B%0�� ߳���M^WJ�1�rh��SK�k4b��1�.��-�5�uo�.��n�
�g�Fw,����>���-g�e��o��{�w�cƹ�.	=�{O�_����M�W���ê
Z��y��z��z�'꠻]�V��+T	���'3�������)e��"�A���ϻa�.a���͓��]A���)W������kޫr����Mhw-�BE� ˋ�%O��zsS���1��b�K������2:�P{)�0����l�i�N!T�+Z�Yg�]�ت&8d[�ۀ�LD���ZD�a��������*�B���io�H	�r9ag*�#@WD�r��p��Vذ�wA���40�V߇Ml�>�����r�5�K�р#\�{bJ2G� �Q�7P�w@,"�邐t�V|^Y�����s�oyN��qX{%�(�Ζ���\��v���W�V�X�-�_G��*�7%�@�ß��0�P���|��ю.��3f���'��c�����0�̡��
��ǰ�_]
��K����{~>Z�~ �p�T-~���X�gD���{�M�I�y0ۃ��\���.]���LtE�#�
����S{1u�x��4O������3� 4�I�I�jZJ��M�a<Eئ����h,~ɘiΫu��D0�����#Ԯn <��9��M;(P���r7��ß������a%vM�8�i�Ռ5Ƞ5t��aR�(��P�m�a� i d𠤋�yDe_�f��ܟ���w����U�ѻhuW�B�Z��D�A#�4mC΍.�������1C%4�1̴I/�-dPO�=��f𓠣iS�l�yey�jc-U�i�
ݩ�G�.�����/��ŋ����,�qUo��7���+���a��|̒a����� ]�x���3��e/L ���៛�1��.��吔�Y<�G��4�(� ���.3�ZM��%��7���G���z�N��V����$x%��I]p�؝�K˺q�OTc�bO��\����R 	�m��"�'�߲U�X]a{&Ѡ�i��T2Ma���O�$��/�`��e�Q�M)�w�G�ӕ+$8�d�q�:.�"mծ�	�~��$���(�g�(�~�������8{(D���k�H�c�
A�D�*�4n��R�TT��"��M��$4��������1�ɼb�3(Az?SRf��:�>G��� W,�>s�@W#�68A�KoԴU|\�������/'����;ߗD'$�)�7�IT"��~��g���(b�
Q��Gʓ�/��A������Xur�7��^�xx<罁�2�Y��$/�dɱx��j3M~����(���_�6r���֙Tj��bey�Q��*�3?rb^�s�oo�0�5P�,?4��}���3 ��g�M+�
x��U�US��k��卓��\9v�Ƞ�����;�f�ʂ&�`~�,69��,��[EV�G��Z�c`��yh��[%��tEF<n�-Jn>��NE�紥�RE��'ޞ Fҥ��$�� ���G�-�v�0���S��_�� �6Oܻ�U�!��1�g�@0��٩�SqHC�E�OL𕒘p#N��Ы�5Q#=�6��L̆����e�
�CqLű`6�{-��M�A�|%A��n�ĵ�-\���mG'A~���Ԙ=I�xږB�&	��فa�j�������!V��o�ȵc�/�3�c6��$�3 r�*��������u��'Ky118[�4�� �_��d���L�|��+�;R��_�P]p/fԁ�I�5�imb�KV�>����ת�%6���9/"����B����?sf��/���S�����1V�[m��r�b؊7XC�E�^E7"�իm+�����bH�r�ߠ?�0�r�����)�E���<+�8��c�~_��z�qzed��gx�R/q�I�<�)�`������[��HD?%����'�\B��6}8�<@���N$�͎~ޮ;�׌f >X��V�th�m��)w�=�P��X����E�a
��.w�!���>�9�jU���b��"��y��JvAJV@(����Y�uc�Z�5�3|�LqB	�eQ�QLU}P���E:/�}�0�R��P�A��A�+�|AV��6�!�`%����񇆻|B�� ��Ò��W��	(Fr;V,Ei���V�, ����g(�t����{[�rj���M�0�H���>�R�B�Qh��ȿ���/ͫP����|(0 7��k�V�Gr�p)�?�14�bJ���l@�k��m�����@e'BY����6��]��C��ڿ�����l��^>棄�����c�
 �D5)ͭ	�����p�d�G��-uu�ò.q7F���#=�:n��+v܂���"a��:>��0c�#>�4�X�T.(�W	U$��Ȏ,k�z����D����f��z洲Ұ6݋�$@ٶI	���鼇�U$ճ�]+yEp��"���u��y�Bgd����ꈏ��^BÝ/�E���*<�kl���x�q���o�%�f��79�+djp?��8f b�1�
*BMӞl<̕}���Ƅ�E����FE����!7O���'[\���p�T�&Z�L����1u��V�dz�Tu�Uv��7�o��l�2��Y��	A�>�� ��X���_z��� ��K�5��W!E��ּw��1I��kL��C���f��`�ʆ���o��2���t������Sζ��]��]���1��
(��ı�o�b8I2�o|���QO��zi���W[`�����P�O8�G I#Nռ�,�Dq'���#���`�Q�x�p[�y^0-����%cs�d�,0��h��>B^Q�3I�H8C�0��>��4�Y����S��h�� �]~�["����� A�.��m��ʉ/IGhoշPz�:�|�Ƽ��ZR�b��w�Z[Ņb��kN�ث֘N�6(,4e�0�H���N�Ɩ��� �����4�2�9t�x�
Y�M���P����}:��S������f������Z��ʥ�_�D�s��K�0�e'G�L#I	[��@.�^�� |:J�߰|�JwZ�v9����cRq�����.�>�0��/�j�)'?��O�mУ��1ū%�Y�oJ���83���w�p�Z����4�JU�w)U"N�h�Z���2<����N��z��-J����)��Aj�R������6��[ޜ��`����5�`�󻂣{�EH}*u,H�?�^�(��	(�c�]����i~=���1пB�Rֺ���x�$���WZ�oW���&E��Fu�Y�`Y��DR�S�W� @ �Ӳ��^m��GtbN�/�k�@�Zd/�����b]���գ��a��-�[f1����O{�q<���d(�!��!�f432��F6�O�P򷧤&>v���YN�A�E"������Z��B��yu�v� E(��%�f�^9Ri�j��������m2T�|Dt�&vF�"�]�k��_�zw�������#�?
0��gV��l���{X��������B���(�n&��Ӻ�u�ҹ��>��ݥ߲C9v1yY�R�Qz	W��d��0��;:Xk��sc[�\���ݼ�t��Ɠ"�祝Y�t��g�n�=�(�٘jX��;5gЭ&(�il���G��~U�����]d���D^�	������º9�0�@��~Ŧm��P�^�V��d:9����n�`5�rřZEl��r�"Q]�T��^OV8�>Ε�sgI�CP��Ζ�v�t�P��[�0BT�XʆI$̤�
G(�m�4�v��C�"��&�@C�-��m���f�]�1�rg2dI�Ii�RXS�RXH�њm��6�� �˩��$��ۮXf�*�fZ�º<z�n����[�g�T�ˉx@̡�}w��9�D`1L��8m�xJʓZ����N��102l��<�%]���Ӓ�C�r�8YϨH���4S���8�H7�;K�ѢW���J���PL������*�a}l��a{J��?��B��L��3�[��
߳��~��1Rb,�Vd��VP��H�VJ����<[+�[�f�{�gN9�b�ܱh�9*wr�cF.�$CPe$�޹m�|'2�|=���Z������EM��.č��1��Dp�<\�-�fg��F��XI#Ų��<@��{���_-C�<-��1�l�=��O]&���	#��Xڄy"Gd
v��"&Oi�8UL�DE��A����R	6&Α���ݨ�L�'��G�)�7��h]/�v��Ӣ�f�勜�4^�q�59D
dcP��OD�:�������׈K�qk�:@,�!T��6 ��&���!m��Y��l@
�B���9���c��؉I��a˭�d���]��y�=JI�\�x��m����U�b�/��|;#�!w�����J���Oe�<�9�р8���{|��ިփ�/ƽL��k5�,��2�-��a&�����)�5Z�HngD��p��ݡ}G�c�g�������n�����&����A���Gstz�ڙ+��|2"�,�������u&m}�J��ʈ>{2����ʘq̵7��֥|u�r�������x�O٫�@@K0]X��1��;�,����rI�_
�4�	0qM��O��7��a�X�tI�蚿��c"����ēY��R�e��K����-�Q���SWż�}��d�p�a�ڛ�7t���jU �!��
���]Xۤ���))�w���|Ϗ��s��]��"j�=[�SN�x��Q���'
h�+��Ѩ�峬q�ؓ�έR}��_�3����N�gM���:�J0��?��$V�M�<������t-�e}����MH��m��߆P�^�#��ҳ�CZ���/��B�f�M4Z�(�Q�8��C�¬�A��-;�r�m-������L�����߂P8^��M�μ�d=�����MdO��2�$)��"�������r��(8U��ݻ)�k��R��%���k��^6(c�"�@�C �\����0Ȱ����E����f6ק;�����Xв�����cJ3Ća�^!�t�liW+�xP�:��s��Ο��d��yuC��;��B�I!��T��h���~G<�
`u��m�;}3�%��\-��w�`�*Mv0֎��LOm9W�ǀ���y(��B�/�X+�W��t�5�{� ��GP/���;0Ka��5��ٞ�䅖�������0���YA��oϖ�!��j�擧D��V,�#]ˀZ~��O����dʟPQ<	r>��h�0"o8`|m�G�^�`����a���%ǰ��O��;3D�Τ�d��&��~�c�C=��'�G㾓�1J�`�W��
Qf�~W �J�Mw�ȋ�ٯ=���|�#à����M#A�Z����4�����'��9����(�7���rR�0pJλ!�U�}n��8���{<��d��%݀�?�>� ����E���qܺ�oT٘k��t�|wP������#ȹ;�����?�u#୴���9�j��c�[>�B�Z���K�h��k!!L��)�� 6��Q �;X�B��%\$5��}�f�B����Y��ӿWR&�ϲd���)��ݺ�����^�|9���p��ma�O�2-���r�5��7#��C��)�����+�%>݉�;s�����.��z�Mr=����BC�,6�O����}�_��W;BϾ��T��',�N�&����*ݶ{��n�o�AժX�BUV&��� j�:�����d]�;3�=}$D���лp���-��{Af[XR* lG��yY�Z�&1X�����-�G��M�v�����ٖ��z4��D�W)	;�����^�_�����.��,o![��	�]�+b�&0m�d��!_2�ߡ����[�W�[[J�6e[����GaɈ��m6��<��e��A�	
mg�tK��yd|(�й����A2�;a?��p�3�)�4�D>5�SG;��o��_�=�yVn���u?(q��(�3�Yf�?J���^��/�=iL(�c�&���/i�|+������T��B��d��t�_�6�Â}��FE{���T(!Q�Gf�}o���/���k	x+ŗ5��Bt�xk�J�R�T�bA��9n�1֔�6?��ږ�t4������f�N-�z���Y��	C��>Jv���v���
U�����Q�P@���6[uq�s�u�9O��z�	��m�y&e���C�a�m2p�vl�H�����i��G�����s�;>U��+�mH-T�s!̕�$Ұ���?.�Y5�ػ�2��ecգ:���>z�ÈvePy�m*jqEJL��<7zFY,1j]�,2E�&�®��=��9k��
Ɉ�C:M�������,��m�Z�]��T*T��z'*J:���7zQ)��H[B���/kT� �����
�E�±+�K����4��U$+�E�� �/(y���Q�����NLyU-��g��W'�c:{�p�8��Tr�B��h�;��iM,ڀl��}8��!v˲�x�M�>l�p��l�p���k��~�lO���a� m>��)�&�[��8�kX5�݆86}�P0���w�O�>�¹.�e��������a(�f|�#��P�@��#�q��Y�"l�ƉL]l���CJ<t�b��w�X��:p�!���_,y���5�S9���<!��/�ŭ���\.�ꕎ��QҺ��{wǖ�-ݞ�T�T���fhH��}n�h���or�|F�Š�u�n{lC����#�c��L:��)������T��6�m���Ez-}+���]D����2\�1�&jM;�z����l�-�)Y�Y��� ˅Uh�*�b�>�����<�Y���ɿ�O���F�;�<}�'&�!��q+����oRu<`�y^jfx�n��t�vt;ۅG��-�0��+�yhM W�p���ְr�W8�.G��J�^�g'���^�}s�90��t$��zh���k���܋�����{kq$�C$W�u����v������#1y
ʒ�~L����w5��XJ?�t����B�5�|Ջ�:�����+���*B�a�o��*�:ǪQ ����7;%B���;r���򜒜hEM��iv,T&G�u��f|ֆH�hb@������D�2:�Z����-���H�P�����o� G�Q�X���Â�͍�<�렒{�&IDӄ���'�-�*I���f���+���
*�~1:B6���f[P�&��b@��#ZB�����p6Fʁ���q1�m���3���/:x�5��O9X��ϺC},es���G0o�*؊5R�Ǜxc�E�˘�׊鷵��0��m���=��T��H��7Ve��o���fʵ��~B;3��W�����o��v�I$*=�J�|=��\���	!p+��CɁ��m��`yM�B���Wk����`j�۩�:M��o�7��"��K��ҍB^�TR<zކn`�?���'�M�kM�ޛ�p��#��6vik�g�Q���4�yNR�l�V~�ذ�G�ҴQ�������%���M�F>*l��pOE��p����'��f�Eg��S�r����#ϐ���qY#��8�4��O��X ��v�!�^~���}a�������V�ҷa#�S�4il �����ӈ.���I��;R�S�}:IyA�LW #δ�x�b�<��tR�\bĨ+ vT?���:�N=J�XM�ˬ�7�d��o�	��Ƀ�@��(`�2c ���s��}�8��tl���"��>�2ȱ@_<���8�.!ރ������Y�D)p�t�=k!Y��� }�� ��U�&}A6|��t���O�_����Z=�e2T;5��/v�燈���|�`	Mo���~�]��D�����ە@�8�9�P��l�!6C���c����F�M򺵻]���)�)&�C�|�ʩ�u�di1NK���� ]�xo㾊��T���{�=`��y0��VOi!�P6��Q�����u���)�$M�&z���KWk�x{�8��wwi���c����Q�����T���i=['Ón��UjJW���ce=�ɉG����4�i��lt���i�LB��)�P��������3����'����u1p�S|7�O�eί�x�ȉ���ۍ(�^�����(�ܤ�8�"l4Ad�� *USݥ�-��p��Gg6����8�}�t%�4��|��ʳ��L:<�2�@�MVz4v
*q�ц�=^�M�[��+%Kx�v��pq�X���A��0�W]�������.���k>���Y�#�����*�)�Y�(҇�{1�Z���9����i��eG��;����6@��Ak!<�31������7�LR��R�s��v�
���^�=���a��وX�!�a��o���":˭��2F}D7�S%�� ZMau�����J�����-���}6�Q����eۡ�"Q��� �Ї(��*�DMb!��>xIf�,�~����DnB��W%*0P�<;���2¨�yq���zMr��=Ey�G�8&X� ]�[�Z�� ��pD�l��Om�S�:+'R�4���D��7f}��!�gP]o���	h�z~�K>NhsʶD�o2գ;����,�o���9���[N%����A���������(��:�`���ZoMZ���M�uUNN��R�v��,!wXz��h�\�&�ί{O<�q.d}��X\�O��r=̯t��L���7A�d��QE�p?�|:���꠻��l ��p�@��Px�H,�Um�wb��"��۪��T����{7����+���,UNÃ�d/��ǬX1}��W���/�a�BJ�}�DF`��:�0� X|s�1VvXr�u~ʵ%/�R��,��S�0S�pNl5�OM�qP��a&��嗌<����Y�
}��r�dw���	�	�JRl��
�(��8�)�]�V�5��m���/��e��A����c�h����*�v�m�b�V߭>gz_�/uq¡�~�VL��mf7���~�_�;�qe~n�E�X�X��Df ��O�{����$gۂ�.c��jt�?_�͞���#�PF	gy�5�1H��[��{c|���JC�:��>N��hB�.�.�W�I�c�����6|�����3R����dY�O����l�.k��&��CQ�W�SZ�J��=
��wA�e=7���fx1C�7dݧ��������Iv��c�����k)j��ܻa��:7)+�K�5CVx��|9xL
���H�Ʊ[C P�mҹh��,�c���m��}%�wx��Z ov
��>,��X �.Y�e;�+/W��d���I!��v�@
�;�nM�ÁΟs%d�����n�d��}?��*D���d�� �W�
����n`�f�zx'���C�4z��C�¨T7/����������^{����F�90#մ��SZ�ȣf(�H�#2Q𞼯�n]'q�g-��Ĳ�恱D0<�rVTE��ޡuȎpJ!��"ٞ�@�X॒msTw��F���1���)����ֱ;�@�޹M�q�U-���O���͟j!�[A�mzKv����=�����2�
���&^�[l���)%c�N�u�j�#<T���	z#���:ua�B��ki"[`���r���y�����F�7����Lϗ��hd�QO�S�����_aح�y@�(�e:%�K�Q�YC8(�N�D#�����l5JB����A	��)k�" �wa��y�p�[�0{<N�m��Ң�-�o�T�}~��Ou�J�w��!����)t�<�0�r;��gm-E��]N�=Y�uNڜj����3݉�*�7��!�O�N��C*�b8<a��n�6(���XG��C �s ����ǧZb	]Lۮ�T��-g$����.���2�Y��6�}�&
�7�*��LV���e|�1�4���L�'��䬂�tf�LG�[�4�2��wk$�tC��I����sN/lM���	<8�HN���E*
�.xY�K�E��Τ�v��� 7���Z5���D�� y�.��� U��{���^E��-(<Z�8�]~��e��|j �x_��o©����GA1�΅�9cZ��6!�)V�Xv3.d{���;Y�%��<��8���������@�/�i@��+Hl�I���:���y��Q���X\ܿ)N�y`��`̾qyub>ȃ���m`y Ҏ�!�F�M�%�k��R�;�����}�]J�}N#�ȥ�ś�A��G�@>�>�s�nɰ��Z_ĩ��{�<�EpƯ�q-ɬ�j�"���;�T��V[�[9K�l�\��C�ik<gu�"9�K[�Q�U�Y��$��S�-~ϓ(����yA�X�:�Bc�};�t��s�@�˫���J�Zf`��>��Q)�_f���#�~. �yU��ԟG�}�c���m}`�s�[��^��6vf�'8Q��[<���qm�|�������c�E���3k�.�����y�=qн�%�f;��i�ֵ�(��mz�k����ؕ�w\(�e��]tNr�񄚼�����,�pG��ia����O� 
!�S&��v�'7�h5/��)N�)���i^jŗ���O��ρ9 [�	1F�h���o��S���������[u�U�i2�5ԛ�jxHNno��L�0��r����J�����㷫B��/�YDܕ+�>,��Z(��oK�A��5�%uؖb��g�F�� ��0�~���;�����<B���4a&�z
�tN=	�!@���丣Q^jF�ޤ�v�6U��|vM#J!�xE�B	}�n0.��[ �2�۰L��UR*��ľ!�{�������0��T�D�d����(�Ě-E�j"]c#a�+����=���eDC���<MrFK��w�&�[�ߊI��V�u� n�KKq@D���9�����ə�[���vL�J<�#!Q�7�W[Ԫ��Ӥ� ��)4eu�%�t��`�6vdXCs�UZ`�c�Sf-sfu�F�.���4��������L�#�5��a�xŰƖEs.-�C���p�#%W�v�]Dqth.�-%��KJ�����Q���v�������g<?�h�\��ό�B>7����E��$7�f��2�x�wt�+z�ci���Y���-Js��?
C�7#i��g�<�����p�p�����;�:KD���x�W�G���ݖx���#{;"c�9(}��n@ �zm<�Rl���{/�=q!K�ke��@��= .j럆���b9h������l�Rk;�x�\G=�J')qda<��c����^1�� �rY�H�*��B�gL0S2c�iۿM�M6G���}�c�
�^OIa`��3�� �"��b�0�b��"ū#p����~20u#��7Ɋ�^C2ؐYu��j���%��%���ćmW�:l�as��O���vh{[�%/c��8o��(Ga#��? ad�n!xvÇ
����m�B�Lw|f-������MM�b��ӗ�ɀb��Lg�8n���r�Lg+K�B��?�0f�T���BQ@�z��2c��)W�Ǉ#�rWȑ���Aˑ�M��/M?v�a���c��ϓ����;A�&����󖴭7i�p���G�Y˳0iRC��b�7Tc��kA�Hȑu��������V�M����9�cϚj�;�3k���Ǻ{u�B�$QO��w�{s8x\�j6���Y^�vb��U��`��A;a�;MK���|Z$�4.0� �����`䅢���y�ݓ��r�H��u������-��E�C�2FZ|s�jgD���2���&+�ZC�=S�9='I��|� �I�⯌�Np#b,��'�
8A��v��&�&�o�M��S��63y�zF78�)��o����47.u'�<*�?������L�&���|��S�U~Z�I暜38�m>��T",�� }�i&)H�k=Ћ���~/.��+d��ZH(lM��S���8V�����W��ű���*�AY��=�ݠIG�!NVOO`�)��#R�tO�"��Ij��� 87( �]~Ҭ^$��h2�Dc͕���X�����ގ!!��� a�d�|��F2��0��P/�DK�j-;g����u�D��4�\9�P2�e�"�������90����K�lD�<>p�Rc'v��[��@�.� �����v�8�s �2�n�δ�`��_0B��u͕3�t[��I���>A�������Hfbcb/n��m�E7���<Qr.�%X�C��i>X�������p����H����̊�|0G��`k��.޽Oy��\eK�F�k���Ba�׼���5vM<
-�tT��N��["y��ðU\r��0�;vG7p��y��Ǭx��o0[���x�~�d&����!O�w�\�\ N�͹W+�R�2d��.����>t�x��b��Q���Z/E�|a���v�Ѭ�� �Z���n��j�dcTW�~�rbV��Bg-������$V�Ȝ�lP�c����\����L�L���oɩ<���_#^I���3�j�l�4��h�� Qεm��������̕�ux)EM�?���z+�'ى�$�,�'-d|�e+�X�c�]N������R���M�C�i0�1��l�^�n _�|�.��@����'��P�4d\%��X���G��]����:_��u���h�S˥�l-���r���c�|�H���
��Mz�� �Ox/��;��b����D
Dj6Q��������SpH�<��dw��򇂟��)�����i�/+�s
����W��_?_ &M�H&�����hkA4��@g�P����p�Z�(v�� "��7�gC�������T^�_��rF)?��D{ϑ��]C�EU|����,�����/8��/ �Ƕ�-g?���!�eu��c������55tK�W�%uX�Eeu0֫��W�ы4���r~�n�0ő��(^9�ϞR
�喱nQ$�A�ò��&;��Qi����#�7�_��aGaD���4wݻ�NŔb��_�qò����>��g?��A;qm���K�D/]�i��H�e�Th�Ll�ct[���"��e�KЎ���pkA��1H�*�!Z9�3��^*�\���\	6�肞�Au"�2���&��R��p�8�}���S�r����NcH�3.�ة�X�é��O9M��cM��`����0�o�)O�'X�]ٱjL������n�{�#'�<���ơvE$�5
5�n$����UQ޾Y�.I&��]$*�G����?z���PV�#�����.�;���岱Y��b	��m�yAx0���$/�XH1D2�a �=C���f�j�c�-4�uDFZ`�r=uO�ƨ���U	z�9�>=_ν=���.E؟���_#�
K�-A��u}U���?Ҏh���� ����5`�[T!�^p�����Ѝ�WZlR��7���ȟ*l�ׁp�����A��l�v_2t�-�t1��x�?)��9Lx�ia���Q�.�=VQ4�?�D"����2��&��H��%�N�q�n����,��7peO����Ɇ?���R��;��ڭb�㖕C�7�Y�!>҉o��U����/i."[�H4�;.N�	df��* iPa2��X�Tfo���I�3!s���se��*��Hu^�*�z�����\E\��R�8���
2|0S�k�dK�X���~r�eyQL-�Q�>��k� ���v��u�T"�m��C�&�3#���!�%��&#2�D��6q�ۮI���M��4�[BT鱴�>��O\ E��W*[��_vAT�/6�P��v։I���Κ6���Wj����Tr�*4G��%�=�CPXp �ZR�,��b������}g���H)���QR���S[6��6���4�4��3ySL'=$�R$����q�٥�}ģ�����n@��>pI�ﮱ.HŌC��� G���Hk1�(�1��B�c��q�J3��2��{J��JnD��dY��t�Vaӟ�V�D��3w
x��Ti�]�ķM��|���6�!��6�2>�nM�<�k��>w5֭xŦ��O�e�Q�,���Ә:;�>��x��B2���CN�Z7J71>�-L�"m"~6��4�L� �c#���,%U}b�޾�[�r�0��Nz����
�����������yy�j}�i1���Ѯ���^Z"YŬ�]Ho\���;cЄ�oL�Ŵ�l�TٲB����&��pҹ�F<��>��U��1�<s*'���塟� ��a�	��X"л� ~�ʴZboE����|���/�j�m3��9&����:�)�T?�H�x3f}E�Xziw���Q}��k{Lq��85Դ�&��i�����g�F&ڬ`�''���ߟ����\TT{_M����� ʯ�G�y(��w�aoզ�k|~�Bz��C�F@]��h3��kE��) ��.���Q�c����&e����I#	������pf��#���Z���6���o[��3�C2
nV]��	�V���w6	R����5�7����,ō���y����#C"���gB�Y}�J�b߯�Ҝ�Cؑ�J��g�[��PV�7J#T�@�U�J$�����ʘ��
�t��f�5������(m��d������ű�t@�:��DV���
g�u��|�/�j2!�R�AA�3h�g=;�bz���� ���U�l��6�+�.`��@�a���eM(I�Y"6N�P��Gp>7��!/�<ȯ��̆���,������
b'��/������S��L�Z\&�~����E��t���ay�M2w��#^��
2��Vt�W��}�A��=>�� و'��a� ̈�����NL������-�Ǳ�$�/�ǃw
h�)1z;��.Zj�������U���m�d�<X���X�����&�!s�:�<�F�J�+N�Ra��q��	�����Y�R�T	J�B���h���+�����ޚ&3MP��1f�m-���DW��(���Ϡ�wߧ+h^��l��p�R����L򢸑��?����]��ax+�<a,&bz��>�7���J��dҫ�A�qw>��b�a��&�i==���}s�|ȩ�ۻmDR㣯�ί���ؐ�n�^�9�I�bǅ��B�:��7�c\���]!I,��,�Q�m��Õ�_����[ɂ���x$�N,��H����	�T��P�E��1����˾5:�lr�#�K����1c0-9�n3���:{�~۸�Dge���7�q���N��Ӊ�h��Q�ƓT�I��Px���oB�I���$L�pX�nƮ����6;s�k_M(3��2�^�'��l���0�OrN���Lay�`����9�N|�O���R���e��H6����Â}Ө��S��Ǐ���x��bs=�Y��HK�x�7,QP�����	u8P2X�z�
F�9�m�� �6��o[��sύg�y���N���N��}�b?.Uj��L�C��>�����r�a�}��{]U�N�Ȕ=&G����@�����"6���GDE'��8��w�=�c�T��cV�UɏA,(~>p��W�\��c5z���ۋ���@i���qy{����������.:�� ���.���9;���0��h&���]ʃ�I}�bfDfyJ� ���h4��V�]Θq>�Y�~��n,�N����N��m�
J��N��1L��O|f���9Uݚ����Q�w�0v�vF�XK�-��A���F���1�c�ȝ�XR\��'����	���Y!I��$>�@�-�]Yl`�:�̊+�Ǜ�P��㜩/Iu_5���2jfש�kX[����b�82��q� f�m�z��.���uho>$}8�����1��񏋿C��&^)'� fB�Z$R��c#<qxQ�c@��nME��V����G��I�B g�V��$���ƽ4�'	�V$Y��3�P�"��0?;.��Ȏ`��`��[�X�ogR�G��EeX�&�/���W�M�a��~b����wR���\`pX��R���zx��BM,����V��_1��	遂�G��̓mC&u˱%6ʧa�ؐ�.V�K[`��������в�haP8����d����v�djDG�X�E�:�G,�%w1$x�EO,u/=sl轳�H�5�brРW�����'m�>[�xOc'�d����F����T��'������X �	n����8b�Å��D�xv�&��'@�(��m��*I�������60��;/h�L�E�_M�c��W�����ɤ���@LK�Яm��\���SK��vB��M���(�pAM8��ڿւo���}ރ�rӦ��u��Ȥ��lE~��y���x�Dѷȏ�i�b�dy��u���&��浂w�,��f���L�x��k
�$E/B�K��e$���t��X�ҭ#����� � U�븄��Ϣ����a�WȖ�E����+hէT�>nJ*���+�a�Fz��ё�r�͠T��h/�!i&d΃.����i����,��v������#��lu�SN���r�jG����5W�Ǔ��ot%1��L�Q�L��i���SŅ�x�T&���"h��CyAɫc癩[��3��!�HH�hH�[*P���*�Hy�Ř��s�V�@Ѧ��NMc���'�c{_�(}��(X�5�#c��_><�l5�Oc�w�9\TP��7Z�|�(��:����#y ]�!�9]W�◛��4G�
3U�Iv��I&j�؃Mk U	<��^�lMLg0��;��
��dӁ��D�8��$o!���F=ڎ�� %8_0���39
k����������,Y���&iJ8����9E^�ɬ�EA	�P�|U�7Ңާ��q�X�_�S�8w[h�V���fq&��N ��V�G^����➥6g\�����J���(�	_��n0y7������M���kD��]e��b����peW~u7؊Gw�;���#Ǳlm�<YtaܔV�d����x�"~)�����5�ϥ�ٰ��ܙLN��q ���:���]A���XUa�U<�����J�) }�8���)���������x�Y��/+lz�f\}נ	�>���;���1��O��[��՚r�G@���3����Tڳ��S��ָP��XQ�wJ�QQ��_ jW�\'^��cb���3�ۍ=�źk�toP#썂�HtqOv c��Du�ͼP��B�}oKঙWx�_�1�5�g�6y%7��#%�(�ڹ�K٣�ߢL�C��Q�ѯ+�ݪ��v�X�9w7��������P��t��l�O��h�����K���sw��;l���f	��'������o0�'��u7%��3E q�%��8�c����H��V�U�������&�)7�!`q�� v��*,�K��C����1�+�j(�j�Il+�Il��Yң0�m,d�X�@�I僺:�ऻ�:�w�����&�q�?<2�����I���=�G@q92H�↵-��ðM	@y�
[�n��"�P�jPD��f֓jD2�6x,��'&���r4����8��\��tB���o:�$5s��#J�� +��j^��^/��gC�设Ǔ{��^� �We�z�y_	I��7�h�;}�~hUDm�NiY`~&[lV]��'�F����Z�GQS�K�~S _N`D,�	����0i����m�2�@�{C��k���ku&����1X�\0a�7p���m�����#���hur"��&\߉j0�@+x�J��6�0�M�)��C{U�	G-�F�'bw<U����ڪ��q��kIO*��o%��q;�����syA�-]�bgI:� S���CJ;���Z�X"�Nr���	�$YA7�(�Ԟ-����5�Hz*�Ŷ��D��zTDF�[��g�����9�T:e�X_$�Zou<v|k�霈��{2$�C}��Ϻ�X��hcb��T�N�"8�7�^u�m�	�������թ��2�ߍ
���Wj�;R�.��e����,F�ܖ��=]|e[��6����:+9�8��$���ĺ¼���ڥT�o��:��(����@�$�@{�e�硏�a����g^�����UD'��͡�(XTPO+���0��S��@/,c�����`�xx��6Fh��*ͱ�$fgi�{�
W��[�\�Љ�at��W@�Dł9�c(N1�P*\�D5��O��o�7Tt�u}�6̺�w�i�$��(��1����/�>�-��CK�(����p�~e��"�̻�TY�Č=�h{.7�@�K�B^�$Z�nR�V������p�P$L���h����C�{�A�
��L�H�8�l����`b��dh����x�����y�W�t��!x��;��
q���#�)f������*�z��϶E9�Q)�|9�	�٢fHA%/�sثd*G�����A`��sEf�A�n����21��I�B�Ju�l2k�z��$d�&cb�%�G���u4	���+)���u�2۳�z����)�#`$�\6Y	��a���JF��>�����^D����z`��ĵ	�7��]]�����Z�wY�skqT�s��t��]qwӐG��� @�*"Ҥ8h����K���$�K�)�)a��R���WgPt-
��C&.�z
��䭸��*�U�I(>!
dƬ�����ǜY��ei����@[
��6ˁC.�b��Р�\΁�PܸO�	���W��i`;������b�v���v��?TQ�=����dX~���ќ4!6N��G�`���yD�;�v���rh�+�����z�q���@q�i;n��UO��.��ԓ��:�߀X<�?�96�_�E�d�*��HY��+`�ɮn�=n��!�'svNF�= I�|�4�LG�J4�܈��sN;j�Wer�ȳ�4H��0��`�����֦$1�l(���*Xiͧ�ͅA�h��@�\����BX~�uW�>���������2ۘ��-�3�y�5ާ�v@7��Q�&����D�"2�6�q���ZCu�4:E�6z`�߆��s6�.�Bfh�
 ��RU���.}���S'#�XCL�J�mt�$[$�0�5�����d�J�z�m�0T���E/��00��w����~��R�K9��.�c=��7�	O�*��N�R�o_��.ǣ���
i�=F���ܧ��w%>����7ґ:6n���H��ʘ�͕I�̞�_}3%	`0���M4V���~�5����Y�=i��޹�(؎s��m�hg/��)���mz<����QgQX^DQ�V[�Ϊ���Xv8u��8�ƺA����+8%2�ɉ	���u��󊏜��0�b)�#��z����T���	��P�d����`�|$�j�\�P5j��r���K�U �N~���m�X�x=���W�+����U���'r=�f���W�navf�v�D��Hs?�j�O�*���7��X ������u�v����60�h��^����Ĵ�	�2��S���f�X+p+�#�6%����ţ��6��.mi�y�����q��8'S�v���ߑnw
)1�^|�%DB��%|6�V���b�m��)�:���.7I�y�:HUFIP{���)�����4�n	W!'ߓ%�_b�3�^[�[!ic��-e�J8��&���\�>�hl*Y���Vh~���R;L��/_��#Wݹ�O��4����t�`l�v<�&%�l{O��$��|��B{S��`f��S��>݉V�! T�@j�{�2���K�$�d��m�<M�R)<����W�Z�a@#j-K1�0⬱(`����j6���rI�puS�:�3��ne"�-��d�j�mq(�����!���+U�z�J��K�_r�o�1��\��P�kZ O��������L1ܺn��B)#�5����9����j�3�o�C[�N~O媞9_��A�X����1���Nb�{�d�� ��u<�ʘUՠٜ^<fw�! ƾ��|0�N�4@෦)	�8ҹ�֪op�^��Y�#��|�]�N�.8+׋�j�2�W}`����7�N;�j2:_�� ��r �ҐG(Q�CG�D���J`������r΄��ߵ���.�^ã�	�.����at.r��N�?��B�ht��$=��y
���*�N���fRD���H�qF��=nHL�M�4��8��>2?R�	s�c�_��fU���}�W��+�m]�F��	�o���Ѵ+�H��JL?vuP��L�m5L��m�U?�-�hM%�+�Y���=B;��F
L.�ב�Ĕx��Q��̚�D�x��B�>]e��2��1eL�
�VH�>>9n`dS�X�s���bt8k�jbX�԰���j�N�WY�=��Á��W�o�:Oi��5�Lw7^+���<Hn����[s��Aj��ej�vHp%��H4����D�X�e�\�Ê�>�����K�����<��d���z�k1��G�gG�غ?��#��Wg��ͼ�!�^a9���|�&�S�a*~��$���V����v��V����>�W�B�U�[�L�a��>�A��2�ׄ�����ߓ�J&7��C� t���b(j���i�-rtm�n��'�P}zN%�k�{��c�i�e�9f��sZ z��	��\k7i��/�#!�k����n���3��>�|TB��r=3ߋ['��/顰tIm�P�X
n���%���Z��lg�(�wJ��+��A=�)>�V)�9���8t'��C� ~`�/jD���)�U�7����[N���=��1�*$v֎VJ�e=�wX���B�������Vd�����F��Ue�Jm18�AC�(@�F�����ή�������)]�vs��]C��x�XC�ȩN�[�A���<��p���B��w��e��!wrdN���a
� ��g�����,x�~G�5=c�I���b#A̔�k1'&�]�UX.K;>�׈�,sy�ָT/��8�ہ��}�>��>9���W�^����(-`��%��B-�L�7�D_�-'��xW�[[UJ�x�_�h���)UӳJ�Œ�mv<�{殖_^_<*=�P��զ��E<(3?�ś�V��{���8hQ�����l�e�uthp���&d��K��\3L�;����4=x��9i� |�b�G\�Ƽw�=H�,:�I,S0 4֙sA��B^r��T���`���,��84{�n!���\�;���{�&is*mfl��~���2��<4��B2��`��j`�S��ɰ�����O뜰�A��/O{:�T����<TV����*L�Aa1ua���!��kx��jƻ��e@̧��M��r(+�xG���P�ͥv���z��3���9�Y$8Z&$�;�Mؕ�~8��cT�v��Cj"!z�u$G:o�k."��,ªP��qZa�Yk��l�b����a7��`�Y���C��"�����'|>��z��A�-����;�u�Vc�D���Q���;	�k�=�J������g�K��;UUV6�ۑ����nz~��k�t�i��*،zc�o@Z�R�cQ��!R���n6��z��1͕��R����W)/��%k��I�����$����\�P�l�3-[v5nu-�}I�?~�Z
 �a��jUF��0j_�p�yfHIr%����iYٖ;��[U-JG�� ���(�(�|k��Σ�r%^��ЋQ$-��'�Eܐq�4��L7LH\�q���T��M�*_X3�/A��&\m��죆���n:?i�7�v-�����3��{,���X��@����u��3��]�؟�b�	�3��%��L+]?�'�쮧���p1t�����+h�� /�2}Ҷa�F����=����E8�$���%�oF����0�S�D�f�S�3	+��	#�9-<��cĳ@�6�D�3� �P&����M��UA����#��(ɳ.�e�a��h-*�C�zd���X+��g�_t>�;�����i�����	J���ⷵ�s�=$zQ��7h�$9�MIm�Ē�	�U��^=(������	�{`�*Q:�o,�R�����	�M35���t��V�S�)?4��Z�b�� �hۋ;���l�������|���M��Z�n]E����^A�a���o�b��0�d�j�{O�� ��9�i�a4��lW�StuW�K�)UҰ��qL�=w�(�m��T��mʠ	H�ֽ
92�{�'s���Y�2��t/�34�U��j�7'>S@,&�Th��kk�7�=*a�SULh"�FU[�@N��nck��R%����x����>�Ջ��M,��i�d�Ϙ�������H�x��C��yau{zF�y3���͊����r�.P���&��H���9l��̽'��"�#U���ZDc­蒮@D����(��M���U�/*�!���;�����67Q�\�8���^̼��ԡ�s�Q��I [�f�Tq-�N�ɣ�������(��<�a�3rH���/Z��A���)�������#6�3n4�}��(3����
+�H�M�i��!�>,������M� ���:e<� ���_Z�&�xg5�$X�4�ȅ16{eZ	��W��曠�WX�K@ߙaw���r�K-\�Yi����'��f��ɇ�	��m�o��� ��#��D�y ����+�~LD���$>�Z�ј�$�v��<ZV%6i��O^ n��X�гc!.S��B7�����;'�ta<��a܌c\���^">dQ ��Q��| ;|+��Q�GO����!���AHTx�AʿA[JxG�,K���T,�p8Q����a�ܭY�]-1ϥ�<�j�IUCG��g��n)��K�%�MD���8���Y�o�R��V��j���]�gj�	����ZI�M��k�#��9 m�>'��s��/�bg��
�#X^����E��hS^1f�B�Km�o��sU�`h7=!.!�e_�Ǵ�׬�ӵs�hݻ����H\ Qʹ�S1�F��>w�u馁p�f.Q�!X�����L�z�U�<�A<��?Y�ó�@?&���@�ƹ(Q�2+��ˋ��]��5�`����XO7U�7[]��I
��a�Ϟ	���`q�#����ᠹ%�(�O/}F-X�ֽ��^�9��=��� j����CR~�t���Fg�b��}M�Z�;>�+��6���4�?���R#������-dJX��7��Cn�j��h"�%�0�'?	����	sa1�W�oF��e�=��̏�h<��f�M�����|S39ԻU�؞������C��>�e�E���먤E�(A�{����c�5TG�z��� ���|>Z�����T``0Q�����)P�ҽx�O?��"�w75���%l.�7���><�u}Fڇ������b0�*��ʼt�H����1` ��?��[���j�����~mY��p�{�yy_���{�=�;�K���{p���p�ˎ���c��M�X�-pE�i�nl�y�B���(Xpլ�Z����l4�ryA�nr�28�;"7I>���J�Y%�̥��s�[nY@��;1V?�ۍ�L����P�.XC��3��mͫ�Խ��5]��$���.B8�}�MW�d�rՍpp�z!؜rIצ�_%�.�g���\g�)�D鱝��^jhq��bRB��aN�s�O��-��{y֮���f�)�
Nx��?��m!gVL���K��mk;Y�DW�6�_��j��eܠ_��B>�Ph�4�b?0p��!ǟ�3�5��m�1>A�3�	��w�~'t�T.c&�ћ�kW?��L��{�Dl��3UDow�<K�@o�Q �=	�q��K�[8����e��K��V��xbX����e.e��85 A?:�1�J��S�Y:��i�&+<(a��C@PY�)���:j�]תe�d�q�4���.S:�.�njB�2���[T�.��Y:��re���8I�˧����U�'���t�:{��Y1��\O(J`c-Z�l�KWf8Х�VƄV_Y��m������t�My��i���'3�KQ�I�d�H�~
hS˘L�E���S W�3��n����}���2)@�\�O�u }A��
��do~9|G�#�u��r��L�pV�+�=�iW�x�<�/�~���e�̇�)'���~æ�z�'fČ��Pb�^���Zx��s�=[G�G�d��oՐTq���b/~�*~�+�u�� 6�b��"��*��M��T7T0���
6 o�_JBh���A��?N�"�?��I�@�J|Nd�s���/]�׭[���{ �.���Jͩ��������8og��s?!�IF�$���吊fW�\h	kh��Ko�Ugb�n�Z��0K8?��6�V0rs�N��dW<Dm��`�9ZݶI��T���>�M�@�淔� g��bmw�T/�9�m|�AN�8g+qŲ�t��cY�'
N��'en�>vɷ'[/M  ��q�2�a9�zV9�V�r��E���%ts�!�i��n}jڱl&�yJ�,"�}��4�SHgm�d��������W߻AP#��Zp��u#>�6RƔ{�1��p�"�V�!���a� ӷ&��7[T�/�-f����ptX�W�@��=)�����m����.�O.x�%��t�v7X�'
��j؂��Rom=nR��u� �2VcKG*��tЌ���kE�B�F�Bť�;��>3���@���-��e��NuR�*���^~$���H�a�-�Y�Wޯ�f��<���mS��8��9��q�����U�pRH0"�&I���ZQ�*+�����?��@l�V�pJ�����NB�g��o�/6 !,e��H��Pƛ�'ru����'��&&������*b��f�|���{���m�׆�F����8���ND<-k���n>�^���sG%������L���$��O�m;Vxx����Vx٧�����.��S:,��>@Tƙ�3.�U���壛˥�^C2�#���S�K:�_�Ate1ґA���m�����^L���u�-����ғ;~&�Y|;D�z�qEH�P��>�O��e8��Э���D�ʤQO=�٩�;�j��f)��C���p{��2�~B�5J1�ݸ��`��6C����h��i�����\�(n�:SLi�Y9De��>)������������$��Lb�ߖ�����9����D�0�m7%��h��#�PX2db�BIb��o�8�qb�b`�$��r�(��z�g'`�]B�Fu<u��Dr������1���6[m��D�m�kغ�����(M!;n�T��)'h����XS2f�Ȅ?��'l����j�&��y`��c����>W��{����S�TF�sM��D$�1���@A��v6���G/��Ρ���=�q�~&T�����.u\R��HB_2���i�3`���T(�_�ކ���Z��Sn�1�++�����Jͽ��EI�W�r,�*����$�!o��T���ϒv�[sf�.��4�78q[��StK�}ä�o����OH#>��pM8 !��ܽ���] m�2i�?���v,s@Q*���=v�������6b�O�Y(�_��&�K+��:��8[�����YЙ���[���T�X����Lf��%�Q�'�ilɗ��R���A(%F�dt��g�l��k��������5���K�0�>&3�.Hc�(5a׶&[�U�aPi�Z�V۶�N� ?�K$Ẕ���0��}^m���Fn�$Vfﱕ.��O�R��W�V;��W��)��:��$}�`f�[mj��4�L�)p�e!�I;�Kw1�����O��-�l�|��ݍ�{��#����@����I��e��h4�W@g߽�U��U<M$�X2d���Zg��!�S��ЦH��x���8|L��x�s��v������2O�N�/[���O��}�
	�n?L�U�k����v7��H�2���ˈ�{{˖4wޝ�겅m�.ӷ�iǑ����D�_�G���Uh��딖Ҳ�Tק۸�Pc�l+��6S���A��X��O�������js�G���`R�W@��%;��1�/b|��Cg���P�����Ev�F�yQ���=9k��e;'���]�@�K`�t����7�7�/>T��{�]���3�9bFc� �b��7;�#�U�Z����ӹd��*.R� �Q�E����y��R�����e�4Se$��ڻ��'?��;�)<�z;������d��]oJ��Z��`�%�~�ol�r���b?���P�-�ώ�G%@��kcZ���MMV�9�,μ"��7�~1��s×���:%�q%�Ɵ�=�ka(u]Fp|ɬ��f��T0-p3O_�a2���n�]���"t�������D��E�[�$Z�:/?��� \QHk��~�s��Oa�ς���	�ٜ�=4׫rl�)d�O��y�����DF��9G�(|�I�&1P�a�)�?�k���P�ALȡ�Jk��n��(oM��o�BhBli��-�����=I_3*z2�v�-�y̳�������#76�vu�˙�:��C���E���&e~]�

����w!8�����{Y)&a�-�x�"���rk��&��Fnq�5M�Q�D�����5�J�� G[�6���/8��JO"��Y�snon�dX�v�*��EF�^	�FW��!�Utpw�z�e�Qv�Or���w�}ݦI�s����*��~(�o�
�X����cͲ�����ࣈ@���)�L��֎Ŷ���p �{ƍ�<>����2k'��!�����`��s�ҢoLOm�G[\E͋��`�n��T[�H<�`����v4M���m�LJ��K�l�X���!D]�<&>!��\�p�&n34��G�����Z�K��r:��������:%@� �: \A��#{W�a�
UN�����\6�j�
{d!����Fo`t_cUM�2�RBu�m�nԼZ|�Y~��f~<2(�������a/�iG�g`|	SX��8 ;�,�_�b�?���U$�ə+h�$?�4�-�(lnu�J@��!-I���C{⿎]�!p4d�-����H���#ϫ��Rc����В�r��m/�

BI4G1izy�����F�ک�	����	4_��'�jv*&��E<��q�N�"ߒI������-�ʖz���Od�3_	�qj������Z<*�B�Eac`!}ʔ�d�6'�E�� �����Y�L�YP<��;~i�KK�,`&{�)72��b9A#1/H1	m�}����̮:�/�}8p��Ң�Y���3�Myэ�-"*��	eֶ���U&P{�j������7Ki<���Q�G���x������3@|��>z<��"�ڶ%�F�C�a4`|���V����~"T��U:����t+g�n��}����[Eo��;4��e�wސ1�P:݃^�"r�:^Ш�RW��B�M�ǖ��s2�PJWJ>��PU���HGx���r����A"L�+0���р4�M�wTZc[��ݶ4����;Ҷ1�(H9OZ�m�V%�z�0����wᕃ=���z[r^��(Y"���S?���_�_s	����'$����������Lzݼl�p����r����V��f���Ԑ��o�����i�7��/�>���w�ϧ��n~�"��'��`�,����U�;^���T��5����*���}��ƪ��Y]"-n%����"@�(��T�X~��J���B狻��b�+yzɏ��j���X���>�/:(5�z P����v�E���[�5A�ףϫ� ���E4��*V�a�6�͝-	�(rtc�da����"*S�%�I
�ہ���f��|+�/�'ѥ�4�?��m�"�q8�ZT���F�r΋�'�Mɂy�%�V���N�&^����Y(fP�9�BXr#��Vjz(����J�D�J����r�!�]ea�5��}S��:�D� N�\.gn�´����h����HQ�E�O�,Ȩ\9�g�5S�U�Y	w��� ]@�P�3����0����돩�x��z�H�����C���߁:����m�N���P��!/�c���vruf����$B��[� �W��A�����k(�Yx+���U�������S��FBI�R��Y�b�̱$ �b��^���)g�'@�s����q5P�ZTw�S˓�.)"��8�Lac0F�>�E�	�oS�sM���zn{%�_odtjs��vF�g_�/s)��<s8��'�9�n@AҭΞ�;�Z�4[1s�5���t�Eb{�;O�Q}��D���~��H�z87P5T NZR��߂w��W��lC���uw�����uM�n�	��4�U?��5�V�����8��*�� �`}����l��BVpN�n4��tw�%���XGL����[gz����F`���A��7v���r�Dz���|��;��l�a:7`�B�t�.ue�	A���&�fᐫ�6�6u��n�	����R�����G}�����s8��Vᇂ�a���d[*��q1�h}=���ɼ�����tn�g2�^l'*�����,�E�+ׅ��#t��G��������^e��F?俇�7HoJý��Ӝ
��������qf��}rdҹ���ȇ0��t��!.>���j_�.ک�N
���`���J.{��Σ�B���Dv$���>�;�y��ūZ�>+,x�O8�9�" 4�.B&8�6�E=�Jʲ�^-C2$E�JE�d7r#����>b��-�`��Ũ�cJ�;�|�k��v}�:�4w��d$��	���\�{R�k�6��h�*��C��䝑�T���M�F�Z$_�j:�KR�U����ϣ?b�UMr���T�{d��s�7&9t��i��B7�yLm��d(o-�"�y��C[q��In���\}���4��k5|&{��O�0��,q��/$��%��wA�4�r: �)@����H_
7t���Y���I��F�x�3U{���6`~�k>S2+qgѭ� �vDa���3�/�Y��
o�(�����J�E0E�1���"�H���Oj`-vJ׊\��u9�?�0W`�\��]E2	�h���ǿQ�O"uA�0�P�ڿ4k�q��]�]ܸ�-����4�O�f�C���_�[���g�YI9�O����P��#��q��k!��'��&�Lk6�7���{^�Z����*@�5%Y=��b�P��z�Nm���B�1[&�	�f��E@��+������ĖJ��b���ۆW��[%��v�h�&�����Q>|4��j4�톬&�8[c�@�it]�	�yiv�.v��bj$��,�+#T;r�5�l��t��ӻ��IX�����r�
9�3��"�Np��=�
e��-;�6�	����oQB�S��`{�#v~#�ͮm��'5i���X@8�9j�� �:�ρ�C�n<L�Nc1g�ⴢ����H�(���g���c�wba��S����Ik�&��%@�>O�8���~��V�8.�E+�~��Q뀷�������e���v+����E�I&���n��wu���r����ug�T�
�$4*z�E�=U���"��I�eA�_q4�0�.g����(�*�U-t(��K'#�)Ŀ.Z���s�9�N�4��'��;�y��*a�\
�8��6�������51���}T09a
T�VH�2�s<��_�#��Nk���M��I>���ܐ��_�KHkMUo@�W�]"t�����͠�4O��� #S��9Χo�.��O|W�J���n5�gG;����l����_`�qrO�E|t�BDp�O�a���|�A�I��	R�?��*
�g�@D��b� -�,��[s(��\�}�5��xVr ��HMH��:QV��X��w�{�m���C�r�bߓ�/��xS��Y��U:C;��h�����7�4�]�?$)GR�U��ɘ��<���B	��qi�d�$��s�n��Wq0�6�'�!�M�)-���ɐ��Q72ٟ@��E�J�iBE��S"愯:��N#	x��p�6��1��+5������-���L������z����j(�g�Ѥ��'�X8HU$o�^�G�r���t�K��>�t����^cT�mwe�A
�pP��5�f��y��f��Ar��ƹ��	R��4�T4�< �� d���������|
˝���ⓩV�qd��x�cF�L��bű�Ը��B�;��%5��#����~�ظ�X�ɳ�Sp��є��μɞtDZi���,��D{(^���f�+�`�A�44�T.p�u�����L���T>�JH��~q�(N�������ͳ���C����g0��Ιϊ�<�d�:��ˣiQ�)1UeX���yH�D[�l�u��֍)��=�s�tZ@����)�E�p=e}���9����-�S���<l��L�Jt����Ԭr5�Dn��2'ؑ0*�#;%�:_x�z@-4u͏(h(I��ja�Օ����X��c��2b��LQ|�K?�W��Û�2EƐ�:@��fi�AC�iM�P�5�K0��MQ�\� �ĉ�|�=!" *�G�t��ƫ�=`�+J��ss��./bke��A*�^h#�B���+����|G��-> t��� 7~*Q�F���]�< �.���U�9�W���T�[�S���y�J�.g9�#�'�
��=paOn�z��$�_K����	'h��4���x��<s�;�Z:�� �[������=y�Q�Uk2�&�b��}@��L�;��wj��f7�[��Υ�.��50M#����!�$c�Ϗ�{�`�zko���h �/�߳�~���|h퓢�(�>�Ѥ�OJ�Ϋ��vvv���7���hK�I�j��e��%�1]#k�: -�#���p�Ϟ�Ƀ�\T�ݮ���mCg8#�w�`}�ī]�t��,*�٥x�-�z*wb�p�{���n��{IU6M�@�2»&ڸ<��@jeTP���&�2F+��b�K��Q�uԓ�	/���ƨ%���lכ$q�)�0:4V�oau�md��J7���Sp�L���Qy+*�U�,"�N��r:�}��c��8V�����0��;<I�C�l�\X��VV[�[���o4�]�����6���#�G�{�#Lx����y�����	y8^͡�_ܷ�q�Ka�L����3�^9
�щ�qU���4@c��$��t&xP<	�*�Rh�Y�.q��ˤN?�;>��ݏLl@��)SU�\���2�Y͛� ��;6+�%���g�Z�eov͉O#�96%���-5��uy��Ŋ�#0Aaɞ���MU?������'�2���ת�EC�z9�gya�}L*0,�3Dg�}�H�N㘧؊�n�pk�� g�6ᓧ�Ӏ\ѡv�p�n���r��nȤ��v�O2r^At����}۵�a�$>�2��S������V�����z;^	%ވ�a?]1y��g�k��ֳ�f�J�5a�rw�e >���x��^�}$�Y�"�qV���U~-#�-��O8\㵼X���kAf�HI8T
&��	�Z��<����v�<��q���in�+������]�Yߏ ���d6�#�կ
��N1��x�Uow}���,�a�]B	]��X�'�R�G⚭:~�ٓ���VGm��z�Ӗ/��= �B<W���r��HPxE��v��(�q��Tl�iqu�m���� �rU�h��4�\�=�۾\��fj��r�`�f�k��H���^�{h6ʬJ����_�T�bVu�ΰn��m�~�|�m����/]|��W����XE�|�+%@7����n�]�V���3���[klLj�m���tf��>gܚnr����H@$oYj���lU��|���dFS�E�=��¾x�Sҏ'	������/�w��E{-I�E>P䰄��� �/�(ϟяa7|�GS��J���.A��,G�`p�]�Ǌ���
��8�\����v,�����A��@�a_�(m
���[^�v��k3�g�������l�V�?�\j��$�����%�H2��c�@_���?yw� avA�����{j��T����L��` [�x"����}̺�<c��Wkwx�Z��o��x5�Z	�ɱ��/�YS�h}�C�q���k:��(JJ+��}2� iw�:o����oW�2��x^�콰SK����N�MA$�c��HHv���J�t�l�&�A�,~EG]<�OwÑp���$�+�4DD��h�HH���cp�e{|R��N�0t�cԵY��b]YB9���T�Kp�2��[G�'$��~!���WQ/��'=�e�A��<׹/��+�`�/ E1CR�C��P��wU	���o�rW�x��1ʹ����kY?�T��/@ROX���ri��8[��з	r�幒�#�}	<�v��v�K� �!��	����N\�?y`�����2X�u��89 �)���X�_�<1t��)Wa=O�a7�L�*��*Q���䩧�DZ��:I�V@����K��%��胔_�VCǍ���o�;�߆�����"m�\���᭦�c�-l�A�8r55x��ͬ,a�M~quXi�"�)���N����2u���8s(��3&�ڥ�x�/���W�ϸUD�=�����c��ֱ &��U�_�Y�C�c���3ũ'�b���!��)��s8���i��~/|9-�<Cb)�	C�z��ڷX-���MN~�s��Km.�33�V�f�o���qd��~�"��Xn�r�?.�/��ʰ��H �J �
y�~p?��}yvI9�D&��8�c��-=�<�!�\,V��o��m�dJ5�a2�Blywi�0���'aDi		rl�Fu��҄�-9\��z��q�c��08��Q�~a�&zrNA�(��Y�5B���l�]�/��hm߅���1���3�~�x:q�{h�X�Sr�� ���*�$���U��e���ײѸ��%�:d�����~TK�I����[��?�M͸q����zhX�����g��[�8��a:]6�f��ܝ���`T0�JP�����}�0�ٍs�u� t�q�c���/=d@�!�d~����$�_ĺť��a��=	o�A�H�~7�Y
��n')�(����������"�7 C3F9KSf� �B��s�\�� )��9C�1�ƣ��3���<u��ԥժ�1�(x9���ר�d��#��V��q�%��; 1*����)��Jv@D��u��_n
���ɉ�����oN�7��k�p@/ͤ_�	d��
Ϝ}"H	{-@2�4XX�`�R�����l3�J����Ӥ��]�2y� �}���ᶀ%L�C��C����Z���O /QT��+L�%��IV�庑��62d���j��坕�D�g<�WG��]�8~�ʔ�(O&��9�xn	�B�B
#��+􂩤������Z	닉��x���
)!�"����L_��k�4��N7�q�Í���I�ƃ��V.*E-�!�ä�����Ygq9��T*5'�+��1��W��4�ҫ�=�}ݍ�Zs������!��"�E�;Y������ /����BU��Ex�"G�D�	�|J�xD+�=�\�==]��A�0A�nV'\f��_�ά�j���;�\��h��ˬS��������_�J��vo�2u�Z�ٍU�#7R|=�^j�D>��͗o�������2�4h�+�U|�긮w��9��]���������HS���S؎L����m�9|뒀]T��.��=eW�s�s��%��Od�U:�8�y[�N�KU0q��c���b��j�V1.�biQ�f�V����nA����RtR���b�P<��|C�P�8�Y-R ���i5̔��κ2��y��OK`�茻��(�|�6I�����6�ư��<*�#��,�a{D���0�?w��S�wi ��) �I_��X��j�d�!�!�3sfZ�	�_�X�UH
O�-.ὄ�����rj�4�������K�uS�G�o7�&��7zX�C?�]���7��;6a)��K�p�_�+|'�ߠ o �:� F�ʮӲ*�q"�q'Vj�ɹװS:`ej�Q�]I��m�����af��pt8�k]n� D6`���	cD ����<��!MM���x^`�,�w�U�,�O4k�Ȇ�=���O/@`Ф@����Wytx-�f؎�m��̗Ί�S����K\�П��R]G���t6s��|�
p�����9�N�7�nJ%k��bڽ6�y�>ѹΙ�VE�?a3��]��d��|y�g"��T���?-��v��cW�W0A@���`w�<�cTve�}��p+XS_�"P_߆V�A�wtOc/p�3E'��Ze��_���Y�%�켛%�8��\��վ2 �w���S����ճ�$���Jʑ�+���g7�h���bǬRV����[�0|��yrG���vzFD�t�}z�ޓ( ���O��8�J�czۻ�%��o�-�����B��	��A��� �#����/%F�����H,���N*��7򋭳q�{���7��6�O���V{����|R�e�>�K����*��@:M�ퟁ���o��M�$罐ܢ]( Pjҹ$���K�G���C�|���\��_EzYp��0�	,�������ɴm
�F8��m�	�N���k�=tۋ��z����neQ˴h���#Q?�|n� �u��i�ɠ�.}�oP�&�:���Q�oz��=���g-�׻W��g+ �Y�E%�P��0s FXA�?��4��i��
�R$;�s��H��t��^��U̵�a(�e��GɃ��z�U�7|��J�d�K0+wRK� ��G�e��Y��Ml��!�2��9��L�4T��4�]�FF�;�f��S�ΰ�m �ϢZ� �g����������`�m�"�݋7#���{�">���/�P��󂝬��mE��k�j&J��"d��]<��	OQ`+�B|���
�	������
���<�3Y��{;<��/�����=�2Tv�q��+�s�����/ZP9l�p:2&N	ߋ�������f�l�1�M]�2f�!5hfQ��+r*�nC��ő�NB{��,+���B���ϡ� T}��#
�f��`��w�y�>�R��5�Շj�������O����sI�&�z@(�M�~
��-������wL#�L�1m��~8d/n���</��A���ł���NS��f�Y���\�+�Dl,�Q�ٍ�tV� o�ߝxЮ�8�r�fy�����U*�S�E�W�PT�8��B$,������K�"r/)�f.ˋB���#TZ`�POAk"C�YT����GwKA�dHM��#���d��r�WK�i21&Q�J�Y��7����ļ��6�V�:�@e��A=�tY=*I,:�yI�G��Тgj¡KV�DυF"e��A���H5AM�~�-�
qxd?���ݶ�Ή	e��0�!��F��	cUA�AL�[�� �螯�'��Mr��6?����K�e��5�^���W�ҭQ5��=�	�o:-�>#=.3��B�G}�����qJi��<?:?Ky\��4v\V��T���c]���N�ߥ�zZ�p��	���n�������J�H=�D�'B���7�lC��l�r�D T��0H!l�)�3��i�w�/1 �v�� ~�(���37�3�l�ҩ�� �w�?�5S�j���`ǹT�Y�0�\zS7��
���I�?Y��cH�'�[(�	��h���MFP��YK>:���Pzi�Ɇ�w=���zk��-u_9����{8L��/M�L<A%ݛ/@W�'媦6/�m�/�xg�C��֣��']7�x-9�Bl?T��pY��u�PɵJH���ȉ�]Y����"L���t�aD]#�5���X�EmN��7t�x0���$M��}�����V�� ���$��"->�ܷ�S!���4<�6Y�צ�6��� A�w�vຏ6� & ��3�(�b���X'>�$)pŔIec�g�������
��)eT��Dt�LM^��ԝ�t��j�&C�f-����$#��mEi0��1�x���R�H��_��A�Y�~'���k��(sm�'�f	�) >���M�;:���� ,�l�m��|�<��ĨO�L�ipGB��sѰC�m %�/�����b������Vd�
�ܱ�z�@����x� C�c]=�s�%��
�=�%�{�c�?C��ڋ!���H�ٿ}�\4x���G�b䇇��U�M��4#�5W�ï��N�Sb�6�Vu��c��ʢ�'�aV�V���������c ����T�R2�h�a\DA��|r� ]u���ͳ��_R4�:�@�i,���Sf}��|^|��wF��"���Q�Q�.��L�8�U�1+(�(P���E��p*E�N�<�� �xw #���P�&_�����y�ύB,/
�`ߴq��� f ���Ύ���*�"�)��YW�u1E|�q�3�����#*�Z�
\L�����L�\�W�O(Ð�1V"!+,�91��c�üo��C�g��j�s�?�>N�5��
P���C��B ���(���g`Q�Q[�{����f��Ɛ�lox:��N��L,���UG�`EVW8;簅��Ϭ�!�G��ʙ�U�ⶰ2O\K-a���q�h��br�l��rVIZt��U5����-��S�+�~yۆ��v�8'Z���8|�����S)Z�G����B��oۻ����A?^擬��l��	��ע9��W��X�=˸��V5ף@��.�f�e������ʳՃG�M�Tb�'2��߽̹�D���tN�'Wcه�ރ�@󤲷�+��l���|��kO�� -kku���G�(�m>4��t�.j7N%�ƅ¶��M� U�\�;�η��M�h3V��}��a����2�����)�:�Y���ZY��c�R1�}�N*n�+׽�Ez�*��s����R��m%�D���n�������=܊��M��
E���P�PS�V��\�q#����[C΋�<"�f0=,��e_gWf' �#�l��ުT��wՕ��H�f�	�h���w�X��}�R|��C�- �En�=���L�~��V�eS��pU9o�4��c�W�>bm;�2���vX�%fg����4�+�F�>�.�Ǔ�/3��{V�`|h؜sD�a��c�Y�X�>�z,|�,�T�D�1K�Ʊ��a�g`����Hɔ�&(��<����#x/f��Y&�"Ҷ)�\E	}lh�ף�" !cI�B	��6e�
���Hd���Uf�>�D���y
�PEr�W^�sb�s��{B��N���!��;��������t
Z��Ƶ�:!Ă-�������Ƽb�!��` Fcl��Ok�f���O�^h�H'�n����!�xm�aU��a_��LǬ[��48�K{���q���<��4Ω~��5�L���5�uWxco��hש�94�/B>z�)ʗͻ~1֙�7�c����U˧ۘ�ų��;��r��V/i?%�p\Đd��� aP�ߧ���gډ�AW�"�%M��E�m��`��m��1�.�G����"�w��6���ޗ�c��@��In
�y�����a�D���$$��,��\a��Q�����꯸���e�5�"�A��-%�r�g��񄹘ٚ�9�"s�6��2����A�G#��گtc&a�#��>C�� ӂU{ZK�O�Ld�']��	�;���5��Ƈ��%����Ĺ��gs*.Y�����beЌ�F��3S!���1�=��WS�ؑG�-��d2q:��YM��?��� ��G�X��uκPyA'���B���� �	����M��+��yѲ�A���H�ێ�t�BWXO�.k���k�����;��}����T��0u�Stt�:����Q���H�؈��Ģj�I$	f �@}�+&g�T�Z�xQ��� �0�/�#1����?�3un	"����$iq�6b_Ev����Y	����bcw%d�J=����Lr����Z����� ~2�ǉW�Q�f���-��Ӧq��v���� ���9G/���uk.�Q2^�[�jeS�)�n?=L�M#�6�\���2;����I�%�a����-'D3�����Eq��%�v%�M_h����y"�� �:��ǯ����AII��r��Ͷ:�}�%�$�^Ӄ.tUh%�s�*�Һ�l����6eqU��H�A:�c4�b�e�+r��1�[�>ž����n��/g����	�B��Z�&xq@���]e��a����'E��:8�{˔W��b�9�	�Sږ�qή�����v!��u���ܪ�����^i,�g����w�0�%��`.!�K ߻�N��.�G���k��9�aW_	O�q�R5;q6��"yƨt�`���*`��d�m�֦���,��RU|�f]<�7U�Ss��d��U��<,!��Kc��d��h�S�P�0w#~�U�EÀ�) ��+"�T��ɰr���!���V�yQ�͟*��]�v�/1#�T~�����VN��&�-�/�����:��V��(Zw��rZ�e�eHC�}GV��K�ЈP~m����S=��Y{d�f�ͮ�7r7|Z�T��	TE��Cp��7�n�9�z�P�KNY�ߵn^�'1��LM=���Ȋ,�N�~8k�sH���ZH���IW�-�A2�R5̖��;��� ?6�b��."��l.�@)�{=�h��q�V�ߤ{��>Y�����ac�jP3�9Y(T�K#����ް7�&�q1��z�S[���}��%wF���*��jɭ��7%�9�A�%�1Q{����v�[��ҲD��@L�A|�_����j���k����Z��u��2������6�4J�D[�-����<@�v�����S�6�R�"�kV�3�% )�TH1���ӄ��(�O#�'Ǉ����d�ҕŐ���_���F�%Ԧ��rP���<~[Zu�	�%�I��P(�Eh7Mr8'џM����}�~Q{�d"H���G�z)_�0S����𩳯�ĵ��M�0�bC0��#cP/�~��w���zA<'�!j��l� 䢂���#nX4�¼�6 _��Ȃ����F���$��_k�H_kJ��Қ���@]�������%�$� Ao����(�~b�x��@@�C����Pʏ�^��7T2��h�k
����+�{���<pq ��a [Lx��o� �E�:rpf���m�j>��4U�	U��E�zi9#Pm��Ȅ�I�\�Sj4��J:�@N�L| �j�E��U����b-/&�@N�Y���`��v�/c�J��/�B!V�?i��!n���(���H��c�8J��Ht*���,�.B-\*o�zH��t��o�gq�S�2_�J��*�*�>�&UQ�g�7g�>�]��J���ddbQZ�B�N`�?E_aS!�Vٞ��!�vÈ�aw?�VZ,kk�;y���M�A�u<k��Z���)���+?�\mb�8>���[�+H l��{8��i�|kz)���,����+�]
*gg��do���O�*�O�+���'�&��t�5>�5U�9x��6)���.�,�|z�L����X�D�%���ya4) |5�7)�	�R������ٹ�$���u~w��b'#=�5و�S
7��#j��?��gx:ᎊ|�M��b�4g�ݸ�5�n����z	���zd�8����c�S�>�Z�E1%��v��LY��S+i����S=В��W<Ps/td�����M9�Ցы�?�4/c�m�G�����v{�.(����)C7�q�uo����HH��'�
1[t��;�`��Q��hvX��D0�N0�~xa��@Ψ��F��G�$#�tǨ8Hk���L[�;��X�����*�a�8r���v���M�<���wK�� ����uT�2lD��=%l������ ��Bɮ�c9���ouS��!μ}pxA���1�f�B�M޾!Iz݁�=�MQ�V8�z���q�*�~��cр	W�L���9�3;���p~�'���,�L�2��XJ?�y�+F�)��tO��Y��#�x�����+.��"�U�K0�}�^�݇� ��Z~� ]�y�?������Q҄�-p:qA�>�Hy�ڢ�H��z=��y]��A��Z_!�2&4�(��э�?`$t��X�&��5�2{�����Rkt��D��6ލt���1R�8$>���_0{�:��ѻcf ��ZI�Y������B��'j���0^�`�е��](;^�ؐk�
j�����a��BS!������̰	�o)�����Ի�׌�z^�~�gbٯno���f�ua()P�_'5���� ��/\�%R�P{�/Q^����6���p�g~��ZLA�W&ܺQ�P*���m��שV���ʉ��	��4r1��%�W5��ב���!�H�8��hݺ´�|a�/)Dqi���Uk|��3ް��V(��Fq����	�p�4���^�)\ G���G�3z��U8�|�9��󁔎�Z��s�2|VʽSj�/�c݂�ܩ7n�q�HP%�6ￔ���8��n	ɒ� p\��xQ4��WԴ�f�	d}c)P'�����"�/Cphf�z���
� zƆ�E��A�ȕ?zhz��3m��M��z\f����o ��G�![,*{���4n�X�s 7gB����ӹ��z����K<B�}آ
���	b�*�x���%�s��H~Nq��8����R�c�W�'W�I18��|5���rw�kK�ݤ�2��&"���U���-).�>z��ZH�"�B��|�e��w#���P�JHš�꼓b(q�f���I�-v}���(6( �?��������
%��~�B`1�+�v�E2#�A�ڹ��on�W������*֧����@��ǩs5ū�y��ahOeiu��<�<~7|�pJ?P�!����㌅�p��7�=�5 �����
���2��ޥ�P��y�Z>����Q o�~�:��A�=w]YpQ}]Dlȸ��Al���,J�'��;9�Y8�C�v�=%B�T���&�<�5�W׮�	����$F-�<Ҁ��,�ݖ�B�:��6�3菏p�DO����?�kY˕��Z�.��b\�Rֹ��Vy�Qlˡ6[�P��P��z�ژf��~p�Z����e�s��T��#��&��z~�KR�wC}�~���|~�wC+�q\R�+EoD{���Ր�u=�����L秝�ʫo��{1����s��â�b���
yܠ�g�$#��G��~Φ��L�>Ȟ���%�C���9x�j-���iR#m-���z3���7�@ݟ�";�P���Lϳ��m.�Fm�@'5�\ZإZ��y�J�i0�C�r)ڹWت�$������c�R�#x���~���[�h��iy������b�gX��#�MÕ{taX��_7HW*K��۫�es�~�D�GuV0���˶.�:� !�S���nD��}W{��gʁ�H,�}'Np��LѠ�@��k��b�9��;��a�����Q����Q��(j_�cm�yjܥv�j�qI���x?Ҫ����Z@?�P�H���Q)�֪p2�.�FC�����y�}�=��J�j��O`��=:��'J�Ŀ�5λ�o@C&4�t����O���;��G�UU9����b({`�/B��y���xd��5J�I�g
dG��3~4�\�;�"��./9����΄��%k��"dV����f��#L����n%��p`���g%�����U��Ek�FDŠ"�-G2���������<J<��Y���I�����w[���S6��x]��q��1�5�:�m� ��#㐯�8�v��.w�m�3/�� M�������Ȓ���:��b�f-Vy��`Y�_�o���� �#��Vޗ�Ha�	�����5��tuN �>8G)�}ֳI�q�������Q��G�$��Kr���G�w~B��E:�Ք��w�/�MXV>����� ���o����g
����Rv:�0����� q��`�v���&�aEW-i���Zw�������4�1D�`!���1���o�׷�����7�����D8��׎;e4��艖��"=eFM�G��/�sS0�y;OC��J;�-�A�l�>���)vG/�ؿ8L�UĪg�"��Z��L�~Y]���)�����ӆ��t)c�u(؂�2Ή1:�AQ0�,i�-ƌ�厽�xM��t�M�jУ�Ʌt:.�5�V���0#?e0�3)��R����!]Q��n� J�u��^N܇u���Vo�#3�l���V��nz��m=�Iۏ���1-���|DR����L�	�2�Sx����%�Jb��R���H����Wk�0o#��gB<���� 1Qe8��|�ڃ*����ܚ$2���v9&���.]k������^�V�F�0�/�=b�.#�2�İ��!�4/Ǫ)�F�{���m6r��9E�GдM3]�"z~�}���	:�aQ!�I��`�fT3		T���;vQ����F�`$����݆?�;�x�r��P\fBj��>u�a�|[�j���I�h�k^T���e�W�m���������NQ
J��"��Y ����2y:)�U�ދ����J[�����W�����������~��l|țwe������Ր�Ќ�aޘ��c)s���Fv��6����F>����P��0���sq���#�e�����9E�L�S�F�r+�I���Ľ�E���J3N|�(��ϩJ�IM�l�܆x�i3�g�ͯ��R���� !��[�9hk��x��!���6�}X)�C�;�K�aP�co���I�+?<K`^��E�@�F�:2'� ��4��k�CJ���xa'_%$��rg]��n�/=�+���桚��?��"��ƙ�D���ك�U��3��.��|��bMrG'	D\j����x��f�I3�g�@��3�յWE~_[	\7�~w�S��uX������K�2�f�{�E)K����D��;�<V��:;�>�A����!G9�x��nuz���`�z|�$<�#r�uyE��l�qn�Y��ro�i� P�yM��9��������1��<;m� ��|����h����!����J��jʒ?�Vջ1QbQmtR3|��[��7I29��h0�23Z�1O���F����[���O-D@Kh��!��Dl
���Rq�����"�h��
�u��굃��,�����r��nX8����rf� ���RC	V��/8v��F�o����~>�!�_��+��ia��a%x64��f�I7�ZD8"3���O=u�����_�������)&N 	��5��{rBF2�M�U�i*�Yn�ܕ�"�Lwɩw�lᜅ�s���8��4H�&�؅��f�s�������q����Bٰ ���� �^V��|��6
jS�b�B�7]��^��3�O�&
p�4ؒ\eW�q�,�v�*�@mr�e��^�	��S���9���Dbe�}Ji(�/H�λ���t���tG�7���u{��"�b�oOh�ئ�a1ꚽ��s���>ȥ�њ�m�@χ�q^%=��q�L2��:�1hl�z�l��B�P�Xă%m�cD�����H������/��7X\U*�+�|�Yʍoņ�T	C�|y�#)"�V�<|��N�tiɝQ�~S^�>��Mf���Ɇ�S�f�	��(>CG=���K�F��������0�Q�
V{�=�]���8:�v�2	�7ُ%��2�DGo�C3n�Z����#��V��qPے��}�Bn� �l�&��͂д(�#���%@U�:r'��J�bk��Pz�I���K-�Ӹ�CI�9e�����vE�R���xO%���V���G�P_�.>(��[��z��\��\�����A�z��.��2�Ջ�8��X����K�c7uմ	��J>��e1	����ʙ'ǫ!L�b�*s�x���'�(�9�eN�GJ�R�:wߪBŗ���U_���q�ͣ�O'���z�FOy�����j��S^�p�ɸ�/xUA���n+)��e���,J,�J�9BwI�L�Q�]�8ƛ�:� ��8@���j^@�Z;\�?���9Of(%1�"O�����uJ����͚�*��%�N�l�̂�Sl��e��xr�_�FPe�NH�����|��Mk��4�`E�W0�c[%�gv�SN�����dBo���T�NҚ�p��� �\Hs���r���=V=pń �P#��[��1b��8�a��ۄ�:5����dе�B
�����̗`)AH:N�9`F&�kH$2�K[w;�i��$}���)"�J S�5`<�_	����Q��<W����/��&Q����=鼢�Z`̿3��(��L�	�'��Q	��췊�u�� TY����0)��n+���"�ʧuy�0�4�|�����⯋mb8�٪Ց���S,u�3Kާ.��2OK�3V��p�D'cT֖M���~�&rQ�0���O�u���dIiNF�X����j�+"d��i%�A��h��0��`t���.�g�l�SrF��/�iC:�  ���*�#\OE�XW%��Xls�ض�F@�o���=gJ?@��eK�ĥ�kǜkI0D�k����L���>�W��v��]၆����15nj���q�������d�!��	�v/��aYg�|R[�r��{���̨eK�g����#�R�K���g`�{�	��<���bJN(�nt�u֭�SX��1���w*?z��z��*��-g���j�x(p�	����z/S��V�Y7�<Q�|�SUd��~��=C;m0��Fr�*�7��t�MKY�l\�BSۧ�t㔠o��EVLBL{���������0P��[�E� ]n]˓h�#��c��	L�R�2
-w�Y�&��w���3_<�8H`�S��#`��"��jcoQ�xn��WNK���[�BtR�΍�Nw3����8��yg�&�2qYL=/�OH��1fZB&��Tl�laB���?1��Ձ,�E_dy,���&�ʵ�Š��&(s�J������c����(,��Q��<��K���	�Ca=\�OY��K~��b �/�9ZYSDT��#mhC.[j8���q��.1v���ŎOB�s���o�>�����Ŧ�BYRˌouU|;[c�Hk�8eR�ʏs;�K�������b���~�\����{��"�7�6���*�	U�O6g�k6�.Z��!�R�)�hft�Z�v���;�P�c����^��x��  ~"N�T�`Q��m��eP�Ș��Rg]F���䃚���JM�!*��U52ȅӾ�L�Y?��&K[�\�/�d|��d�t1�h#F����� �-n3�sti�a��/W��ܻ����6!�K��#r(Id!�6Lm$��ӱ�1���|�{3<8�����x�ksͱ�Lm�[;�"�c:t41
�)a�n"�fJ?���p�B�\h ��I�R5�Ck��K����}�"r�"W\��=�xv�"��5�^Aƾ��ѕ��#A�dW3N@Ek��Y�^�s�c���,����-�/ SQ��sz�6|��6�L	%O�?{s�a
Y(D��G�
[وI������L[.����r��U|w�.9������GQ��
����'���4�+OO���h\��E�׏����:b2�U��k6f�h@��"s�������H��uK�vCF���CU�9��c+~e �zP���Ebq!I5�\�d���:p�-
�k�-�����9�}�U�k����*y�w� g���6i�j/�U<�SQR�5E�"/F�n��^+�<���Y������Z��͟�tn;p�u�S�J�M�ן��e�+��ܽI<B[��濺(�Tw�`�і~���3f3����]'6	���Ϡ����J�:���f;2�+�f����68�ct�P�7��Lf�rG�u<���suI���73C7N��K����ce�܄����Mc�bG�C^�

�9c�1��"-��Ŵ&�e���j�D���%?�b��L"1Ҍ�LR�"qm�*���n��H�¿��LJ�Je,yl�U���ܩS�%����tG�ܮ��'���b�`<�L�X;�J-�i;*�glq���}$�k�'iX����~`�$~R|��m�<=��>�)I �f�[�f�_'��a����OcVg�Z�`9�N9s�|�@�ϥ�z���#ە�]�{t������������>��V�y���RU �	�~�l P��T1�@L@�s��^6�2��}�D�Pu�W6�R?�����N�2 cJ���M��FL�"�׀��;�����h,��'/�n�$��w���n^ܧ���Mg@�M��Ԗ~�E˟�'�u�}A�����&�")rn6�^�����������8�*�����>�<���?l�$�:n��XՁ�`�K�vD��Շn}>u}<�����Z9K�F�:3h�Smk��z�"��]�ξ��z7�p�hM��+m��,%����n�C�C`�·�a��_B���x0w`�Qoj��ܩ��c9?N_bɵ��Z��:��( �S|auDƿ
�<���j�Ǔ#�h�M]q�8R�G�&A��Ȭ�٤�w��5���PX�v�BͿ�������+�#7E���N�����
���L�@��!z8�l�z�I�A3�6�s_�,%ի�G:�8 ڰ�C��y���@8u��`�8e.J���I��z��#�Ͼ�0�w��_��h:�ND��f�����%���E��2Hh��I����l��r_Pra=)*>��/�˵���wX�Z��|=_6�v��?������"=��e�s5��sʙA�1LBA��ɿ���X[PM'�XMuNB�q6�"����j�ݤC�Жl|y�>�g��|{��r�Y5�Ĩ�(2�zX�Q��1�]l�Rˎ�U��ZPpy�z
 �T��y}dI���E���^6��Ǿ5,������p��]%P���?�;��.p�]%�`T���a�D�3��%��ї�o�w3�����lI�tuԛ��v��۽<��X!^yH,s���A:E&<?��r��M��۰.(�?(4͉v����_�a��Z�	�й����n�౤l$����At�$���U ��h�^����})����9iC?���o�~~x�UR�6d�E�Q>��+���Z�޼2k�,� �������m]��^<�#��OY��|�r�,�x����ATMx� ��^w ��I�ּ�}��)=�[@��cJR���<@��#�X��΅�4�)o�C��;�2�kO[�c����p||���~����+Sh\pC`�#�>�,�8X��|��%�FN�����)Co�I'���؂�o��RGX��Mb�R|Zg�K��[��@�V�gl$�C��(����"��Yg��+�����nBt� "q|A���:i�8��M�О�t��J"Ҁ<�FWC�:���q�5	�\�w�(���p>���T�g�*p��=�6�>��D��w$��L��C��t�y*��0�51�9�Rli'Ϭ���R�'!aqԒRݙ�)/��Nf_p�� �D��K���<�T5��du�-�Z%�d�]��&���pA��(�g5 �qzD�d��r�¯>=�������V�皿2jh�ʁ�%E�{u���L��z��8zN�����t�mdra��,J�y�������{5�ݥ��5��X����!:I|w�7kL�?6�"�}���?&�����>&�7��A�i�g���*V� �A1��A${v6W�F�[콱~���Ć��+)���r��!7vmI&O�v̎��0�u=�m�@#G֧�g¹�,���N�p7�(
z����������&��[{ZL�s���C�I���G�@/�E���N9�5eɶV��3)<é�/���Yc�]� BO3�zd/dp{P,գ�EX���x�m�7o���zr��c�6�u�D���YUC���<q{�>	qd�90�<3�ul^L�?�Q� ���ѝ�vx�� �ix�,�n�p��Tct��K�_�R �v��6.�R7B��6�d��P���6��/�r Zު�̴����_4-�K���L*}"3������H|_&��(�����-L�@B�D;)H����cG���^*����^��>�5���Q��"�l#�A�����U#v��6��'V���_'+B Ǆ�Q�΢
w���Ʒ�o��"v.|��Վ��"k=��籘Y��@��d���N��ML��-J�O
�,��0*��JĞn�!����"�������"�_��v�q.y��7A^pB=\[{��A�ۡر�Z@[��8��ډ	"�D��a���Pgvߝ��+�y{	�i���JK��]q8�W�&<��w��~5�Pb���Z<�g)A�g2���(�����86��u��:3{=�_4�H&���k�ħW:f7��+ZU�u���>��m���t>-�9��k-t��z!���e���\b��Rķwk��z�-��$�oVi�����[>�@LP��Xs\�@ި�@�-�Y��j�-���&m�Fe�K��� J���ZN��k�I&�#Jkg6��
���_��j�%"�^+	��(-���љϐT�f��zR��z��k�3�xԞNǧ�Ed�μ�� i.M�fj1\ڨǽHC�׮��	K!%��F��Q�J%�z�.���T���̿��A(P�����%�*x�u 6�OV�b��q���@okN�<{�k���\�������O�uH��y�0�Tf�r����n,��I��0�q�j����0(��/�>,�	�8:���,�ӣ0��9*��L�Sj�b�;��Bfg���AYy+�&I��J��\�D�(�G��u:����aY�0u�r�f�
C!��3tv�����s�l�-ڑ��%Os/(�#7G�G��1]Rc�f���?`�����3y���F�e����yh�	��: ��Fܺd�I^Gq*�
�R��X���u���0'C��ڪv��~��@�?7qK�>쬔�vш������]u�-�7̦��Dw����x�v?�T�@/9�&ݴ�1�;��dV�MP�.�q��Zj�A -�Z�L�f`Yw��$P]��j�"�5��P`�OP�+A�/�d�#�f�?�x�Y��XC����4�UN��w,�J�	6��{,R^��d!�o�����}I�6������@l�4pްޖ=	g��;��dy�?��a8l��!�B]�O<�N,�FV?kK�&D��;�����vȡ��������m3#�P�ձo1�����Μ��L��Է�{g��~�N'�w	��E�?2��		��#����5t���xr��8�
z �PQ)cT�v��Jѥ���9�\��.�`�w�*���<(O&���S�"/y���m�w���땔�m��� �fP!�t��~�ox��l���ˢ�����֡4�-/�Ϟ�
~L�����K��G����7��@�x ���z�Nc�~(�Xo���$����fReS���E�
Ps�斐�c�ʹ��i�NG���}�����:�-9�w��6���m֮�8�}0�
��/5��X����;Fd	�k(9?��B�����o�?&�\g��I�w�ZC-���;�|�����:3��R�n��x�V45F´\�b\�jUD��\�W�;�}_5ԭ��`I=׺���8�$��-!*c����r4��¯u�5>ֵ1
u�e�廌��%*qoD5�.�\[Rx��D����(E'�c��L�aq]�P�YV���u��0�u@��4���`h�G�~�c����v_N葷-���f�=T�P�9Qd�P�����uOi����<V>�R���Riꩿf��0S�
���~�ץ�k��.R�����H#�j�	C^�Sp8�~3�N�O}1HRI�%v�
��Y�?�9Ǉ����}�c��/��$��'[��6������Pr��
V�{���%���M�~�t���~�y�Wsf9%QY8F�mк1s����(����ht��<�7�>ݠ� �X���H�̙�/��@W�ʺA�5�P��p��]�Vb����<�1����+�ŷ�r;s9�Zz��̽��u�W��u��Z�yU����� �g
�o�l})�1�l��{���x>���D��M��8�������|�
6�_��s�O��vv}j�E �ò=z��ۃ/>k�-��f��T=���#��Q'5=椴��tI5�=q&�Ǣ5��ݔW�J/��o+�e���(���p'����+=3bO�k,�W��!�~e0�#?Q��N�ZZ��qJׯ��A��-��J�d׽_lƉw��՗=ev�PB'�92�>�6Q4��e�l ����͉I�R1��m�U��{5@��	R��t�Mp@wҎ}<��E!@�Uz�QL=�#�$�Rċ6�{����u�i1��d�F�.��v|���'�9$���ǹ^܎�����gr1���_�H8׌�Όf)��Г>��?�Gs�F�ȳ�N��{f���E�p�qZ~8���X��*�ؕ�Q�)ér��f�'�p�U�����Mc�ˈLzq���n�(I�u� �K���Fv<�.�e�����ӈ<ױ�ަҢ�yc�$��h�-	�f9�fz��� �E��>T����slL��h�Ӝ�J(t��ŝ
CӺ��/����}ƶc�B�+����^��lw���@����=���&����Y8�R���8��'������z�N���}�����E_�;� Ȗh��C!�r�Wl9ݨoH
�Գ��l�x���`w�G�� �x(sUj��^�9����9�^ 9��iz!4Ʊ٢��Jʟv���esE���i�.�-U�F���Q+��ښt �y5�l�\�ZAAW�7;6�zZWA�f���Ŝ����32Z	�l��� ����*�n�T�(���
jy���s q�l[ȭ,P��o5�*�@z����X���� �]���%�w_=Q����?��]�ā�a��ݰ�׌MBd��_�B5�]@륇���yl��#�� yO�6�{��y���	kc���s�1��Q܋�����z�$!�_fW�!*cA��T</��)f���$	���1�𞯳a�0��}�vJ޻c�d~2��&�Qݰ���O5�.x��٦���p(`rXm&��Rr_���������"!}�z��&$�w&�x�_�;�3���^�X��@؅�s]�0 �����סJbB8�-���w�I���Ě��i%u}��!A�&��0i���e`�lm�D)$|�0�l�/k�������/I���X G��Q�ח���1�a(�X:ޓz��hGk;,P���f1y�{ǿ`叆T ���9���\�p���d0DeU@($�<�=�
���Nf����/\��6]��XM�U��~�����\�A:���B�I��+,94uI>u�x����O׾l�$:�S	���kM�t�3̿S���p���j��6E���cF+����]�K/�Z�����i/k�� BS!��gQ�O9�*��k��SՃ�� t�LǙҕU��
��<@(��.���6N�J"�#�wr��嚖*��ṜRGѴ~��/�j�[k ������]�����]9�5�=\v�����:���2�bZ�u�¥�h��/@jn��&���g�rϢ�ϊG#s`-a-���UC	�"�70�bI��S�����N�c	EFy�Ϳ@ͨi�H1�u6BDI���Z�V���8[��办e4��:�H��l��	%�C`P޺�K�ش6�]�?�Ȼ��������y��Z�jyY;��޳��2n��RB*
T+0^ND1Z�
�G�$�Of2@S&SH��wF8�ד }G��"��EY��|i*m��1����)���2a�/d��E4���y�q5S�,Y/�j=[%�<�qB�է������c�\�ąk���x�N�M%����b�+���1�u�
���v��ݭ����DZ(x�S��J!T�v�X�W�>g�����f�Fy0�\�L���gg�韍�սbvYFߴwV�iӏ�Z>te^���`����m���W��`R�;�l��͂�v�uk芾��v_�(~��h�������{󾅅�%�i�|Z}R�Vko����% GB"ʘ��v�EG��D��+
N�T,Ŝ֫��l����=�U�������~��{8�8�W��.�<L���A��<짢���]:��ƫ�?������4���	Ã��(��k�x �.�E�W�\r�)�5����.�٠	3���p��}!��ߦ
��&ʓʏ�g��K�bOD�צU��W��Q��p���\�,bP��_���\�#�9��"�
Dź�Kb��EY���@��ުs�O�A���x.�4u]_��Q@�5��x�Qc��/$�1�Z���K0t0�J��gaf��Β���4�n��1=�	��7Doy]Y(��P��ǚ������>�j��,�|n�����[<�r����u9<�P���23�ok���q�#��/�x�� ��� �
H��JIʧ� ����'�FIU,q��F�?��ˠ�>Tt�v\����It�_.+��P�n��*���U�t�����O,�)��7x�Gi�W�<A����)�� ��4r�mAba���-̖	�LT�LAw��$�o����A"���'�g&<�\������C:��:_$G���4ܮ���A)aB��\*���+���^�*�w+�pQ�X�}B�@��w��~�Ɋd{��H�.Z��\�嫰�W[W�$88g�/�/^�\ 	;y�a�mg�ԍ#�r�2���L�"��o��s����u8n��/E��錰d=HI��T�J�E��P�v�@*�a�ӳ��	^��7��3�9n�c��8{�SP�Z��S��H��'�à|� k<uN�_���.�9_,�K,��%sA��;	GG�o(��w���e�6FvjςL�Vi`��Rof����K�
j~����(������!%�"^i�����C�kI{H<t�:�1�5�Y���������*2���.��D�Mx�;&b�Q4�h�Q[�IW����(UӦ�lq�l4��v�^6&R�,W��Dh�������Ɖ$��W1�6�#��-�j�hB���J�.��+�9�7�V^�����C�'N���9!=@�g:'���0kq�#�������]J^@�<�g��h��Ӡ�t��GŮ&;�"!�%$u�t���3�FN�����0~i�v��aۈ	
<2�h��ω�\0����wA�]�Ĭ�^]�B]��H���R͵�r���x�N��Y���S�'\W4Z��v���n��*V��p��h2X�K�a�6��*�_�A�k�g��տ9rs䳸�cRu���� �28���K޶��զ�kb��D�@�(�c
^�82�s��Y��E��Ǒ���smA���P�\;�Hv��>��*����s���j���JJ�f�c�R��^�/���L�ǯ��2�b�����Ƭ"��M|�<�E��Fd
�=Z��~s��C+��i@�Xv���	?le'�;�b*`�qw�\ͮ]�P�Ui� uPiѧ�N��ʟV�&	��'�'�w��G��n|$�$�T�d����^�/*�Z^yb_�9�3�a=�$,J�7��Y�_���CqI<wzE��� -̈́U����vb���'0�4���%��W�ՙ̡�����s����1��ic{7�Mږ�~6�w��@���[�֑x����K	4��a��0�϶���}9<�m�S`�@��o�|f�S�Ǎ�y:�U�+u�Ke��ˆ�s�9951<��3�yl�(�8sƋ��\v�����������vB.��B
Ձ��ٓ�;/RK�7�ī�|m���aǟ�b��d��|�P!F`5��
�6j̛0�`
�!H�����t�k��`���)�Ad�z�A���!}�/)4��ùo��u�����?;[���*�7�M�b�HjW8V[�f:�
�yN��(�{z��k!�¤�IZ���0g�b�ޅ��$�l���!6�H׍�J�V���lq\Ύ�iv>]�dk�0�A��h	��&��)��l�$
Qg�gk!�\^�!�!���32�/f�8>Ę�yqhw�;�
a��sA�����[.&*:�����8W)���3�`���p��F�͌�u�|W�l�}���9�o`j�+��cp0:/e�Z�+L S;��� ����@��p.:nd��*n Y�G��d��x�:�R�}j�.��fK��>|���-�G+E�#�y?�p�E�؛ M:"ε�_��Ed�<���x�ڌ�O?
��[����^�;;0�o���+_Zc������u�-�*s;@��hWK;���ψ�Z{�}ͮc���P�(�~��j�U�h'�uooV�'%��
�l�]�'~A�j�gYLM/9"5KH��}�1���tZ��AC�f�G������.��&��C>.P;jޭPRlV�\�g�4�����p��>�%���������n��`��!#��&	:c�D�پ8K'�fOD/��ӱӞD�"��Y;�i���ܳ�D��x�-:2>�=�	qy��W�tJ�V�PbM�Y��>�vI}��	9h��'��l
���R1$�q��m%�m�Z��J(n��CeJH�ga�JzΊ�\c�Rf�9�lz��	Hr�Y�En�
 &�0"}8�e�u�:�|����ҝpWp(3q�%/�ݦSI(���Ds%�Jݓ2���/q�2l����_k�E�!��S�O~Gy�~�)��W4ޯ۳C)w �ׅ�](�K�&m�iޞ�J�hv�&i%�_֊*�CPd۰�Y��X�<�hү��@�XͺV����Tkd\�22u��f�è��t��4֘���6�\�Վ������nO��e��ܽz��bl�~�� �I�;9>��[�=���}>�7;�<��(si��/'�Ĭ��P(+!�b�Z	!)��:�2�}N�c�l.x8��YS��v�-0�|�/S�=��=�QiDdR����sn_�OI�3�\�r���_���}a�w8����/�4Q%��&�>.y�5;��A&������6��H�ύ4ߵ���	�eIo�R�#|*�L1������'"M�N���ֆ�A�Lm \AG�i6m"n~I�ZxmV�M�PT��7��v��6�̥��ɷ5�4�Ӓ'�U5��(����F�r��P�U�r��?Q�?�����L�(r8ĥ�[�j]p��w�Z)���=I�aA�{լ�|mk�V!L�A��9�{c�n���ر �n&�[�49���r|�d�_ÖӪ�sY�]�q p��2��!�歑��	ژ���uL�mWƋ?]�A�cw.�7Mٗ_[γS�1�8e!�if(��͓�������6!���Ţ^5*Zo?�ǌfGNd�	r�^ؒ�p�`�g{鹙�/��hhjk�Eb�������.��@���3�R�ͤ�Dk���Ӑ�E�B��ڣ4œ0u@�I,�������%(6~m��>V�8^0�jõ=��z�g�K
S�5�{�p��b
l/�8px�H�,�5x�$h�ħ���R��7:�a�����7���7���k�Na{���%Aãbf�s^b P�	��Q��g�s]�@�W�v��p8}�F;w�g�'n�"������B�Nx\W1���^i]t"�s�h�~X�����M���>m������b�&�q<����®�OYkO���^36=�S%G:"��C���� �x�D�z��ݿ�T�ƙ�A�r��/mɵF��ѝ�t�h���g��fA���Y>2GMaiF�!���x�~Pv�)npKÚ�[�)@Q�#���b4478x��CP�)
U ^�
d��"�-1LH#�S���(�w^��wf���D����&
20q~�؞�ޡ��#���������։X�v"�C�#����5gb��e�A9�6�������\6L�!�/���R��/a��t^�*�A����י$l�q<���'�i�rz_]���K��}I���S3+�I��-��>��M��D���0�M&s1���%�F� �M�a���ÏRO�z�<��=�R1�[Wv��=~w��{�|fz���TF�P�O�2=X����Jܨ�C(�0�ގ5���u_1�A8�!w�9O�p<�&Djic�Q�RL3��H�2,�3Gӝp;w��O�!>��šB(n�Y6oW��VC�$/z�u�Ǚ��ZjHm�$4�H��ͺy��lM|����(���t�X��|��U�qZ��#UJ'L�p�)�u��9�nv�+a��]\��!��,�r���fS�{���4�c�&���g�kZyK�qz�K�)o���/�ǒWʢ��ȏP���@�POC���:����d�H,����1��-\����EIG��{�]����L�=���[$	�6`�<���1 Q	?p#&�[?�o��گSj#2WS� m-��3d\frM��)�X�m��*��^%z��Y�Ʊ�鼺8k�m3M�Ol��}�8,V�Կ{�
�)⡾m�,W�����g������O���*@�ݳ�Zu8��W{�h�u��ܕ�t�	\ T���ߞ�&U�6��	E�0Y��4��'G	�J�D�̍�t�C������.�j�������r�i'W�_�8?���}��|8�}2L)���|�
�#����>AC���?Q���W+�l�9us��R�U�q��V_�7QWt�ax�6^�Oōc{Z��,{	������g�c��z�� Z[	�Ѵ�J7J�1�)A��͛�1�v���o
,h�@�؄y��S8�Q̣����!�u��i�G�5�G��z���������h��$�6�hT��K�X���,爾ͨwJ��")j�
�ͽ��Fq�����U�c�����dB-mZ�|u�巹8�mÂe�Y�,������b�T~lS��̿�jO�I�����]����5�X7���2љ��tҞ)3���~��CGj>k/.�u��>�����H�F����]I�=�A�K�u��e�e!KZ��<A�ʠ��68�1��W�_+�}?��"껈J�
7�ˣ��PG�)���ȣ2�!1�2$V�1,#f����]�8R�8�CҰ�/���E������k�^�-�U:��)T�{fV�pT�����^� �O0(��v^�~+��^G�M6�}#(ŔT�5?�����p�-]6t��	У�j��;�ܿ���K[{)�P��~����a$(�f��l0Y�6���j�k����g��n���m��g����������V��u9�����>4�eǬR�7B�����>{6����K���H<�^�]@I.j�[�C���s�[J�P��^�״迵H���t/IpC����+dk�O�z���ӣ��xr�6�&��p��_��Sk+$I�s�=7��^��vy�̗@��j�
��𼆽8j���7%|
!d�$JDiC4�9��K�9i�6X��0�G�Q�� Ì����Ҧ�8�� ߺ���� OR/�Vf���̟��$�I�������%�F<�����m��#l1���%�m�6�`i��7r�+����;�9�Y��ˌ�DB\��^zE8��=zH[�[�6�I ��`�a"T�&�)�w��k�-�|�. RR���nC{���(��1C��*�I��~3��������}�6A���c��d���B�6���en= �O��^����y��/%��e�_��G��$�,�JlieB�I���p�/�-�sG0���	,ڠ�3F���_{M}+!��U���%�vm��<܀Bn��Xs�	N��ܑ�q|��߯
~K�[��Jua12��������r55�*�Z�)6�/�\�1�o	���yfj@���}��b�X�W��a!w������!�vV�ރ�2��s�`ü`RC?�R>�=���9���(@n�{lR��z? /*?}6)�R0��"0���b���S����U�<�;�/���o��E�{��a�U5~;z�N��O��Ɗ��Rt�T&��Lh� �2���y{�6�j�֎�3�&39����\4��=9�Ψ�H�iyp>O���=�B��%��N���`=��}�b�:���l69��pWue��a��f4ο�'�x�k��뱟��=c_o�sa..��N�v>�(�_����8��º�}����5K��>_�����'�o�����I��fqL�q�X5�":ض)��%�5�d�|�D�tT��GA��a`��a�w.B)oC&�A�(�rs�b��T�jۙg.s6R%�9lq8؊!�w�J�4�̗�i��T���%ʹ�P)ϼ�MY�4�s���sl�`����yz��י��F��`�~�>ɛ?n��1���������άx#?#�M�n�7�c��ȋ�;v�	a�k#��*W����J��_�܄21�Ү�RR�e�� T<�[������q��L�$��Tn>�~�q���Y�6��;���
�E��Q�?6k���� ���ʋ�#����t`oAha��}9-yʨw�"�����zۃ�O���*�#�-hN�
�U	�c�Wo�bE:�r_ʿ4�UĀ	rD�2�h��?�c]l�t]l��5�V9�Ua9MPc#�l��+�7Zв3�
 1yk��H�r�����E�yp��-�(�R��>r��s,�2d����!¹�J�e��sxys6`���������Gw�a�K# ��Y���BaL[��z��}1�	�gܿ�ě��k�_���1p	}��m���]����1� �4-�_�M�ȷh�N�mx�T�Fm�p��t�J�5͜*)�~fx���m�S��N��:>�0yނQ/n�'ZQ�~���U^��h9�߿,��ܹ�g�&���cc��M�M왈<o�jы*NU�Ǳ:;�1�4`Y,n��/=%�oGp�c����<���0~�ID�D���� v�g8Eh���fO���n�l7��N<�T����a���1O��jR޵9����R[L{A{�<�b�c���Ӝ����g��������W^)���.T�k�5�l��̀8x��J�U�xH�R�����L��a�ѳC�����$���"�EG�P��zp8���!R��1�t�u�T�.}}w��Z�]N�}��t,Jܔ�sJ´��!wJP�%GB�jrݕW~�upw��O����?� @2!xd�0�L��8�3���g�<n�jn���LQ[��b�^@>N����7H�~�WR�����Qӳ�l�`ژ~c�:,�S@m�~gҗ,�F�n��_��9���H���"2-�񄾱�hq���6-Ɏ�۬�����_[3xj�^�Q�"|��<�p,>�4a-%LL����W��]��uG8�(�>��`$��#�qK׶%ş	O������:刍K�WB����'�����E��nF�r=������
q/H�,!�%D,�l�k��:I�$(�O�J�y�y��/��s�뫞w�G_���D�YP1g����HH�+4d��S���uػlm�� �d���Fyl��W�S62)�n*�.�J`�"3�"����������;���T��.�52<��Mx�P0ؚ ��E-�$brW*�:�20@��h���jzξ �R���r���O��i����������I����O��G7irt�i�=N��m3^�FE�2�+)un�K�H������?wI�<Uhx�k���<�'81L�L����Ї�J�y'�v�U�^�����qmlz��Ŵ���7)�>�ʄ�kI���,3���*��$L)�	���`���%H[����γ�_���nԛޯf����u�2��i'+���6u����C���3�E����h�v�A��L���$��EU#"2`�B�2d��P�_P��� �F�A^���3��`�=fV_⽘�1�k�X�N���r\�%&�ݟ������q�ݯ��n 4�b�*Ӌ�\r.`��W�,;�E��k���$H�����#�YV�W�w^�%5L�g�f�k$5]���{sr+�4����x\/N�0�@�O�jsel��=� #��^���+�?!>�Խ��v�gSӇ	E�]Q3L.��w�yZ��R��X���f|�hP�/��ǐ�P>��������zXd�>��6�t_a5�ly0�ޥ_�x������	����~��m�)��hP�+&�׃�=�8��a1M[/ �$� h�l�5�D]e�n������Pr�.�[�rmp�Gc��s��1��6w-{�U�X�3f~�O�W;�s�	�����+�*=��U�����A�h������hY�^خ�)��L�� i�)�~dt��8�]�5ಬ.3�1�|!�G���w���^E�RGxD~�~��G�a(�JS�K{�+���	X1�zu.��H8ũ�{��3i�w2GA���hXOv�����]��T��Eqhl�����}n �ه�S����|c�2�=B]�K������+�m"��'��Aq���b�[��A��]2�!v��k�U�8s�+@�uN��9�p�R�4#��ʡ����ik���h�(*x�Â�V���}m�L`���~B�M�9�Mm�We���Ag��k�@1CL����u�b$��s;����uB�$ ��/�碋�jO~[�j`�F�.�b�ޮ���J�?��(������f&-;�i3������Y㧈�����,ЀVXIK��Θ�v}sHZ��+p�,,���K]�"�ot�*�X���ɟ�J	��eS;U;W���yj��E�0���OԞ�!��+��;�"4ڬ�� :{8�[Y(C�8�|�g@G}KE�T����:&W^(�-N��d_�m:�IHT4GT��sm�D�W=h&F��@eaؔ�����&�D�j��t!��cc���Mg ���	"�]��	�?�h���'۔����R�X��>����s���h��սoha�h)d����"F����p{2�r���D���:�H��3@%�/ز���*s0���s^�A�Ǥ/�2�g1ͼ6�s����>hB: ��GQ����o�Ⱥ��^��,'#��������"�H��Sl��~<vdv?h0�R?��Sm�c���%!�JR3��D��r�ߌ�����q *fg�җ2i;�:+l�$���fi�t5���� E�=��mm�t����+%�K���Z,!��M]��G��F>��O����vG��	��z�-��+:	'� ��Bm�:b�Vg���W����jL��x������-*R-����U\b��N�D��{�F�1��|�YBԤ23ZO���]��F����^��|���=Y���#����NIMg�l�ǪJ�$��G�iwy����?4Y+M����լ�҉�2�	Pwʶ[�����|��~�1._��5}sY����hJ�`�n_A�;)U� 7� �QGM0��xe���i2% �	\���[����^��X#�㬷`>�Ъ�U����m�4�#^�o�Jp�S�L���>k���iB�����D^�_�9K��;X�@ެ`�,�Ol��-2D���U�Բ(Y��c���d�R�XYcU�G-be��C�cը-|5��l�A,��*o�܂J;8�#���+*�&ץ)�����a�A!�CU��"c�~
�n���u㼃3�D�:�m�Ĝ��U �Ā/�9�Ñ'�aJ�ak�SiL�er�,�U "������;u�'�&T.�H��2�-]��!#���8��K.B[��8�
��f��< N3k�\PĚП�XZiŅ
�A+����mzţ�+F���W����:,�.�sB]�{�5[��Q�߉�I֬j����ä;�k���aY;��~���j�>��"I���%pN�a{*����cҁBAPl�xҾ��U��K�[���r4hmy���F���옍�L�>Cz'��e�2Yť]楡j����"���VJ�2�Msy?ʥN�L�u/�y%"�/'I��tM(�Ҩ�yW_?ds�
{I�dy0W��M#.y�<�F�%�^+�Q*�6�T�܏Qb�������9]���zF�&��;7,&��'	�'��ߦ���!F�����Vy4�.�'[x{D{��������WUd(�'���'�t\\�aP�:�ʐ���hf�g;6.7�h0y�w+?�{`�ᵧ�UhB5良9�louW/�K����_�0'5��2��6X�E�^ ��`��)�앆�Ac@����|��ⴼ��54M$�{*}��z���cp�%����⎙$��-��;p9|橢���ou��~�t�)���mI�E7M뚋�sV����8M����X^I�̉=�����9���a>t�ͬ����xv�mk]��L�[�J�k��m}��8n��lW\��\���FԒ�ޢ�茸K���
s#-�>o{�]��cƶ��D���:S4\��j0!{oe��ά#~��P�Y���Lv�K�w��hu���肈��P����(fd[f*��t�iL�+���� 4l0&�P�0r�Zj*�7���ƥ�a�׻c�V�����?�a��0��Ĩa����V3��/9�萛�1/c���ҵ���6$�<��x�3�t.�0�i�y�ܭ��35� ���|ż�|�*�'�j��$�́
�*����pq߱�'A�{�CB#�X�N�%�(u2x�F^j.�/���/�tT�M��wanR$�+�q�C��&�0�H�h�w��ʣ��`=F�(���9��;�(Y𵵰�-����H\^���H�5��-E�55�ciUjp�k ��/��������/����ҕ�%�q"���2�{Q�<�XqZSf��"
�o�rP��y��^�ξ�] �R�#�D5��>M�+$y�JBlHI,B��d�?V�.4(�C�,��w��ǹ� ����S�^�'�rsɵ_a"��h�jYX�Έ���Uu��n=<1�͖_B?*}>˵�/���&����Y��(
?�]V �4�r����:�NK�kP*s1E�����q�;r8� �}������Ȁ�3}n� �g:q_� 7W���j��+�x��5��7���H�Z{����5����T�N�1B�\����Ѥ����b/����~N˗n��p���]Ǎ��{���%A�#��\J�S~
؆�ŇO�ːPX�BK��C�s/�o t�9�����4�S8�gK�A�D��jI�#\@90���L`�Q�>K]ߡH�.��m��f�>M��`��"���Zz�y֭:;98jZ]�`��<��eL�cH��37�[�ځ�99�u^|gٴ�ͯ5��a`���oDs���RK:G(��H�K�:q�x�\\���]��	��9t}D+{纗���4+'��{����7أ�1=�`��d
�XCO-D�Bl�dQ�|�I���������2�p[�-	Lm(�~IӴT�\L��̊��|�9R�6����B%q��je�\�w�wՂUQM�(��v����ެ-��	�'\�7��Ȑ��L?b�/�_ �oJ͎��4����A���������8הW�%
�<���s���~5��"��pҘ$���'�,Ei����b���̛{�� �ԟ5?�~UWQ�*�5��Q0�FrP�X7Bw����KYkt�A�Y�yA3�Ռ� ��%��hw������Ո�	�x_��9]T�&�u)�xN���*n|��6.��4a�r.�\Ĝ2��.����W����l�����8�����Ok�8{#5�L�,�ϓ�6p!��ik,d�.]mQ}K����2h�����[��!�p�v�`h�d�+��z������~���� [�N��I?������j�51���6��(���WU���D�Z�k<���Aԯ���(IQ�Ak��|2xz�_��@�g2�`T�A�!����"��ϫ5{uƯ&�r�bS�͜�Q4)�h/B�ҁM\'m(PQ_	���*Z�l�(4�Bp�nʋ"�*X�Q�߫���@*�YM����5 靼��*����~>E�&�O�خ�B�t�x�/o��U�&3(��k� �}��d'4�B;Yֿw�:� U�e�C71���ߝ\�9��09�ק�����eA^��M���q=gW]1I��κ!�;��\i���m����pG��Q�p�ZH6�
*Q?X~$��XO E}��c�o.ea]<g�
N9Ј�Z�#S���Ei�J\2<�#�I�e�����~ �ڞU��"��4r5�g�<�mH��u'_7��I�����.����eI�����d�#D$.63���3����Yث�n��s؋��8�<�orY�g��$��BБJ��wМm(|��_�(`���fZ�-2������@6�Z�I�b�~t4Vc
��c��!���C-صP�GF�����O���lh���a�醇�ᶓ�;T.�G��)�OK��栢,�C&��n,�'��:�E���Dw�_;��`{�tr��f�իpX�îhBcUJ���T�b<Ң��cW�z�����(W��/�!d��Rr�}�����RQ��3f��'��{+�U9���Z�QA,�_��A����؝2~����Or����h,�^�]%�K��i�|�Y��s#vuxo�vw<��� Ôvi����0�+��/�֩��=����Q����Kc�G`�b M�5��N�xQ��ݒ**�}�O���JN"�y�3G�ꂇ5M`�9u���T�YT������Pw�'��1"}0�$ZR��o�le��3�fd�/�#�6a�{f+d�;���!�|'�)|�C5�\
���]w��95��MQ'��Jp^}e�����L|�ۥͯZ�?]�:e��O .N����|�a+ւr���/�r�EVL��J�Y���������K U�@�7LE���(q7�9��������S����+Y�k\�p�3��I��beP�w^o9�E����w�ڶ���V���)�8��"n.�mc��(I��F#�Or��"œ��(���d�R�=�)�,s��:����� P�M$��#S�<��E��v�=�D�9m?��%.�I�ڽUp�h�\'�	�R��4ХX�.M5�øk+�+t��7(��(��c�E� h�/��) ���&u����룓� ��|�IU`Lc��!�}�g���=���t��j������È���_��y��}�$A� +�q��;˻�I,��v����a��܉�2�c.�D�;VO	�*�w�[`��>�Nn��?u�/��vB�?%�W�O3�y������5�Š���In����ܷ�0�d���^?��b��`�?��*�Y��h�ݘ�y���^;�L�q�@�����Yns�l�x��ϲ�R�P�4���L0�ۉ8OY%��9�j�mU�	�����hap��s8�!k��ffz�H�L��Q4���bl��e����-��?�N���~鯐��!)�,�s�^5�4-���@��䝋���p�5�bᱜ����ZU�T$���x|�	���
R��#��o���O�q'v�:$���ҡ���\�Ǆv!HMVl�wz��Ĥ��1��rf��c4�uu�� 2��\��[�]}��SJ¾�������|��4M������`T� ގ��f1N�<�����S	7߆��Ɗ�z^q�fH��%Q��Q�^(�����#޵F��0�o���;�����S߉������qD	�߉�F��Y�x��2�����@e��e�M���+�s�f�E.�05�#�Tn��K���I5�u~`���}�a[�|c�v#E@/����������;�w�+�y�zuX���X��3KC1��JR�4(�/���o�y4��/i>틩E�¯�׺M�s��d��ws-4Ev�ݟ$)�/&�E-�j�2�zE�USg�����лyE�~M�\�ݡ(��i,ջ�߅�����z�)�lл�V��wc�s�>%2�V�,/2�#�݇����ƭ���=n#3�:h�Y����$���s2��9��A�k!s�4���%��D���������,X͛J�1���]A�3E���9TVkx��j?�{H���)���&�X���LʣAe2�>KY7�6��'������iG�S����/���~�w�9X�D7�����}C5�F��Hg�If����z����]��ۣ/��=�[���U�O����S�0�V�b&�~	��Se����)��'��ucۉ�8��Z�Wh؎Ǖ���S�i|��w\�� � ���eE�5,�.UR�.�[�<�,O����]DE��FW�۷����#�9��V�LzO���CS���Ok�:����B��ZPj��V" f@#��*7�JGJ�6)&�!�S���s����z��,� ����e5���̠�t��o�f��Q�YL��#��x�X����S�D��T�G�ۯLa�0U�픫Z����י�]0H݋�K���ڒ�<�;A�X�2#t�������U.3)�ҧ�⫑=��3��EA�������B�,�3����b
^�ז��pMy���5#������`]`��NXc����؋�[�a�l�����	X
+�V['���J�.7�Ƹ��~����w��S��E	m��)����� ц�Z;���3���٭X����q�v��2�~�����֞$1����z���V�^ɳ�IDC"�����U,�� ��9)�>�fW�{�pW�q��QZ��PxL/�|N�K@/�p�lo�5L�a���R�e�ݝBrXl�	9G��I�L����>-zϺ(=����]/ ]�������Y0A0|��1Yͅ���,.W9{� r������7��f��1o7�p�hmJ8��
%Um�`�Z��RSI��6���0��5�������N�Z�Q(Qr��[��_���˖LV���f����	[Rт0��Oj8f�M7�h@`ٓ�fc膄-?�"���DԔS�;0.��ښ}�Z�s�~#��f9�[6���:�_͔rK��ʊmE���҈#�ohڛ�HX>H������-��*��4iX;��&_ʃU�6 ���3��h��&+հ��*6�z2���v��zF���aP�K���{{O�� �|^0�x٪T�>'C�۽vY�����v��QG�+��=jܙ�E����<������<�rͥ��M$��Q\[iU�'q��?)>��¯*U=�'k�I �	��͈R't_��VHl���	d��,,��n����x�y:/�1��a�'�fη!�Ė�jb���,���1�LI�Md�AyRw��J�õ�05V,��0dBr����S3��nL!1AH �[J�ϫI�8��$&�A�N��
�I����qNl���"��1�k�z���X"z8��V�HC-x����"��O僲��(���g.A.��[�B�K�i��>���M?�n'R/���j`��e�[�9X,U��'�R\�bN�K@V��3k}F@J�|G�(����ϥz�%u>-��͚�@��*��i��)��U�n��ݤ�u:��p:R�T�|�Fby����M<:�})���+C��,Dd��`�,�?1v�\��L�Xm��D���e�+-]G�	Y�1���0t:q	��eH���t�͒tm��xZl���η�"P+pld���C0�c���3! �]������Y�&�7X�@࢒��;^w7s�ō|���h#����td\�,^"m��hʍg*|�$���(��Jw�@ȣ��`���ЬQ�$8BaGd6%kp1o�(�=}����mq����7���+J�mxa6�葋��=�d ��z!�����AM�&ƪ���_�A#�!H��pK�Fn?.c��TB���'v����-M��L)��'��)i���4�}�w����$�*��3*S��呶j0@�p ��@���銥K��X���E1�H΢�r��>t�A��LFK��F-��+O��8h�W���t�z-s��]�נi��ɇ�}n�1�J�<��I���_0�K���/�]��QU$��8<�}oˊ�&���������u�KVCpah.(5���M��b5ps3r���`Hw`���v#�/�﷩@,r�P�V6 ���B�4"��fJnp��#���j�P�iQ������5@�z&g�J)�h2�̨�>':�j����5�<s��Z��(���G��)���:����V����c�"\͙���<��8���9�� 9V��U�롃�Ԕe�EYO�ܙcBm-�ɿ5��kT��;�غN(Ь���T�N���O���a�y�+�J��'���w�5뾺�{&e��K�
�S��ˆ��'!� �*D7u��6�T������Zx��/�e\)�a0�k�"f�<ɷ�J~�b�c�t��F��� "�WN����5�T�lG��������n��9�5a_X�4����&c��� \�F�>
+\���� ���� <<�l�x����=���=^e����!R9�gA	:��;������d��:`ԁZ�-��_�K� YY�h������|��M��T�5����?��z��B?ko���r��p�0g��,��G_��q���4EQwB�Dh������e����y��eQZ������kU�%�B�>�ŲJ)A�G�0�[ǬŘ����c���汪5��_��}k��%� �P�{�2~��?�]P�Ky�Eu�G�f$GT�蹐�3�2V��B�"zq�1��
�����5< b�cn��%�ɸ�(�=v�8	|d�XT�4��b�w�0(0l ��v�
�ϟ�pҴJ�P��(綋BQ�>Z�4ͱ��".����#q�<qeΜ���fr�ƪE�nN'���}~F�b�;�h��ϱ�t5��tNw?���:��p&/B�߄6�2��lK�n���M	/��{"{��wP�fg�~�PHC�y3�9���/e�S`���3�<8��Š( ������MP��؁o����Q]m4q*�|��Oh�`[�3%d�k�q^���?-�)�݈E@TR�Y�K0~[���X
b Y�&H���_�Xi�����6�(�S�2(��LK(���W����s�;��`a��PM�[=���:�8I�<�]�vW�#��q�AQ�2ȣ���~3����Ү%_�ʉ ����?�/T����>�?����p�ſ;����َ%��5g�;>Щ`V������"�e,n`OY�1P��9o��	�u@�w�YM��Ţ�Ԑ%f��y�n�] �,��n�ӆ��[Tҩ�k,�E���ƣH���^SVW�%��"}���h��z�� �%J"���cnE�_qV��v&ӊT~�v��J����B*����c�Q���#vph�2�-���4�v/�X�Փ3o6�/�L�i���b'[K���.V��UZ��5�/X�i'9:�cj�6]r����rq���Aһ���9:�8�}��J�jt���Vgi��	;
Oe�*[+kY�*�]������{e�1ܐ&R9��g���1�HȒ�������Q�u��^n�]nt3˳�W_��./����M1o����3��($�Ŏ�i3�A��B�_`~=3�*�*�t1��J�4i�k�$��&������&�hB�������	Nj��������mxU���b%&�A�$m,�;5�JZ@��C�F�?l(�����f���m"#�M/�$7�9�v�2�Zj\�7�ȧ��*nF� FޣY*���!�L�T�?��Z(��ۇɆM{�~p���Zs���Py��p�	�m`|�у���;n���Y^E�F��h) |vv��#x��� X.[+�)��X��u������$���韾ј�V�X*�H��f\���*��J&!������'dⵅX4��I���zY�7h���F�Q�R�T�0.(c���פ�_ث�o'Ut�3H��j�&�d�u��ڌ���w�+�^�:��#.����þ�"���YU	�/ ��P��?a��J�5��*�v��G���&�>η��ǃ���E7��K��F�6D,ɥ{��⡩�v����6A�C�;X"}�5T���`��Њ�����f���PI�L�t�\��?X�9�
(3��Nz3�`��H>
��fWϡ^}tm�rQ�QnD17.XQ/W�x�iqp {��x���m�y��Spة؜ I˽7M��	V䝅C=ZN��C~�JrD6BQ���0���������C������p��v>�,d����`���/v.; ��=ax6�a��V��4l�U�tnxkb�]�g�I�>"��c��+*�h���ޕ�u<g�@��o�s.�~C��}�5�%��p-_pG�ό�U܉é_y���ߛٕlk�� ]GL/Xڳ�ƽn�G�^�~G3\N��.��0�F��g�I��RY���a�y�6�r�6��kC�M����������;��L�\����d�\�E/R@T	�rw�C��v��aiyi���˝n�i��q���W�6�Γ
�vg�]0����골��S��ٛ�����o)|�2078��$�kW��<=��A�,�c��i=����u�����|�<���
���v��	��
F�L�z�`a*�t	�csە���\��h�z���3D��H_�Gŷ����#SM !ơ;,�z�{§����ю`k��}s�H>z.�:��% dV�5=ve��C�n���J�!�h��t��A��|L��P�(�{���X�Yw-��i͘����է�'�0bf�E���v����KUG����)��T�ȩ�9E��8�B|�gc׼4g-��Fn���������t,P�1G�TK��Ȱ_��W품���ٺz���O��J�8���&6:^�n[��AzI��O,r��R�U{b/M�' ���`y����gu7GxUc�|@�� ?5hŝ�ZS�H>��y�����Ȑ�'�mՂǍ�8ͭ�ע��qG��Ifj,�����JY|
M�(o`E[��B,�P1Jt��m�	?�,�vm?��>��ɜg�����g��y���@�����2�:y��NX��ͭ��m w%υha.�A�TS3���gz(E�	5Pņ�� �P�>��E�i����G��0�Ùn�6�>�Ef�ɚ�qލ�VH�J*��~��8҉̋�v��L�21 Y��Rt9�����Qz�"�E��O;���&��!yN�/�T]΃��u1i��aƢ/�z{-�:o��3ҋ�؝۫�,2N!2��0{7��8l-c�<�_x[���/�[u��
�{����2���}ie��v���mu���_�N�ٝ��0f�y�\��1׃�=�wBIآ�R��}*.�9"7)�N�֯6Ӭx�]��D]6��)e	_fb|�ǒ�vي�0L����?2����p�wj$z
F��>�^j�}�����Fsk�RQ�Jc�{���q�!x��k�:oi&�/�����'��R�2g�F�H2�m��e��3�>$�܈�1��0\C5�Q	��y�W�N�����\q �2�ݪg�?"`�E���� �Mb���w��	A�d������A��	9&3}<\Ҕ��`���P�`F�����^���&�%ms_x�B�x���9L�Ƿ�ss� 4_5���e���O$�}\4��eH�I������d�Oy�'�A����4�(0�Bމ����,�L)	� =I#�ae�Տ�DZ���N�6wkx0^���w���ƽ�+���m8��(+-_�_�\�
w�T($�Ajk�\b��_�z$�I�l
)k4�p�w{�r�) ��T�G��`��,&"������hRV.vg�m�kfp�P�|��M����v����6^m���$w�os'��4��"M�"{R�G����:Bv�40^���*��<�~?L�)،|h�ht�lEk��-MP"
	�3�ؐ�ʝawEMs�3j��ac�|�% ����A���S88�`��(�Ѧ�h@`P�	<�Q��eF�����I�/��N�[�KZ)Ttљ��-��Of&6�pB�z}v��]���5�8)���c�6���^�#A�)���G���l�Y�#vcMS��*����l�j%��6������tߘ��\q_=���##��Up�7]_ρ}IjAl4�?x>��.{	H�XC�������'�Q㟽!S�ȁ���"�ejŤ�o���1)@��Qz��u�����֯n�'���$�,`ى03�L���{�X����J��f�o2,LH�>Kg�]�Li�ǂ��|L�e��h.�V�XH�{R��s�P��!UM�k�Ӣ\�/�C��� Ǖ�?d$3�L��ꇜ�������.^[�B�����
�k�>�4F	?�O��J�s�-���ִ�,b%�"�B#�.!ϗdx������Ey�%C�am�fm���eZk��@�
-|N2���6eZ���Ai�-�P77���|�OT�a������S��'����亂(~r����g��\Y��8�<�Ahr�����&���Sv�|)M���Ұ~�@ǵ���4��~zK'�M�}
��XC��X��5�%�]KˮH^䳆վ<���c�\��td�Fצ�͜�'?�	�/z�)��Z���-u�*�Cz"�{\�2����q�iS�)���jǊ�"-Lϡ;:�ڒ�!��'����s�@]/��P��jB�&�Zx�� �Eݠ�v�
OM�`�/���a�u���l���!;K��Y���o��um�C:	bH�L@7H�^ x��dʽ<�ɑ����G|������
�����Z�)Z4�&O�� ]�G�w̜档GP�.X8MC1]^vN^??E�m*k�/�����Q~�+;�ϥ_Cy͡�;̦!������K�>�0����".HȨ��{��N( r|{Ύ�j���2^c�̽oc�Ie�j��4Ra�Sx�z�i�{Zn̒'�0ڶS�� J��˲B~�� B:C��F ��]'	-�<�:�/\f��7���6��	�XF�oY���hWh��"��Sb�
�q�1Ǖ�(��UR\>PB8��?���m8C�����l-F��
nn��?���U?�+��<�T��+'T�]_���nɞ���E�7�p�K�p�1�L�|T0z���I��[<�X�e�N�Fv.��
�N����� "�C`!�<�l a�	?Yv�O�b�7�"�/�?�>�Λ"���{k[���eK ���i����Y���vؾ�)��rw�����n�
ZG�`�VC��߿���qr�h�L�s�2y��]T6���?�����inc��nm��z34#O��ù0�e�$�o?�{�%�� �
�X�0�Q�f�r��[��#m�uLޠ-���E���"�m�!��m�u�3s�L��H�d�-�$%Ս��6����N~Py��b����l���Dg�8�9�IcF�ݿ-�}��(�����Pi�7�GڴGM���~03����>������x9���0z���y�"�2B�N�i�Z� �������`�$�
�珷e'�b,��;S�� ��$T.��B::Qw�,���,���wXeCP�y?�b1m�6��5}�8��S��Z=�`��k�sS>�t��Ɖ�W}�yo�3�)u(	ub������ܘj�^4Z�9a�Au��yH��'~�)�|b�S���I˾H�]R�} 3�w|���?�d�΃_�w�^﫺�HW攅m����G-���Y5 �"Du|r���1w�k^�������k�L��GO�<;g�*a`��>��H	)��
���������,��v1Fl�+�$��.�f�ƙ����]�r�3�`J��P���+�X�9u�L)��.�$�[b�}�%vA��ȴ�|iql�#��86:Q�;s7�qH��S��������/X�߭�Y��$N�[,y��!�|�Þi����fP�nt^/���Z=ǟz]� Y�m�%���aYDJjX/`�Q>����t�X*��H:����^�Y�� ֠��	�r��7�4Z�μ&ˤ>�%G����kgb���3�� ܤ܉��L�]W���%]�X��ھ��}t��Hh���_�,d3�hj�h���K-<�ݪΝp���=+�f���I�SG2'T�f>�M��l�k'���w�xߤ���RI�{I�^^-3a���^��MD.��H���Y�Q6S��EŪ~3XőU��䅜Qd��n�C���~��4s5�1�w�~�*�V�VwûJ+�����{���XG`��ly�š�p=���qK;�4ާ�ǭ/�zP ݇��B ��	��u�����]��L�:$	�Sz'�G���H����Md�����5���>�#�TJD�]�E��k�;.^�}v͊<2ZGN5������V0�I�@��o=S�<Y�(������B$�\��').��o�DM�\�{�R��^Ձ���2F�������9�-V���#�K�o�8�,���1n0�4�]�d��+q�a�������X��<4P�2�t6�.�30n}nD��m� �F`I�d�aI��cdi<�er��GV�ͭ��뿚��(��l�/� ��Pq�+�����n����Ǘ�~ݯ���"��S�(j�� z�7@49�X�^��s㟈n���|,�d�g���o��e��3�X�W3�x����kf:-(
��B��
r�)�P�)N��+7�F좆-!�6E�K�Zm~��1�u��cF����ߛps�F���5����D�UWQ�1�>�9� lK9�^�c4��!P5���F�]G?|B)@ XvIDm��,]���!��o�Hӡ�=sꗄ��,�� 	B��U"1�Ŷa��fn�
6�ğ,��:"�!�H�� C\U�~��6p`?�rn��ƚc�r����|�?�����.?�)�.�-1y�t\i�}�Hb��/�P�L�Y�X�(����SZg����3����6�}d��Z�������X!��q�er4f���"��pM�Z���ed_4����MɌ�iN�D�v��ý7�d���P֗o'���T���K0B;�ą��b��U�s�e�'�i�z[�8��
sǫ�,!~�e�7c^�dS�k�1��_"$��
iaDb�	o�{�����f�E���J�S��$ $��`�6�h.7�J�T�A6-�*E�=* ڜY�N�Q/B_���库%�wj|�{3� :L����r�K�R�jH��J�?�v���=�����v�2�kXk�tr8���������C\.�@0m~K	eއ%����(&�}�q�Z{���:���.�ʌ�O6�U����I��mMg�B�E5��K-|���o%k�����և(z������U����)(]�r�2�f�Y�)f���?q�J,Vt��<����b�[�D��[�\�!��a�E���j��j6��w����ѝ�ծϺ!��j/[]��-�=iԌ�E���O����6H�?U4/�⡃ץX`�R�+[_@� v3��w�������Ё�����K�3�-
"��	��ɐ�G(�	ooX�u���?<��rv��E���$�j�9��P�ÄlY��9�M������{��[	����C8q|��m�@���o÷�!Ų,T�<ekb��ƀH�d�����v\�*�K��Eh[398�pq������������UO����o>�&@&�P�E�ɒ���^�œ���]:,
�1��ݖ]߲�(��5X��K�q)����q�6��U6։����?�7��f����޸�EO��X�]�u:���m� I�']�b�b �@�t�ю�`��d��x,֋��]�x�~(��ڑ� ���p��`;2\T������^tآ��F���1[ڷ�pEfX�{B�i)m径��g�|�#0C�֤l�\��� Xs:*A{ϭ�ˣ�"�Vq��M���3z|��՗�cNQ�
�5d)+�j~1��y]���?�[��;�&Z��F����xTc���i��zOz���83���"�˼�}牊��E8$O�g��l}	�sbEmU&O��WA��J�s���d�
'lUkځŜO�G"_�����������vW��[�R��d��&c�jFM���k/�t���v��+��U�u����hG� �g�f�˱x��~W�^�QV��.41ep�IM���dZڎ���60���!%�����b_�p1��ÿ��b �p3�qN,���Ll40iiQ�5/��U���&l�TX���a�����㹊�J�E�5��t��M6�N6`�mg���n2�cM�;z��O��TKef�|0��t����={(-��S��{(�]�� �5-������`�LG�@�g]�x$�#y:�xzhhΒ�.	_o�UK� 
��g2��[w[V�,,�A��	,�|��'2:�nw�� �#,q�t�w�n;,�?А]�p��v�:������Z+��D��ϧ8�{�/���K�>��S  i�0uZ&���u�bP�9�㺔Qi��l[KJoۏ�bϻ0��u�	B&� ~_W|y���9��X���:��M�J�p��,4w�
o�ͨ,�=J }��G{���
�o�1��C�.CӲ��=*��)f��n��4��D^�w�T�܇��J�D���Nn=Ԃj�&j7$ᑉ��<��k[b�jW��"k%������}E�3}�GE1BԱ�o���V��g���@��A�)_꣼�'.�ҫ��;3v���΁c6��w�*�=gF���X����ztO�X@]��c���e#�U�i��0�A�	�����1�1��(W���X,�����{2Կ�W�×)��a$�D�,�͗U�!*���lu�U�>W�A�nґͽ��fN,�/�df��W���*k.�mb���N0���8&�o��WKA��8� rc7[fǮw
-�3�\�Ӹ>�*Yj�!��p|t0���`�a�>k�d|1�ѹ\d�^.�z;���ɞ}
< =	�F£�À��=�f���ɡ2�7]|��=���ǯ>!��*�cu"^ <N݅��q;2�Nf!�<�H�U�;��=�_�I.��ݩǐ��Q�ė��ަV�ꫪ�����>.�T��kC+��F(C+ o[I��FXZ����3���P�w3%Y��ե��S�,��{u1�����쾧����XFJ�\�(����&�9P3���c�(\ݓ:n0,��mM���գ�!����U�� �|᷐3�h���j%�fG�U_��� 1}u�/I\Mr�nN~^[9U��(�H#�%0��R��Cr�r��^��2'���!��j��������CJ�?V�"�A.Cķ�?�(�`$i��J�@-t���y�z�����k����\(B�n�b6���[	�B\���N��nl�^O�xd!ڽ�S�����HtEŸ�j8ۄ�'�}Z�~��׼x��)����J�Mz	iV�&x�o��b�.{(��}�s�8��Ң�������5e�Z�������y�-�8Տ�׽T0C4�I���S��"=Bs8_�:��Y�<���L�Lj%�Y��w��D�NZ�[��f_u|[p>�ԟډ��8|+��}R����]�da�f�\8H�'KX�̰~z��� 1G��J_���f�B#Zew�T:�����{董$F�'���sϚ�[�Ѣ�of6�(���򜄹�u��9���q��K�뿷Aj,��A�8�z1��&n

c�p2 ��ހ��D�L�m�1��>��0{���t�/��yb�PC�5�_��|{�@�D�<ձ�Kb%���l��	�����o{�v#�$�uAx�+���zM����@����,��^�=�����3��V�f����"쟵P�VdxXϜ�ۯ ;�m�6me�&���!ӣ �ז��cQ�~Ǒ7��_n�]E.x��Pi��z�*29�)S{YFtߖ�]�G������#�]�ܠ�Z����	=�#I:d]� *���o�9�r��!�9��W.6{��	Q��,9ʟd)�e�����	o+w��<~G]>���`b��P��M���V���X��'�����˄�=�?��,L����*�d��8E����ϗD���ܾQ9E�yM��s�C�/���!�4C�	N��&��?q��C�H�G�ܰ8�NF1a�㔭^�[y0����K����k�,[T�C���ζG���-�J�ѭz��;l?��>��sQ{r�	�ӵ���z�չYй��#��z�?BB� p���w��6ņ��L� ~/�u���j���f��el0x���A��+2&F=I���SV'K�q��^���/� ��ِs$� ���.c;z�`�'n�=G�3�-�Z#P�C�vA�8��?�������i.h�d�v�nN�h����=�$�{�y�0jN�'7p%?��w��j�m�6��*2�h�c,���|�
��O�tG������}��y^ض~Ҡ�\67����˼���k����l� �;�����2T 8+dE˴@o(�]�V�3e�*}����a���h��J)DIޥ��]��Bf���HWIp	��k� /B?�x�.�n�"kѸ���D�t�I�����I}gz�p:y�t%��&?n"T��59����S�!�D8:��E;d nV��sYIƕ�齳u���|Hlt��`D&�'�H�C��c������=	�+ErX�8bӍˋ�/]l�'�� ����J�4#oOD���1��r���c_r�g�Q�h�vXX\FqTJ�4��8~Vf�&��ŶO� �KM���U=�q�o�k�=ׇԦ�vau�6D�4G�[$�#o@�%����FMc"�3y�we�c!��o�1u?�е�� �p��7�
�C��M�+�ֶ����	� ��|U��o]Z���l;��Q�"�0�"���0wp�Ȼ��4�H�7�,�M��n4�A���
b{���������М쨸�}]���0���d�j�g�$u�\���=���wA ��3xMe�$�)J��M��pa�ͫv�A�FF�1s�����A�^@^qV�����O_-����y3q�����Ku�@�,�X��/����2�������qR���%�
Y�b����:���d��Ɔ1^u�/{o�j1� ��Y	q	����w��$�r�1Q���u�Dhޡ�_}w�ɥ|������n����/��t���5�B�(BH����B�XA��>�_Y�W���A=~�Ts���1ը��b�VFE�[��q��ؤb��c�7\��"�k�:�\�m�ZH-�^����}#Q�1�"w�uϓv��gj��[�� hc��؉�0���A^2�h%�9�v��epO�v��F��Hr��ZGɎ*oz�83���X�_�ĪޢqD�\S�w\u �a��W�1�u)˪�dFQ
ǦS��4�D�����	f����g��H�ϕ��s�@1vcqXY�m���9��<XO�z~����-\��v8	�:s�uu���i�������*�ɔA
boqon�~_l��k1�=�UƧ�/&g[X`�R⻮
�:��
W�Gx}j!*�D=m:S�A/�!��	��s�<��*�)v��f�Zt�iV���B�:C���q;�-|�&&��(�����~\6
��d�{��R������z�Xh�gR��U-m����XO=,&Jl��!.匬�e/;���!(l�g�k�3U=�#�����"� ����c-DĻ�N�+kx���D�A�)\7�����^b ���-���hH9����H�>�ϓ�ƒ�4t�p}G��f�E+WKS�w���6%�|���8E@��8��3�� ,��>�d���Pk���'�e<1��9��.�n�+ǃ��H�ču�q�^�q��g��׮�mbpm-�����K�v�3㐓�ҡB��ʅ˒�\�]Diyx��>EW{Sw�33���Zj����6�;\ɢ�GW�'K�%3�^����/^ӆgX�0��Q���t1jދ`�m�*k��f!�t�m�B4BG�ΧLO�m4ސ�������N�B�	b�1J�5��;tw�[�����f@�9��NQG�JN�T�_���Ϲ�,r�푃���LX��6����:�#O�:��{������}�M���q��Hj�郬Ȟ���&�Tʿ'�3QL	A*ӕ����ޡ��s�y�y׋�s5\l:`q�W�V1_����`�L���#:�!>޷K;���n���q�4��]��5��5�W�{c9�p9JOx��C�"���@��Df�d��%�+����)9�2�F0��M&p�V�U�UO���v��:b�]f&61�/p������C�=��|��c�s����K�{F�s�/��U9�>�$<��j�:\'����<���Av-;~�?�?��Yu����z��v*�fu���6����e�Cq�Cm@L�q�DV������{��b��'�H�'�չ�����!�TW����%�\��g�X�x����s�qTMwe��=�5J��K����:��67�u��)$�b1���
�EK�^�ۇ%۩(���n�/?�O�O�Mf�sI�h(r>��t�g�������\��{�Rru(g�3�B/�Z�����|��:si^�6��E:�$�ǘ��8�hM���}���8�`i�2��CE���~�����;Ěת����R�_$���a�9k1R-����j�V��ju���T�1�Tp���#�ZeW
�K�K��J,D�n�@�v���P�L���c����0�b�҈O��jiq#uh�kZ�efO5ң@��f��O��1UF�	�+�彧d$w����H�#隟&~��eQiL��4$�7��_��Z�t�㳠�<[~����?�Yu��\@������Zf�oFγե>:Ԏ��5�y�?c*�,�����p.ۅTA��z�?D��]�<.қ�� �:��{���I��y�>�O�F/n�	X��� ���2�^�����vS(��!���H	��f��4,��$���r��oD��ܫ�z��¿�Z�`�lwzb��tk�8?����4���w�QI8���_��z1�삘GS�g=J+�N���CmrB��N\8f̌yl�Њ=�M�@}��f,=�h5����a)���x��+i'�W��фOQ ����z	680RQ2-�!�F���1bY�{tˬ�j��$O�<�>]�\���"�G�m��=�cDc����4.
�>?x����g/2x(5�T8��H�|V�T�%-�r6 ��Ql��� s�4wt�2�~a(`��5��2lE��)�9�GF�b"Tn?p�,�����^b₏q�&D�.��]��3��;�1�l0�)��`!�R����5o�=���2��yF��ZD&Zdco��[�&���[�	s�e�j�5�apζf�X��Va�H�-Y릁2�W�E�+ٸO�ND�U�/%l�1m��VG��.NuAߦ0��J�d��h�ցb��A���>U��~���'�����pӛ�)����	Ť�.�V�By�O�	G/z��Q���#W*(�Ou}��r�
��5�tW.6,����笼�X�8����	�>voG�"�	�M�0ԝ�̠��a�Il�w�S4\#��H�ˁ������#OK���ӥ
N���h����_mʢ��؊�I�Gi��u{*�9������05�����?{8w�5) �]vN�Uvn�'
 0Uy�F@}5����wU�s~l��^�^_��d3�Im�-�TK�T�,]Y�\��D�@���x�ie����J����X(����k�Q.{gyN�a��W��49H�y�A-�h��U�("{�{��ko���IW��m�/a�_���m]Sx��¹�P`� $a����
�WCr0)3<��Ow.�8N�7�D/���+��
���5?�wC�$=8�Ez�?�����t�Ŕ��|�6a��.>ٍsQˋ���W���r2���΢i}�溍��.�g{%:F�����?R8�"Ú��s�77�W��xF"�����87`'��d��B���BM���.�Wb��@G:��Ɛ�ݼ>-":�޼�&����8�^ZK�4��ŋ.��ˀ�9Y�)?ާ9��z"��P�1>8J����d�S��yU��|K#"�DAw��e{�=s�O/��F��WU*�� 0=86��N�Z�N�̃/�.6�lv�X�u���O��R��Ć|��!���%~#����[��x���}��������A㘒�M�W����d�JF����`��Iڂxb�Ck�w̭��E� G��˩X�d]Z]�D�Wb��1ܓ�wg���|�q��R����,Ra�g��߰�%,-N���~���Sp�S�y�>�VV7�jW��R�|(\�����Ε-��E��zOz�4t����=
�2�U�qՆAǳw�v쟅!�oL��K	�{uv<���oʷ�9s���N[�g��/vڗ��|~��ՓS˕�o"��4�!ȼД��t����`��6Ѹ9���7i��s3\Ҩ�'3_����7�_mvN�\<������711�s��a_�L�,���f�}%�d�Gd�@+���W�֮#~�9��|;;�fK'���ɖgt���]��[5$�/����>Pw����hU��6�<!��w(��c��Kn%ٔ����B�I\ł��WL��an�I��{w��^�1�eJtC�>Ƅ(d 1�ak"L%IL�rNA�j8Ѧ~mT�)bX)P��P|B�r�B����Y�>�E�q�у7ֹ!_OiW1�ߒ�,w/3��M�H$3���(�$�fry=�ŭ��@����K���Z)�8�n����@�������2�:t�8݌xDK��'Xidq��Jp? �B�����I*�b�\h�������ҒY�xDz3h����D'�w �1��D��e~8���N��I�<�T�����\٪���r�i��\#�,��xgʶvo��������q<>?;��A) J��ݥ�˂E� ���e<4����ϳI:#ՑxG�a�t�=N�7�K����O���7������+FZ�
�SF���r�s��')s2������zM�!�vs���!bC�*+Rx��7�@�g���[?8]CDKU��P	=b¡q�y���"���M�z��ozv�@N�:�5V�'�v-|�qh���ga�3�� �"h��@��Yc�p�v�ˌ�P$bRw�Ɔx��� ���������_?�z�Nۛ�eA
�~M������;)��v�;�ƚ �l���a4Y�'�4�&T�E�ka,8�W��sI
S�����̂&V���I�o�f�'EK,c�+u�\�y�]~�$�g	�ʕjZ���>[�&g'���Gp��7���22����.��z�F�$�W�_1�������?�����|�m�KiA0tB��u5P�p���(S]��"�',����Y���[4&	nګ�S��7���5-�����O��s���?W�}8�����=_�;��o����"� �B�z.��W~�2�;i��^}>I��3�a�_�f\�Y_(aEzq@T�����E*����d� ��7P7�|��� ��vz�(Z�+�]�9�׷��z>�Ԧ�l��<�����;����f��U
5Jrg���u�2»� DL�>�)9�V�~xQp�b_'�=�ݱ�ˬh1�F��K�c�L:�W=�p�Z8rxt��,ս�-��}K!<'K��F`�'�-���=���y�o+���2FF�=H�D4�ȅ�^�k��VDA�����o�,f���z@(_v�j	�
4G��J�2�",f��b9������XW�ǖ i�~��_�e�Q�,c	(�nzm��iO�WY��`$�o�Uf�v%.�uA9=TG���U^)�>�[=�}xe���j�I��xmgō�k����ھ:��ш�&�Q/���`�����W���H�������zǙ�%��X�?���T���IR�V��i)ah%_e
�@Nmh%�1Jr��yr	-�N⟽@ h]��fh�P�2pYi�܂f/�h\���5��h�=��������]Rp�Ĝ��	p'�J�!a*8uu�_y^slEжih��a�%K�X�'S�����.�x�x�+x���]�g��¤4�(=V�
s�3��W��K��g��W�`�]S[���H/������W�>�9�ɢ��D>�$�,�
�����"����,b��j`��8���.F�V�%�!?q���>�����G~~�@���|�Tn��'����2�CϪ�.��+S@Nu�Լ�+;0t����Ⱦ���7_|�����0T{�F}-�b�4kJLqgw�n�A�6e/w.\e��n���O� J��,���&�N'���$tIs��Et�������e�ǬHO���&Sv�sF\�Ī��� �:`�Ew\��{��*��@��yQ���N���k�Ѹ��3�af1!�y��y������e��}yTO�=C�R�<�4�QO�o8�(�0Y�N:_t=�)_�׋����t�N4O�3��9�J{���!- 0�H�b�Kؐ��Ӑ���A(V��;�b+��A�C`�%�]���vJ�8M�d��?u(w���Q`.�c�U�Wp�3��g$��A��魭P{ț�/�x���dqA�©��b�CyC�?V�+������r82y�x�$���@_��o��^��ˆ�h����!u�������UAm{���*�.�8��Z:�k�2]���W�r'̒W�Q+�Yz�_~y�jPވ"?�ϓ��r�sz���jP��79���E��e�|�(3Lw�ml�=ߧ���H�4VTb��3ʬ-w���f,����N����ğ$���p�����^���Qn�&_���5q��")`�@��<�gRQf?"��N��
J	��/X�Ee���Ybz�}#�.Te��
v��/_��̟�:�7�u�����jR�T/5E��:
7?7s}=�<�ىJ�'����;�؆I%����w�?� �df\��D%zD:���]h��j0���\�ɺU�����]]g�}Lv�"9�G(j���`��Z���U�b��':O¿ֶ��`�巺�@
H�0�`�>"#��$�xbQ�|B��d�S���������W?�Ğ�:�ev�=��c�dR<������t߱�
>� ��hG,*r%ʩ2�A�`��W��^"셖	�]
�O |� ��л�^M�|�
`�2g�1\eش�.�hH�9��)ye?ıd���i�nV�� �j��M�f�� j!Y����]p�5�C��@{�����<i�����hA��f�[ްi�溳w�h��ˆC�M4���cmZ��h��÷��:e�W��a_KFk�{�ˡ�j-$�G��C������ ��"�-�L�Pz��b�]-ٲ<���Aw�g�͋���X��^���zϘE�6�r��/� ��[J�*'�-Gx
��j[���Wש�j�}����*�&w�ݭ�!���ȫ��0����T�ᢌ��$㗨_�M«�M�� ����*�&syԪb��qI_�K��^(% $��6cC=މy�+C���i2@VO��v��b)D.�|}yR� <�JVI��,`or�kSG��z�$Y��t�.�������M�M/��~�v^EM~h�����]��0�<<��\�R'X��3ۂ#Q�q�m��;��SI��v����X��+�jz4֡�>,��ҭDD���� ��ؤU�8>�M���V=��\eg��7<�lD/uLy_�J��?���jT�Hu{.toԛm{-%+��K�<Sx|!$(�R�d ���݉t	 h�F��2�
c�Y7#�(����8�S�rJ�A!��
�3�0����%�+�[.����.ft�p
�h���ܣڥ�3�"�CN��WNm4ٟ�!Ö4���[�^��8d�y��=:�<w�z d:���Mn�R��3�6�%�>m���p��\j�w.���X/!NY��#��+Y��H1�K���9���mG�� �_J�ɍ��<q3��n2��>��û��A3�y���:��!6�ۨ"��|��k�ܶ
wW1�ĉ>O�1GN#���rb����k�6�ɳJG��N=�°��,�� ���#��U�[L�+���ˎ͜�.ֆCfPjg�V�[)�����ئ�M���b=��Ap��\����λ����v?�"�Q������2��<�E'y~�;8��,�����k(��z�S�\�͹��T�w9.�삏��XI�EL�t�(z������ï�4�uŁ�H
c�I�>��Ħ�ĭ?��( �Za�#j�L�����u���^4�'M/��6���Gȟ�{G�T�"��#f22�Z���-9�[Cx���Jr\�8�;?|�_��<g ��w9�^�0��{}�ް{����|N�a��ۑ���ً�Y�'��B�P��' ʮC���O%��M�l�(>��.F`�R��N�Qd)���u,�?��A����}�~�h�@Lr3�4%��I?��c]£c�^mҾ�g��&Os��� ��{;��N*K�6V�I@8 �OL��ފ���!�nֺI% N���l�X��?�+O������^n8�V[�/��%յ�5J�'vC4�Bwf��'��c}A�;�:�Z�l�9a�?M�hV$1��?魌.�T}��	�}�o�&]4�~�}���uu����ʷ�YY��8���9[��{��k�{d'�}y���N�^S�U��?�c�[�<*����Q��`��y�棕D���&�S�*�)���W�&�g��!��*�pG�6<Cl1&h���w��#Ga��׾ا��X.y^-�I��LǤƾ�X�׀��@����FN7,l/��������y��2�͞�8�`�
��?�U+��j^�[�G��~�d�Ė܁�ڃ`�݉���#
W��I�B����l�d꺷�إ�-�)K��BU(�rx� ��!�[��f�e�c.�XJ�GKEl%g�Q�����%E;������M{�צwY�Y�7� _��t]��������&�Ľ�����Y��#�	��%rN_<���]��:�Y��X9�ǪJ�e�K�5I�J�lXb3.#ޟy�)�
�S %�r�
��!qjLH�v�3��v���k�\b\����[�Ql��m��M�^��o����T��QN���6��^@�_"�3茓5Y(���x"�F�n�������)S��*��w&���BJ-H��)|�^��t\:�!2D�Р�K/B�L�4��F$I������iΣ4���~kS�m���Qv������X�i=M(+�z��C镧���BE �v��/�(�����DO�t�� K���Z+�1b�^������ ���;(Q�xy�6j�����U]
x��у�r�\��ܫ8e=$��ӵZ�<'�Wf���W��mqώ��e�2%=���n�M�@�B�|y� k`�B
����UmGru��0�fKvt}�s�MT4�k� ����x�S�d���av�=�E.��#ŐF�%�r��QH�;3�}ݓ�e��A��I<�p3�ӛ'��2GP#�~��D�z�/ �,"�hD�$��=��p��Q�_��O)��f�%��^|�be,��a
�-_���}��_��ȏ:M,\اCa��iv5MS�ǈ/.ÛC�m%n�.���ڨ��^6)�r��rl��Fm����e��R��:���㴀�o�H�j�%�X<|�|�B�)��?>��l�Ә�k�@�x���פW@i�Op>3�']�{KƓ��>uX�pBxG�nI@���c�#�ɀĒu���t�"�9� {�%X�4��C�@�T_YF��3ſN�B�#]�!G��~��7*�\��89rA��,3B�����Jh�j@��C�Id������A��R��%N��m�:z�n���*�\�<=�;>��QvT@��j>�QW�y�_p���\9 ��	���>�L�LC�}zݙ�3�J蘵�(�J�R޺�Ғ�O��ېa�h�<3�Q�S���E�V`^/�-��� �F�ElU��n�$����/ZI�%�e��=U�i��-u�ŋ�HU��&�M��K��K ����~�wW��:-�I&mɣ�~c���T_%vBA��HK3<|�Lyx���xl`.�3������zJ����+pŲ���$�s�ޡ��M���z�ݵ��ךRz3��KA�bq���kȶܞ# ���B��Qi]��Qz��ң�/v�i��~暉|  �����؟_��O+�Ƶ��!�E�mbTq���ތ*<\�-���~���[��ѓ���+�Ѿ�O������Q�(7"�y��\~/F��I��;X(���	�j%0d� �[d��GA|�~a*�/Ch=�r��8�Ih.�:`�5��X/p�g��]ben��M=7���V�&Cڤ�-dӪMm|��V�+,�N�ϕ QW���r�f��7��	�	�2tċ��m�-P�s��ޢ�T���m����G=:g��*�jC9~F�����3�g��W�	�>K��ur��묍 \����i4/��R��_�P����v�^%�u�K�<?��«=ٯړ�\�5��xB,�n�9��R�R��HW8���A�_I
NȼE��P'�b��3�oiu~�S�p����#��X�m��ƫIݨ{p�Ӥ��ԗU��y���u��Z:�۸��kJ���K���� ʓ������`�{͞���{���+0ں�|G\�Ж��?W6�� ��yh�9� �	�cmbZ��0�Jh|�6��/`�Hk���ΕX)4��P N�>q��f�6ջ�G�߳8��  �k�L�^�O{ �C��n�~Q/I �Ģ�\�dm�7I��a	~2S@�p�>�
�?�e��z�E<��,T��Ap���Z\���΍��5���m!�h�ӽfT7������w����S��ߑ�Ϡۏ�`Zj�<1׬�`�w�S�O��_ �H`u��h�,䍓�+�jS�vQ�e��H�mG+��ڙ��.���Z��/{��a�����lԡąn�F}�1spQ�Ꟃ �a��e;,J''Q�G�����m�Uv��B��1<���O�t��?��J��h^M����"��;6����r��%{�2j�A�^^�����dk�?�x��pM*��A�YS�������x���p�Bŉy+�!HO�XH0m�b�Pp����� u���g�*�f�/�Eʌ����]��E)��l
������;T�w;q�N9|oZW]��2-D�\�؄�~&��h���e>��);��z��i)�J��O�U�ŕ�4��D�aX�A�hb��7؆.�q�sc�H�d2�x�P�y�SȎ��9��'���@~"�����A1%g z�%��i�7�"ʾ�IXC��j����|[�	�C��$P��>�k�z�����@?�����q4���3r���#�JBDs!�9���5�!�c�`|�Ø�#�)wcoֹ���̓Z�F% �>�`�2��ގ��j��5��V�r
����A^�6�z+�������)�=������s
����`P���p���=�/V��nwW�A�@_�^\Y{P�["@��c���}x$��'-��
ˆ�y���f�~�"�m�!��_lT�� ���jp���*��Bߘ&v.��B}h?!���i�n����cR^�W�d~Ϭ����-}(�X�h���3c��pm���)4���b�Ԭ.T�V��l��}Ã�hD����% �;Ɠi6�9���~�������ǻ!/�>�� <�;Րn\�^���n�<q�������x/����#_��#�-餗k!��D� 
;�s�	H���o�9����lJ_��j���|�(&em"�l!�ݡ򀡥a�b��i�&�����=V���
�0Ͷ�]����0�e+Á9*��v#�/�k�f�)�2�=~q�y��׌������H����-*K_GD��Ǵ���Ȋ��R4��T-[��@���\�k����Ǉ�uU�wO,z�ͣ�F&�S.r	���x���R���~)�#���σf㢔W���r��P��α���[YMY��t���;�m���@OrRp`۝��NCtΫ͟���=�������'L2K�{۟��g���!'�W�&��1yE�V]2����6�x���9S��vDz
���:|P��g�ک���Ŭ5�%E���b��s@�)��R�����83N'��u�8˱~#iy�2H�N}�j��%�8��߃���T.5$���a�>�~�*3q8�N��$цD�g�x<9��+��k����,��,pB�~%��fG=(U�R�F�&���ƅ����n������_Za��@Z
�*�oU��?8e��l�|:5��r��3/�#�yxрϗ�J�sd:��s�2�|S�;�`�j0M
�g_�ar�,�9��̯8�`���/�)�h���-�N<-.���`�-`g��C��9*�J4�O��U���\Q��|�������Xƀ����݂�|�&R�%QY��
�����ߵR�����|��px�rM^�4?�m�x�f�G]������l81��.�4�ؘf����Z���x��UQ���8���L�^����2��)����p��݀b�lVR�`O\�n�-�S�n7_�/�u�y��U*8���p���I��}�3)4�-�T�ۣelRuA�����#��z�}�"�Lo��:�-z�L58zH��9)Yi�[�)͹)�J#��MR��Ĥ�\�=)��6�k8Zs�H�͈��'�6���@����<�*1�<��q�E�,���4�k���]��lr��V�^(N<T�>��&�[Ne@�X/�gjKV4MS�r	x�G��Dk�^�3� kYgƬl�Gm�����Ҽ�������E��"��A����ŠeS*�Ə��b��j��5o�Ь����u��y��z)��mu��)��0��#2�u�lY'���Zh����˥�MB�� nA���08�U��3��F��!�`	�br�ڝ����_�:�R����Y�󢬱0������%ҁ�Nچ�?�)w"�x_��fPh0���,8h�Ճ�da�պ��a�]�(K�pU��}W�?ş�p�ӎ!uF�SL.�]���4�e�u�L���� �#E�CtMQ�&�e&���'N�Yjy��������19MP�E����w~��0Z&�t^��l��>�ݦ��&=�-�Mp�k�}M�\9r+�N%�t�ߓ���4�%x�����b���`w7밍����GQׯs�{���8}y钖6��K�5Sh�͎o����� N����*zW�Ҷ3V�	�6򏓁���r7����_[kV	��tp����k���"�]�$��L�}U��+,�	��g���v��C?3P����
��[a�m�Ή6Nf%]��"��i�Or"�J/h��w%���t��bE�)�av�m�󊡵�0x]�^ �,ԩpL�s!��ş���E��e�tu9��t�rg��~��I2K��3��V;�_��飨ŴI��&*����sA1��*�؅X�n_ ƒ>F����b�u8.=����a��[6�_���q��^P{�.#$Bq�?g9b��c�R�xFO�dŌ��Y{�\�8��>q����%�/�t8�Y?J�_��)�f�:��I\�ŧo�.�Z�Q�}o/��d�T+	5qF��s��ui�"���\h,��/PL`��I�\���R���+uC {p�$.m�;��@�h��	a�]��h.�t�lK���Ap����&0��Dޮ�,���F�+ _�U| S�d#64���]�b������ �s��n����7:������z�l/V�[�i�YI���ST��ះ�M��`Vƚ��WyV��9r	n,w�%`1I���G ��-M�'0� �Ѐ�Ud|�*���Ѹ��}���X7��n�Y�wL�D���9� M�Rc�e,?��[bI�$���b����H��6y��5:}�B�I�5|\ so�A¯���Vx�zu�LT�\a}�j�y�DmmE[UwT؉�q�����m�=H�k�	��HJT����C�:�mjn�K\��?�e�e�5��U��&)�nD��^N�|_M��U�+3K���.oo,�A�pI�Y��0���#��U�_�1S�$�<z�r�P������"�0�ō�@�|8���s��y�@��N	�����g��L��#PB���-�AVB�v��b�a�̮H�i�� pt1�g��d'�z�o9rq���:���E���(�;(�h�����M����9��r�F[�XhIݥ��~�d~�J����yo91�]�IYF�%�]|��uO}c�/��So������5�b	�Q�V���*?g��� ��X�a��H[��8�H.[��qc|�e.f,zWߘ��DU��I����7L5���5��=ֳW�Q�w��{Vy��_����#��S2{*/�����V���0�3���1y��Vk��v��<�٤B]:m��o�ˑ����E5�e��\��/O������zO�dc3�cy�]�e���)�	��ݟD��#@�l+�tu�R�ԍ��҅<���6it���t���S��xaZw�ֻ�;K*(����Pɚ�m%Y�𝕐Y�����O$9�1A�U?r���U��+����_���E����y�Yܱ/q2ц�z�	e�W"�qb(��|�q|`m���)�ң�����@����z;�ե��ݛ��і�YQ����z�gأՠ��Ё��0�C+���m;g�d����)̦��U�B��wg_��4�?O=O�Wx����?���q��T�Y:�rP:�j=?���p1QW�:KԴ�ߐ�4[eģ}L�[
`�D9�{b����D+�i)�K���А ؆�O�G1�-M�P�	RŮ�t̄D��~6
������Ҷ�;�@&�u��D����g(6}a[
�v&"e���ʓ�/�U>;^}3�ݍ>�ƀ 2b>%x�?tK�6�o珰�"a��#Z��M�U����ȭ}����'\�S+%��G+��j�p1�~Y=��!%������B���RZAz��
J��l?$pH�J��zV#�C|C,�>���5u�~!�JcN��;9D>L�3����*�SȜ��Ͻ�}[vc]�|��e�z�`6E���-{��/�
*.����W�	#�)"�L�������v�����ٿ�3RH��`���TJ���>K�{��wl�n�4В�N,E�n2	[�Q�f�RK��	V0+�������V"�V~Ĕë��WkWgh����F�:��*�`�ԟ4W��'v��lQ����C[��nx�-�ou�P����%�*����kv\'���5�_�M�a�	��X�/�.�et^#���'�f*�  �t��놸�l=��h�3�����-�	:���n�1+b-{e�	+�ӹ��|d������é��f��9��NDδa4�a��_��zT�֛�]�m�"7M`!g/�d���27��A��`KLZm���ۅ����}+����D���VC�PlA�����O���PI��k{?D�f��,=OGؗ�h"�iu5�s�ߎap�s$�H�lZw`6�^ᇋ��ٿ���C	�AS�7-�3��zq���İ��iW�U�F�n�Y�\�)�<.y�6j*�x�Y��ٷ�K��9-��Ǹ[)�d�"�|��Fhn�#��ŴA���D���+�k�ˇ\:�dAR��QoQ�s��a���a�d�d�j�0S�c3<��#]J�񣖕��D�^˝e���̏6����-��y&3�[��ھA�~����	cߤ������ƫ��X��A��	��)#������yius�'�@6>�RA�$*�g��7����
H`�C0�@�@��|&]1��*�g)!\��R�Bcq��+X�2���Q�Ox�a���Jd�	/���Њq����\k'\^f��+��%������
�0�TgX�(�D��a��P�{��X+�Y�vEp#|5�����4i��&eU��rv*ʍ�m�Ġ�G��2�߃��qp�!�gNt&U��_N��q�������*G��a�^���,{#��C�-��/�K#���9w��Z�����s�:~��U7��bI/r��T�t�k�8e3yq��2D��і�'������28�6�3���V��/u~.���Ү�v�9<|j?+���s�b�/��{�~EqC���}�)t�ⶔI�*Z��26�M!+���.��Ħ�����z9r�]Dլ��*%�S���=��+vV������0]��V���{�t.'�����]j��
�.�U^��9�ױH�N�45�2��Q���u��M�4k7U�a�m��ʦ���:%����}n���坍�sN�飂�Un�B F� 4�RB��ͱ˄V�#\gc.�����3�B�J��?6�N����PG�xo�ݠ��pȡ�8��.�[rB,H���@���O(�7�����b-�5�
3x�l;��l��������W�<�K���,������O���\��k�ks$W�Gr88����ewXH������u]Sr���m���ϙ���$.!B����gku̨WU�ArI�k�!�Be(�:��:��ȵ˴F�կ�A9;\���;!�T%���e$� �,����Їl��x�"xw�U'y�B��t���Q�yx�� `��u�N�0W��g�5��In~��S�i�S���*"F���������D۶2����Y~F���j���͢}�(��	��hokq<ؠZQZ�'���!N���ӊm�"H�Q� ��ԅТᶕ�F�SVJ8X���ob�2��C�-�g+�,�{a�#aI�4p^Zm3��k���:���𰤨�/J���%�b0��?-Uʝ�Fm�D-!e�l�4��裊���c�ި�&�rMOC��,�&��EJ���acV��u�#*c���o�����_��g�D� �'|�u�A�͆N�P�,�\	䪑b�ZWx^	 �t豸Ick3�y�
�����)�@ͅB�_�H�Fo�s�Zo���A`p���1,��$�:P�яIC�����؍�ԩ��O�-��B*�4������(X�������ب�CϘ��Q�����R�ݡ��hA}�<srL��Z��/�L��#��e��aˁe������0�|S/��"Vm�s�Q&��=�w�m���$�h�Qז\�Pc�A\5��{�gqm��=5����o�Z�ښ�H:��s��4�����;r�t�&�9�L�~5(:\f�L�_�@���ւ��hEw6��½2e��_��ڲZ�!��r�O2vi����bٚ��ǧ%LO��ˑpHj͐�͘��ιQ������5���Pg�w����<�1D���1�.
�J�Uz���c�r�-)S��,�`J�!%tA���&���˳�Ӵ�����w�cL\��l|K�a����?AX:��3���J�r���	����"ьu4��ٸ�hc}]�4�X��RV��~��&.#�W϶��у&ohr�@������A��E�`"�9 �0 Թ۩��#*y*#��1VRi�l'Sg�S��4S��p��%��H�ư����4���F�;>��7Ic����;�S�'��V��D,~9�_7��)��������.�]P�3��9��횞�G��2����f�-L�8GDo�D�I\����4̣�$��LP��}7�_���6Um��RuI%n�Ĭ�M�AP���x�U�0Na�$�I�|�+��T���t�5��Mm(�����m1��ȟ���Jz�o�S$x�Q#�M�d��b����."!�b�:!�t�'��#�{,M!���k5XJ��z��f$�b:�T[������W/bX���Ge	�� ��&S�S��u�ԏ��՝�@*��-�b���0I���Y.V��|�q/ޙ5J0�qW"�z��(�����f,�&c尢��2K�)�q(�^���&��fY���]��_�;���/�鍣u�TE�Kk>�^��S�AT�_C�����<�A�U���,�^6���C ������)���D:���sJQ ѢF#�a(�_���hej֗�)�G7	ؐ��#����l4se,Z�<&:�:��x�X\󨹍��Vy�N����n�o|x�╋��^6�K,�;����F�S�����X�ø>�"O���OA���N���gGtL��Z0�*`�{�M�U��ΟE����U������$Pr�~���4���v#�� 6{����8-�Y�F*��(@aL/pA���:��d�:�9U���_�[o*��	���/���}�`#�%~�,���3m�@ਪǖ��yĮ|�w���OP�����#ؿr����&�,q�bf���|�1i� �����O��r��*��	dv���;��ǓE�Yc{�	)Y^^��$�����X3)��ν�"ɦ��9t0���iN:��;0^�f6k�?@P�	���KB��L�&We� 5�yI]�f$v�*�)�����B)��'ھ5ed��v���+����6�/K��#�ך� ���'��]n`��)S��j�����+yR�6]t�l�߅�kKWc�A��l�j����Cс�yw��B���7$��ߋ���(��ak��ZE����������5�6A�kaV+Fo��ӧ�!A��F�74�x�J�?�"T ��P:��k�M�.�7ڤ^n�vws���pѾ���Dk:�oe�S�b�
g����T cs�B8���߷eU)9��^��U���%�8nE�T~K8�sc.c��2C����D��i��	+��L�=2��O=���M@q�#�z�_�į�sj�]��T)��b��%�'E��_�S����L=M�$�w�5�'#�2c;z���qY���K5�q8٫m��SNa���W�@�)�>��UM�� ��O0�SհK��;+5��b�'ޔ�	T]��sΛ-`����.��:�XY�A��'���x������k'�	b����R��4J��(?�`�lʎ7y�)Pi�aq�9q�����n߯�S��[Vz��c	�Y�rm���|�/�
q�w�ٔ����p���kRK"���0j�R]���[8��1��5\5�r9���� ��8�{�c��xXS|2�>�*�"������Mp�����n��rꝌ_�)R��i��9�C�-v�<ܵ���q�:�lq��)jlLU�W)�ٌ�!���I�.-B�a� �d����kf���c���V@��`dC�b�
�k0�^Y���Kj���~=t��F�C���Bլn���ˁ�.W�-����t4O�kFS��-�ٝ��f�|�ܳһ/����J��2D칋�4���d&���@�&����=�4@)��/{��aJ��w� b4�>7dgd���ڿ���4˨2:15�K��l�XM	��nNP�w�В-D܀!�eMZ$���ї����]4�u<ʏ�ߕL
o��������o�.Տ.W��ZMZo�Q�Oj����qf�#����4v�_�5�A�°<n�*�C����& ځ��\\��\5��Z��Hq&�#��ӂ��l��S�+�>oŬP?X;c� #������us�ѱ�����nx1��}ݾw�TX~��Sg�ÍCc3�;���(.)O�՝����a�Fn��&o�U#�i���[�p���[7���+T�x��|Q�`l��>*��W�^�����W~8����>�ql�D��`�m��������B�t7�Ҧ)F¾����&e��l���� :T;X~��:��-���'��rՓl!m��$suX�ӧ��2�Ӓ���jt/���O���E�)���ofYM���s�%�M�׷-�R{�Ar���pٰq�&,M�L޶�Ҵ+wq����5@}~��zJSKgqŐ#l�G�T����lk�4G��@롽�{lڤ

ጌ��|��l����J~d��kK_?Fɠ�M����n�%50]���J
*�hQ����[��`�������,��`/���ɽ1�j�~���}UΘz��UL�H��~"_g�b����Aq��_�h�m�)O�ZCr$��W�l�6�¼��#[�J�(B�P&,��c�v�nEG@l�H��1:DvQ�������&i�+�n��UH����14�������_�xZ[�/MO5n��$5���!ڌ���3K2]��9%����=�7E^s�4��x���࣠*�#�|L�I��.�;s����f�X̞Z�M<����&�u���E�t�[��xh/��_:?�*���'>SW��1�)v��cLȑ8��es�22R�z������e���J���Q�U�qA�������b��6��΢��)ײ�;��o��������_�·eS����)H�8O�!����MN��K9�t06�ψ�D IU2Ě,Yi��>ʅ�L��A�j��t؍��Q�,���>�����˕��@?�Q�>��<6l������뙭|\�#%��KH������t�:~Mx�,4�{��[��%��BH��|n�<v4� -�_�x��t�{v��N1Iy�>1()��9\�;n�XM���Ilm(Pj	�-�+�R��^0����}L���[�o���. �����$8 '�ݣ���h1 h���SWmRZ�i�3����.	1?�����?�OG�p >�V���	��Ա�U�>�6��H�_�?٠0��A�Uy���)�����c���s.o"w�L.C��� ���F��8��1\��-p͊�Ԫ:J���;��`&7����Xq�^ōX�ש������,�3�u�gca�N=�%%hg�0�P����3��i�����h�\,G�P/��CJ���.\Ή�FX��B�sX��J:�J���V��ˡ�����	o6q"rG�w3��|iR�]�.�����C���B�
B�|S�l<�'WRAEWp�یڑ�j�0�a��s[�EQ����4���ψ\��E��K#6��2��������)����J1�3��\?х�����5Cm�y�����v�LSE��2ub��Ϧ:1L���	l�����w�ԙ�V����as`Zҿ���K��kcXd$X#�@�ʚ�G����H'>�]�O���9���c��Z`:{�(�8 m�4����tO�����+3Ψ���2�%����ߣ:`�?��/e(��C?4�J��*������(�p�XQ�Ny��҆g{2?�S��Tן�N��b|$_O���H+��ڽ�x�e���s]��l��*�i��y&j$��٨Ҽ4f6��M�iP�����-̎r�i%��u)�Z�I}��7C�mTf�-�;&<���a"�E��,7�݊�Fw &G��Ty�g^�N��eQ �뇮��,����~�i��{,�;����ݧj�i�q�"x27�<�\�8�L��������|��s>L�#�ؕUW�L+V��Rpc�s�D {���
��N�#�F���%mf��v���Kd��{�Խjt%C%�9;�0���?f�������/y��2��P�<�l����t��P��r�� ���n�>�G�
È��U�����V���Hr������9������4���:�-�z��5?O�sV��+�`8j+���Y4ם�ZÒ��V��9��IC���y:)d���[8@ാ� �Y���Ik�]p� ��Lx�B�N�c1�kf�(��h�`<��3`r
q��C{>�������������2��@�3���Ɔ/�c����Tý��tZ)��>l�)���5K������t���S��v����ߖ@�?Z����@���T���<���ٲ����k!n�g�(�������I`�<�_��?p��hP�	��_i���aX̾ʸ.[-ԣ@��i��Q�������s>Ԙ5�b u+��|T�xr-a+�VU>?}�������`�[*�2��`\d�M�¯	���&��2{��@}�j����,7;)��Џ<	$jv,ɪR[+�f�d�G� ���<eNOA�#��*�}iY�ÐAU(ᡎֆ싳%Gv},K�I�v�I��� ^-���/׏6���~$����C��ύ�<(f�/h��y��Bܕ���0Z$(�	`7�om�)Bv?;��%c��4��T��e��$v�w�E�Ї9���������ė
��t�����)	� L�f���nb�\��E6����g�*m��i2Z�S�� CQWo��Z�0�h�O���z���E�$B>�'ba`��k�&��z�q-����{�����̵�M�.$�������X:�����^�:}�-�FtG6�6�|O.�JV�����mo�V�/����#�U% ����Q@E��A��h)�D+��}��f��EGӬ\����O�܆\��-�f�g��=�!�L�,/Ɍ���(ס~Hf��+��8�;1q=z|��OtY�e�b���K'yf=P�@;Э�\��Ԃ�+<'��ϰvC�������X��Ԑ+]�ҧ#���e[�b���7h��rL�<�W��c��v����gz�$[�eZ�b����Z����+�rR�]��.�l՟xh)�Zk���,n�S������֗8�k�H?WEl���]6p��W׳�̯�w��i���c]<R�g�k��� y�>�|�6�g��Ĵ�ጹ��_7���n�V���I�^I��N}[���n݃�j��5�J	���a �@�K�Ό pJ8�c��7�A�(���'G6�i�_���g22�>��f S&��]�S�y34S׈\�������M,���R��bm3�a_�W�C�q3ܻ7Nd�.bc�4�?�)�[gy�a �Ⱦ��V�l����_�v�;!��2B�/ڮ������?:|ʼ~�1�|�
�AY:,��U5�Ǫ\IZ�P�D�x�|~' �̈́{�"2d��(϶���G���i]��}��5� N=z+��K�l�3��s��r^�M8s
���b��	'����"SWt^=�b9�p3l��$�.#x҃K�8����ͭk�UJog�=�鵼)U�,A�n�P��޽��jq�� �"���̓��	��Z���yu� ���n���V�� ��ٷ�d�,��k]��Ly��Վ�ಎ���cG<�fb��fdY9_��8æ%I�7�^��:���~Rm:�{��%f���>�s�q��]�u�x�M�ƕ�5ngb�'�]��&v�y�M|೔d���؁E:��n����%�1�*)�U��KS1tYډ ���'v���؊�8"�k�(�xb.�Z9�y�{�d�բ-�>Z+oP�n� ���~�7	������+I�PVa�w�$��r0�29���9����b,��������z�N�� ��R�.OY�gѪ��E�4��7�1���'�I����+Qt��0NPz�K�5I���_�K��a�������Δ�	���J�a��wT���L�mM2����z P���k����M3�.#׀@X�K�(�q�H�f/��A�Ain�to,>�q{�f��*��C��Y�Q!h*�Tx1�6CE�@�\�����$�<K	,S_;�_�j��X�ItX��|j�-WF�����|�6�b�}Zv��~MR�o�P�̴%���:�YUӰ�q�}�ɜP�J:C��t&o�(Y�_�Ի{��5U��ەS��8����V����� т[�<�5�w��U�I�b�*A(�ϕ����`��z�c�6��w��>��=��_��ܛ%Cx��É��*�Sޫ�Aot�n �:���ۜ�J��p;�{�:����;����zcd������+F����hɚL�Y1"�CS����@��d�������.+<6;�;���`�-��r��/;�)?�	8�I��XH�)���M9Gb��y�(z4b��	���%�����;X��V�@8jȅ��Ȉ:!n��䘬 '�p��:�������w��[�?B��M���Z���e�M^U�d��^�gN���r]���@�s���k-��3kW��6M<ݛ\��J=�W"R���!�{����ʠ�M��s:!θC��NO	WhtR3�w�<���_v�g2s�&��ORyjg�*U�l�������d���L�I��74����6�ݤ�8�V�;+���$�@r��[�*p�U�\��� �½a�����^i��0�A͊��${��1$4��"�I��R��	�Y]� �hv^��Q����-v���H�E�@�ٛ%�6)�Y2GGݺ�%����hQ��Nܳ���Rjn��ɧ��pP�/2���#;�B��S�q��BE��HA�c�E�R�8���։�ઝyY���I�*:n�d'��0��D��x8�JAOA@S:N	tnmg�A�:H����EG�k'���])^�7�(o ���aƓ[��%Jut!�g�x��XT.]��baY��a����$��O��_�hVVW��L�<��Q�٢���܏�~{��:�_�|`m���XǠ3
�][� jH_^$�}�3޸%���G������O�	Ƨ��ILY0�xg�������L���t�'��u���\ž��kiZ�c6h�ވsF�s�������zUyh����xE���}�!	tX('�:�DƹO�XC5,����̠ ]�����)V'�s���yL'�u}�WRʢv����A�i�ŤC��k�XI�����y9���|Ք�8�N���i;��iG2Z���ao��!u�����S���a��>uo>��)D�r*�H�Ȕ��+ϘZM1��@t�᪸;�d�l[���CNP��Eg'�;G��>��A��T���nKd�1L�KBmh�����q��
����w��	P�E�r�:�E��p�����&S����ߌcԅ�T��@h}�+���#0�c%��gov��{S�50m���#�+G%��f���Gc���-ś��)�X��F���+X�l[SQ��q��8{����7�jA;����!�����8���1+�I��� �� ������ X�
β��*�<�E� ���,( ��\׈&�Qyx���mBAE��was]� ��ve�4�����]@�q��UY�8um��פ�O6���[2O#��x���Oq&ͻǚT�z����� &���*�t�ue�
[��Ǚ���u5}��Y�b�IY0��Fқ�28����呰��I�V[{u�Lqr���ICs�G��Y�i�`~ٲ'�A³����.�-hDc\�F�u���{`݂� �>�ѩV1f=�y�v�$z��C�'�^��d��eB��]��a��HY,��J��S���Դ�|d�����*/�JN�-�m/���x�]�5)���}����k�[�o�E��γ,���Gۈz*�O�8��(���솥׀k�ȤB0|.A�rf]ɏ��h=HKZ%�C.�%#�ӷ�й�	��V��pC�ˣ�?�]��O�O��?�$:4x-g��@lN���9�&!<�O���t���E��#CңsxZ4tp�灭�ƫΘ��E�r딾Ƕ5��i�K��!q�c)�ە1��O:d5"k�\�S�ɞ��H�g̫�eʶ�����N-Zt죍�O h9��qn?�e^�冢�x�YC����io�hfr�*�^�VR6-[�y�^�'�Q���ܘÛ=2�D&|��k����v�k���
?͙���͠�K�F��T�"]���&�&�(BO%�gw���]��-��C(�W��s�>ީ���_��@���+�Q5��ey�Oo���D��n�3�P���3� �qKǧ�������K9���uS�vG-�Y7��'^��Ve��>�'7��ǢJ.CU���Ms����M���񓇍�6�t��&R��1�#B�"�6����q!�z����c�vGq�Ϭ�}�H��a�;��1Rt�]>f�=M�M�:O�P_F$yD�ڥ-Ȧ\���Zҿ��BmW&�G������,q�;�6�x���u�)��(����Ψ>\�B����{ �������~S���~�-���5�������r�����n��ϒ�-�����G����#�y�Zr�c�[kk=v����*��u?���l
5�'��Fy�` �e�?�[��Z��;s�`��Nx��R�	5���
�Y�ZU��� faVs�k9Z�����Y��U��B ٥��
����\�M�\�/�o�����^x�s~8�9�6F��:]�IlF���&�יּ]�Rn�$Bd�e&���я5� ;l=ե�ע��^r�-B˼z=��G��0֜wg͈��0�3#����'$��67�j��"3�&g��|�:��eO^��v�	y���ب5m�5.���0BL{ib�����_�˰ �cU�UXP�]VN�yљ�zUQ^>!-�f>{?=���oYg�W�����͢Es5��~�*��Br�`(S�j'�l+^
��=�1����4���$ͣs�A�V%:F��A�t��KP��x.IA�\�պ����P���9�իj��*�ʠ���}��2��W!`K����d��Kq%f�g<��q���N����UhL��V 4��>k0�:!��[����⾆]�� L�!���y�]O��S?4_	n�dѿ ����2A��\f������iH¶���?&0�#T�����A�!����kt�<S������$bY��$�%�Q�DK���&���-8�U�Χ��}�L/v&�	��0oN�W��~MN&Nl�*�2��*q	"hEj���e�tFj�[2t�iޮ�SF�km�Ae�����VN2�N��*��7�W&�M���caࣥ�<K�!Re��.�b�����\
t
��ܟ�璶�E} Vx�B}a���*�wBb"���8B�]�ҋ�$6F�^� ξea�2�{6̑����R�~�s_��
�vEJy�.�eXX:�,�g�O�Jz�niǾ+�	�ڇ�$��+j��T��ysK&V�U3 W:~�c@I*&��nR��\��,��)����[D�J�{m��%̌�$W�E���:��d/�Ko)2O϶P�G���HGA/{P\wOo��#1Y�=ѝFU�"�-tk�o-w�,|:P!Z߱iP�T���bR�	1� ]�4���A����@��aN�s�Z�Wa��fL�s�R�+f����t��3TR �j�t"�W.7LX�~�#i�����&A,M�xdfY�]<�%�e�rR\��1�XzJ��g���+�c�O�7K��C��{���>	*�fG<A���-�jJ��bk��5�����{d(��Igs�v�V�POA����˔㺮����vk��T�<�U���Uϊ���Qgw��g�T	�u'^x���$��m�A���$U��YМ�#銭p�Y �$-{^ȸ�3�ŝ!��J뷶�>�H������eգ_l�O�S��]�8�,��ݞ��F�k����$,��>���]��z̜
��&�%H���[c��r���o�!��z���P�]���"E�4�@#�	�/.�pm��a터�K�A���5�%Q�Ve� 8d��C
	���ȃ�x�R8E���X��׈��C@�H��H������wCY�� ~Y��Ȉխ���4͖��y-�`�]�ʖN���jƺ�'�&F�L��Ec孔�c~����
�JFw!�QV{�ƨs���:ϗ��4WYޮ��)�u}�&�vET3��z)!u����Ur��[�0�7f^z��y�r*kX�����)�r0�!{�(����T+��$H
3�����gW�כ���21��Y9�{�_��[�%�����JF#\����>���_&�Y@54�M-����`�[@	���o���^������L�Hmx�8��k<��5��g)��:�	S[�͟���$��s�Ұ�G��K`<�"�����G���`�p
y��c�f�Օ"u�;���cP[�F�d%�k��pg��� w���BZ�Y�c13�*\K���#�	A��ݦ�M�bӍPJx��»	�Z�:�R��r8Ns]]��Ի�}��
�B�>l�R�����v.Y�&8��V���,6���~�ך[u=,+js��y�����ۗ�7���N����R�E���Sa��K[�����+[3��R]�0Ý���������m�^��j��Ю����%7�{���0
��EQ۠��o1�4��[T�1�٭i���@v9�`�`M��+��VuI8dɛ=��}3���[����ų�-���}5b�q��#C�\k£�Aż�<���WƂ��<Q:�Ғ8S���/ʂ����#�4�3�+��&�D>Z#��s�R���z�}ـz��v'��0Z�pL>P���x�Q�o�z�[X�w��S+(����m��}E�?/��Y���^�և�=fKY��!�ff�J�%��V��)�������vQ�7{+�uط�J�}�T�����C(��,s�=��B�j����#�������R��j1�Co"J�Z���x�>��I�Š�eF���~R�)�U�'i-���Ŗ���SB;�7t��(�x:m���b����.�rY�4��~�7�^���-[? ���B����7�.RddT�d�Ѳ�Eʹ��E�x�����i�7��q�3ɐ���S�2�;]:��kSǔ�$���g\+{6-)_�S���!*����t?͞��Q��=,���F �b0���������YR��R��X�.@v��Ԟ����ko3�_&��s�P�⏠�E^&�g�fk�Aɚ��=�η=oj�b~b*3�E�ޏ���[���Iˢ�� �?���`n���+���N������L"����{=X*�n&H�ۡp�� �8���#� �$yjbx�f(�pPFHr�P�\e�<VhɊ��i:~�j�nw�A���h#4��$x��U���4W���_���I��hs6�oc��]�4-�[v����Ik�$��z�Y����o_��*�O�
��&�Z�ʊۛ쑲��@�MJ�O�7�ϟ��L������Y��?�Mp�q����V-}�԰����iw;�.�~֮_����-�~�{�UE����(=x���p�Ȏ�����i�*��v/@�#�H[3�3��"�,�'��y�������	�����+;� �~��6��̹Q��nN�L�Py�nZ� �#&��Q&��ot"���8K[\j~fE�7!S:*��uB{�`��;���7��y���q���A��?'��FJ�3��(O�)�iP��}��[��l��Λy�,�:�n��}y����{��S�')H[������ ���S�����.���SlF���r��H�S3R�;�%��,�Zԧ\�f[ϜR��ʤ�Lp��)]@J��=��=�G�첡�.��F�7N��=�&����z��Q*K�Z�.�i��%˗�]�Mɖڡ#����g|�E�T'�3 T���[%�_��͏5ڵ�N��x	J]�(A�_���o��3�Ձ��li׎���-p$R⒝+��b��l����%�����s�IJ��t�����;?��6�lx�̷�_�|2�V�Ι���>�&��uuJ�������Kc��׳��}�� �^�L=c�?%���&�e����7݌�D����O.�0�|������.�����A�����!Yګ�@,G���-|Kz&��|o�� q�E����n�z�YR�Q{h�U2�τ�:~��~ȠQe����h?� "��̏���.�Asqo��!�t���5�T(���.�!��X�Jx�ve˘V�
�й��%E������~�nTjAu4u3�<%��.�7���e��<�'��n�E��J�-�(��t��i��C ��������bK�EUQ#�{k��^.��%���U��?��, �q5��:��P%�#�0ܹO_rj����},���a�����E1cr��5ͫ�>b�#���� �_W����d��&T��5���k�
"���A�[಄����:���uh�E�R�Q$4��i�S����V�ҡ�HJ��f4v�tdy�4JG�<b�W
��N���X�Wj}Mb!އtAE�;�bM�R-	����W�t��m�0�n��"�~���t��P�kJ��X��N�F���2_B�lņ4a�����吒���Ô�B��Dw�H�8��(5K
��X��%A����q��D��'0�G�
 ��h�1�˿��6b�'���,l�t?�M"��}a*w��u�#`u�HB��|�ÿ��$\�W����Y�s5B��0v���A��Fp��_�6c�Z'i�qo�D���b�;�\1L��Nr%�X�k����6����P���{aE��y2�]��k/;��1�C� �lЀ�u"�<�@�q�cjW^1;`���VyF � ��j����;�fa��Q�!�ZC=��46 
�y�S�İgHˁ&��%o%�gl9���ʉ��Bu��R'���Ic�M�����x~l`�v(Ko���O���CW�F���$���a]��Y�=Le0}�0n�Ј*'2"�;^3�k�j�TIdf��(����2OW�#7�Rl>�˛�F��*IO����j��A#�lGr�N�6�;�`&ʇ����T�mD?=�F-/P�S�9�m�{����]^=.<�~�絧�繞tF��¼�A�K�]�9�d '�{F�w`�ftpE��x���L���M?���U�1�`P�s�q`��
"b�i�S{����r�����+د/�M	�8�q��T��/��x�_�
�O
NDRoD��::���i�L��" �&�F̡�q/Y���Gh��["�I��^�IK�H��#��G�J�R͈5+;�YͫlOw�5�����	U�E����D�����,��S��iă�k(���RMc���8��WE���X����b���u�V�?3ؓ�pW@��z6.�S1�΢8X���G-��q�_�Z��=�6���a;e֖���j��������޲I3�zdp'�i��� ��֐����n�\7z�� �)�LtN3�8K7P��2��h�h̀J��l�� _9�D�BvA����/PE �������J �q0�+���=Z*ZD��7J�`����z����˧��+�(�� 8UHו�Y���P�W��{�W�Q��{gȾ��%Ud\�Ė���m?���>"o'��F�&�����+�ֶ�R�Q�m 5�E���e�%zd�eD�]\I�5�K� �������RP�&�5����� 9��H�rUޥ�l�R}O�"�K�FB����4�\��L�.�N��r�V�ʜ�B�j��E��s�N�r�#�z�U�5���D��lb��z��5�D���3(���}y$����-h�1�()\&W	if��H[�&a��=���G��DR�J	�hn�ޏ%iD&F(����kM��h5��)"���(	r�M�`�N'e��2��8�u��N�O��(��E�` yY����3.ؾ�j�y�煝Pcn�y�@�\�i��.���5NL$5�AxY�u�d8����♛=��9 brQ�M蕗_s~���(I4,E�X3����*��C�ˊ��ʕ^D�0V8{� )�P�*�WK��/g�����|D�~��D��W���
ԩ�X}���3����b�EzZ���Jh�Y��zːN#������{
F�� �H���1�"HM}wl���q?XU/��o��̟ �@ϛ����Bv	_2����#�L^?��O�)���~#�� �o�$ ��-������:���!�,�DF/��J�������ja�{RrS�.J=J���;�9�@�ծYi�8	���>6��dO�m��?��a���~����#ab����֯��Ws1]Ș��n����\��gp�������/�)Ћ���4�Ҭa<H͇jI�kc��AKJ*W:"�!���x+^��&�Q*E���a�	��"a�;'��)jxj��}��]|��,�� x��;�9���9�})షܐ�5㾈��\���X?�'B	�g���O�;?��(-���c�co�2��:Dh��جEkzq�t�{�%��VK���B>� �-����:rw�\�ˀ��r��`#��Sǥ�M�lt}���IW�����(K����?������=L�����
%Yi���>m1c�l��ǅ��>���%t*�JAh�L�����X���
��\VU�O���H���rcd�4^�
{��$l}v4]-I����(���1Z<e�j���c��C�@O�c���c�l�qJ��H��О*�����u������4�Y��W���	��yi��W�<�mwy+�.,B~�l_V�Z�#R?E�E�k���D>���T�!=��G9�p��+�A��a�LM4�vڽ E�e3M4�l�+cM��h,d�1��[���Ɯӹ�m���E9����G:x�|��)�3�Or�Y�v?�@#8q>W6�H���H���ɤ�/���P��ZTY�|A�q�{���N����C��Ȫ��pe���7K&	x�w�S��`�41=D�5ۧVj�f��� ��)�f���B+G�j�g�z�gYV�LJ�9^��z����Mdj�C��I��52�ޏ|�D��f��s֭�觝�"8�^����M�XU��|C��Qr�(P����p'����y�'������c�uu�"1�WM0�J�RĠS���(�����:���x?O	��B���z�j�8L�Z�0.��hf6Ts���7H�Y��s5^�N�.��.m�\9�3�tԸ���n���4R�!��I��*�ew�h�84Q~� ��JW�jl��	�N$J���Fq`@��׶�n0Y�3�B<+�Pd �X;�[+�j�0E"|>q����`�v�Yr}l��	1���q&�o�-�r����&iy���W���`�_����-���)j4�gĥ4���7�ճ6A9b%�x#��/T6��Eg{ST������WgMc��t�ޏs9(*r~>tg�v�5�BW���t��a��� j{hP��|0���0�E-e���g������'Ǔ�R�ŉH�,Z7U���q�)]���<�$�����<U�M����b�(��4{����'�A7���C
�q0�M�� �����&��7P�Bu�|�2�N�T�݆�!�M�m���4�G�f7���5��&Z�������e�K�O��p4�w[�"�������[�$x���+�6T�
�i����)9>�SN� �7ӵ���i#q��q���Q�É��ʞ���`V/!�;�H�$?�A�T���BU�9����+��7Hգ4��RW]!I,��o�(z����6`�{�!�����%D��k$㓥:�C��Q������MS��x����5�rQ�?[�sA���ļk����8ZߔT�fظ�H���x�Lڼ�^����~+<�2\p�]NM������&%�����%q(iM�R��;e�M/]UQP(�.�f��I��J��R����7;���*�߉�Ƀ/�G�%}�'+�^��k_�D�,�'��ȬB(��SYZ��<���K�]���U���y�{B�%��9�Qf���R!��De�y���j���Y^!Ų�%ZmlL�.4o��L J���9}G	�"2�^l�YU�W
ǣ�e�z�48b�:Ѐ|s֝W<��D,�~��m�Yv�qJ|$����	�YkG�ݖʆ��:�0�$�a�='(���%Pmo�s����������k�v8KDz����lyxp�ǰ���I��х���Lכ��P��g==����(C�AB >�#�vQ�[a������}-�2)��;8ElޞQ/��wұ>u�^����=�"����_xaE�	�t�O��Y����w�̈́�qMW���~N�C�&��'ƙ��|�W��w-�{��1��xx����)�#�$r��0Lh�A�O8��Y2�ZRW��͠_,Ʒ��LUz=a,�c8fO逘Y~�j��f�^�F  e`mUIW˚$=���Y��]'V�C�����h_�u.��q	4S"�ocKz����xX���uj=���9�����aMԍYDF�NyS��7D[% �#�?&*�=p��))�	LV_ap�к��<.d�<��yʧ���Hx#��c>�.��3C-�������w,��z�>.xSy�+�0���s�/��JpXLd�~�$6�]i����Hb<�i��N���I }ģɉ�6X�M/Z����>������G�i�����=�zh�҅4#����բu+H��a*̐�ց�⼈�JU<zyK��2X�q�oĿ�>�9W8��{	�&�;�ӐrE��y�&఑���Ķ���o�����XR��%O�>>�w�tcq>�)�cpK!�c9sg���0����2+����2�x��O��R��:33�o�y��p�*7}��s�Լ�h�b.��s��<@:���w����Y�eg�LR��B� <p�R6#;Ǝ�q4����4��Yk6���h[����B��7���uL���i���?���'�,�xl ��A��0�k$�GI �OP�)�	չb^|v>U�  br����_Wĺ�݇��7$��u�SRk�,j{����k�X����[ف�'wz��Z�LZ�S��k��s�;0O�Ob��7�}EM89��s��z�K���e&��t�Be{&��I>���"h��EXj�:��`No�S��X̏r�ꍂG�Ji��j���������o\Z���Վu�V#j8mo]���6ݬ�K1�a��x) �Б��?��GR���XD��ȗ��-����7�aj�"`�����k"G�D���>�����ey0��.��^u-BlF��4��~��h�]�y�A��24����]{�-����
��O�"�3���z��9+�o�����o%ܤe�)η��Ll�P�@y7q��`�:J��0�e�S��bn�75�Tw��/�:�bHh���r�u1G�dN�p>>Q-�G[�c�L*��eJ���p&C�:&�'Нy�ь�0E�PJ�h�!�H�O)n���U�Ч�ޱ��56[�f5�7�#��y���X�����N������Z˙t"�`�[,�:�XD���X#�s�m�Th|D%q�l[l�I���j�N�(-@xi�~�P��6�RG�n�
A'�uqӅ#N��C����1�E�.�f�����r��<�7@џ�[	k�z��e���c:	�6cu��uH0R�^�W���]G��& �+�m���O�u[�������]�=
�X5�s1��lfhq/�iҒvi�� ɔt��C5(k�W�=σ%t&}������t��pjTQ�=r�٪��녙�,�@o����^�T2�����9�/��{CϨA�zS&m��Ҹ~�N�����z���Ѩ�y�4��b���+a+pn���C}90$}^���<`?�:���.(�.�[7�%�<��N�) ����H�:��=�|�Z��R>F���%@���p�*���V��,���/���|���=W-۲�'D���76���A�$1���/�z�7@%���Z���|��8yhP��q*���Wx�ղ���fG��� ���R��Wη(u�/��:��HE(j[�z��!����z+�x��	�*�V"��@�`�ZHTe��լݥz�ji �nO�Y�#�Q
�ZG�+I�/qu^z�,������g�U��*��5�4-h�L��vO�rƝ�vK���o|�N�4�&�/% �pr�C{6��l%���3���|#$Йv�%a;����F�(`�1Gi.�{m�P_�^��������R�T�A�a�����g}�M�z�J(�Ӡ�q��ϥ�9n[��ƴ���4�����ܒP)�z"-��j*EL�?�S�wvJ{���Ϲ\��P��?R�/S���lg�	a�Bin'C�߁<�&B�ܱ�n]H��r�ӝ+�,+!��e)���8"bʟ����������h��8s�̈���K�5�����_I'v�F����L@
Rd
�cM4R?�|S{�7���Wkt��6+�U{����N H��T��(�
�@�C���^y������؟AG�/.Z��+# �T�o���B,G1��)�,�+[��p7�j��l�g�YEn��(\.M��m����8Rj�m�����)@��@�!�@���^[������t/]�և��AB2��P��Rb�ןlWV����_@�O �-��^�e� O�)XIv��)m�9LfM��et^h<�j�7S��@���M�ceE�{���$��T����Ȩt@Bϗ��i��L)�Gm�V[���Mk�5�qy:>%B���U�Xlc)���i~�R��+1��Ϣ��5�ŹhK�X�MSA������U?9�ḥ�ˑD0U2{S���h7]r��<-�"�SSCF����ߊ�H�7R�P�)����S���;��e�k����Xi[t~�
�V�tFs�r��ӳ���!�Wn:��%�|х���9��_������$�ۭϐ�m��\Œ0�T ٽ��%%;������B�HaY���4,C���H�6�87<����:=aV�aԎ�$el{�a��x��?�+	�[�(����a����J>���B*Ӑ��	�(��"y��
��f{3|�gA<��T�N9:\������I"6�qc�A��JK��B�9��M�wƚ�����j�H�$����s��2���~�`9�Mv�ԭ�7���.����&�����3~��BrɎ6S��g���vdd!r��z,O��R��_� �n�qB�">0����b�\-���
%����1,��I����J� �7^`���L�.��P�x���E�ЌV�y��$D+H�����~�7�[;��.�OhQN%Z�7�gFO�`Fݲd᠁O�%��S�1���3eޮ�:�b w��o+�LZM������MV�S� 8D>�|O���ڬ��ȑf�yՂ~�;��p�)Ө�z������X���@л����mSF��S��,��A�s�^����4gӻ�Mv��4�����7�#���71Kz%}��<�.;m��&y�%���U���\��H�$b���w�?E C���Ӯ;�8Q���w(�����C��)E
)�aVc3��sX
M3�|�x%P��� v���,7S�� ꨚ�����-�c�&�زx+\�H%E��Q�d0��L��'p��6�����"mn�җ0��A��k����ܯ��+�=�!�^����(�e�r/�߄��f���:�
�R=Qr~��L���H�?���%��FL���#�Q}<J�y�M�r���+?)ܔ���39�Pϲ��-K��|�E��flY�'sF��_�P6jc�y�VmD��ۼޤ.����T�23��5�鿤O_m{�$Ew��xh��`�3P%�k}Tˎ�:t�@��B�V&�\,c�`�����Xu �+7K˕3�bLa�?�M_ܺ�\a��K;VEL���|���Q�+Zpz�m��-��@��������o���UU;�N&>
I�����9�l�j�i�`��r��%���x��	��,��i�!`�1��w�<���fEQ��u/gP:
�Ņ� �jJ�U�mj������Gy>l��a�]¤�����L�Q�Q����cem��&N����N~��a� �����_�|)�f1s������>���+���R�"���
�˛�a���}�.�1���CJ̬vfD]d��v�%�(�n���X���	��)vT��k��~Kٌ7b�9N�߂SZ9���F{��9�E��5$*�˅vɹ��dU��4���k��}��'@���ҭ�	�vqfo>166.�#�R�g�����_���������r����u��+t5TX��/t�t�f��4%v��H��V��f]� ��V{�hT�|����ݪ���Sب����zY�G�[9 8�T)���i��1������*1����!=�O ú8��'F����eY1R���jh�-	6lB9�p7�TB�fK�G���c�{���4D���� �`��},]`~��>f�6����ےl��>��%���#W�Rn�[ =j��Q�D����1g���F5+�i�{��F�˘S� 61��<>zV��1�g��2/�
����n��ĄQ>*��O��>j�|8H?��z�k��ai�:u�[�G�j(�����T�]K)[�hܖ���d� ����9I[]���:�"��*�W|�{h&�9�<����*�>�
��!��9Mx5#��C@��ԋ�K A4�J������YN�DI��+������E�i7������S�^9�Ұ��$��f���&o��_���r~|,�\�_ 80�
�<�����|���H���z]s����-i���`�]m��)a\ڵU�5C�h�純+.�_�/�P�f����0��S�Uy�h������a	2g�ÿl��3˒];��BR��*��y��qEC�ߒ�V���a)��O���	$ԭq���\C�SI!�h�%.f��$,�������2���y���g�P�D�����}�k��`�js��p��3e7�0��2���/[�HWDv�w��z�Ï�ɟ���uVIL�W��K(LP����i��b�J�N}��+������t��r�B���ˍ���
FP�1����m�-�b��Z�s�=!���uК%�Z=,��!���	� � �z�̩B���;����Y(�f�j���Y�f��%��c�9��\�v�Bސ��r��T��p;�l�2qQF/9��e�+L�!N�� �; �9��2�a4�>x&`�#d���Ċ��{�aO��lr�����2d;��&����'ݓTg����\0Km��^�PQ�IXߴ�q�����?���Y
�D�i6Z&8����e�.�l*�0��@0��Mc�
H+����l|�������x�-�����
�����f�`m_���K_�ކ</c�k
6v�9_d6!K�-l	n��G��t��b�[��o5Kllu̥�n�O(��w��w^&�6!(����%R2�T.��uHN�K�I���;2,\=�|A��E,h3�!p�Bt��ʹls�$�[O��F:��X`{�����əo����aT`�,��,��q(�x��)����*t��[���U���"}�Jy�H����N�#~�1�R	ĉm�u����5c�\�fH���rߧ��3�����S=��ec���U�8]=p	 W�8��S�/"�
��p�|�6u���nPJ�7�0�}Dc�9�6�h?����W�,A�aR:	�OL���'������3��1u��T֘n��!g��U�������S�#���y�w�� �p��$!��R�a�@���w��(�TG��y�9�b��їtbn�J&����7[ˬ�Zf�����p(*\&8q|���Y;|�[Ζ5��I -���W^˖�L4:����
�������yV9Zn`1��Z��Xo-�q�jU��c�S�T� �a�!�Fs�;,�6��v�M��E��h��bH����f���U	cŠO@�r���3,��I�mC��1��4�ѳ�liBj����#ף`��� ���Lo���ri]�XQz�$|b���ǘ��#�N5c$�_G���Po�E����6��dw��
>�i\����g�m��ې.ũO~�^�x�%J³f<� 6����
:�G�9����ZH}�� 1�Ӌ�2JW��Pc����v�(��/��V��;���k��#�6�����SȲ�X*�D�㊜���)�ء�q����j��+*zo��Y�EգD����r�]��W$|7��������;���y[.�r��dw0�jI�� `͞\��nM�O�Q�����/�DU8��iS�z^�t�zA7����U�ju-����g��x�7u�L��9�e���̇�~��C�&�Ͱ#F�Y�S����1�@�ץ���D@f ��w��ϴFj(ͳ���������[�����½���a8���08���r���\���"�@������.!9�n�B5ۚ������D�KO�������]�N���ͨ��[Ɲ�$3����b;R?�Fr0���:�Y�7�%e+o��7k	y���|u�G���S�I�v��/:VuM�8K|��as��B�>L����|u��3.'F,R�뱛��-pƵ��f�>�B���O�T��=�g����7d[�/�B��Q�:bo&C��y�!0"�U�Pyˡ��^��P�*��~�֝VF���M�#�z��>ΒOg~f���I0�3m+�ˉPC&�:<��wb���#xI,��V��P�8FZɳ��~*��A�����0������s��tu�ȇG��:����Ӂ�>��UG-���U���gK	"���K��{�[��f����KSd*��� ��*X���ђ݁�BC�r���D�I�f~�م�#�-�0�E���BiqdL ��G;���zw�A�9Gnq{|� z"����Ve��Ά,�}<c��ǂT�R�j�읈;�.�Lu�@��|�?�%��[d�	� �?������z���?��mc��
��gS�c��낍ɽݗpz/>�39����Ty��t�7v\�Q�RF��z@��ܯ�Qe���w�Q���-�*���<d�f�C ϔl���*\x$!�.N-���n���
�F�w/�J/���X�r�;N��Fw����!��m��`؂��S2=w
�j�'���E7��^�F���1�C�Ԓ[����䝿+�Bi!w�_���SY�f��#��T{�vs
#�<pztCs��ǁ��(4Q��gn�}��\�qU��8�~I]�{S#��7ؠ�A"�r�,IrJ��M��oZ�gq�@$��G��(_�F~X*E"Fi�&�U���E�,�������z��>���2b��À".wh�X;Ǌ�����������͙j��i�)��yxL���H0f�E���5���!\�!?|"�cKZRFÁ���.�M+����������?��\�!�^	��T�Qo����_ڳpQ=�ǷT�]`^4؄�K;��뱔��ڃ�q��vs��>�4�;�hp���Yx=d���봎���{�����j�GV���I�X ���e�0�}8�L�<��ˈP���iI��Ð%�Hb�o�<s-�=�^'����弆�>������
N�Ռ��5�A�8�����s�k7~"Έq�0��f_6��Q�)�IG��s��,z��]��C+�k?0(�M3$����:��iu������J�@�C;�EMd�	�AP#sd5��]�̆�/��X*8���u��->����gτ�̱K;b�b ��ү��e�]�	x��3+�B͈�U���ҝD�_e;��:C!�y'MFA4�ԥn�^�m��
��-�E���H�	/�x��M���5W�htpʷ���-�u��389������ʭB)�$,KrR�]�5ˁ��܋M9J凪���ӆ�5Q��Ʈ�Z���'�1�aD�P���~��J���Av?xT���N�PE����0`Qӭ�k*�X�wr��Иs��'��[�ꫝ�᠊�1�QhxS,�4�v@�m
q����X�j�� �H��WɅ'�C���[���V�Ibd"�n��m���dcx���sH���+�r�O���cɰ�B��9Ɠ�J�q/OڠG
$S �7�7�xf�x��v]J;���I��s˭�0@ѣ%�h��s��h�M�J�(�`啶a����e�iϴ�9�H�����+��=��Pb����bE�$wZ���n`S{e���x�µ���T)�-E_�u��
�n�J�V�9��28��`-�X�A䴵����ߋ ���2��)a�^oQUJ��s	;(�d���E���v<�AT^ĭ����/=R�̗�PT�)�<:S�r���a��@�������OFF$a�NA�o�/&Se9��� ����߁wU����M�����/�������PҞ��r#�Vڅ�B���3�S>��q�#��Q�89�)�Ì:-�c9@��3#���ҥVuD�H�������g�Y�v�2�NZ΄�{����K�0� ՙCx�r᎗#����M:F��.���N�Q�c���U�W���SpN��=�F��x|H�o>h#$�ym����Y����l11�ꠅ�CG3!A"����
��*��	~�[�cw\�H,�G�˷��[��+��̶A�"aZ����=�x�U��#��Y!ۺ�\�K_h���1W�������[%|Y{������ց���#�dY��@���f��x�4�>��y,&]Z�X%V�3ۖa>�н �1o|5�w���D�O+���X]������#%�Q;��n_��A��p��3p�0���f� [��0�(ճghe
�L퇯���$�t�}����vFX7���Y�Rя�jtj�k�V��� ����U�Ԁ���l�"�~���E��^bJrm���Pml��ۑ
bK9���Ry3Y��,�P"����9��I�e��@|�������F�[ݖR!q�u�~7q��'�!Avn�[}��i�s�UU��β��܍"H��F� �6/�X�Q(��w� �Lt�*�LU�B_�X�hR�3��g�W�xN3s�NWBu>G���ތ��ͫh~���*�ݥ�-׼�û��Y�EY�c'� ��`OX�kc�1���$�p;�!��<�V����$c ��e�j���{1<#XF�d�BF�ą�gyj�)!CiRLY�$J��:KD�1R/ k����Ў��R�Փ����	G#��No[�������kf�*<��a��ݾW��a���)N���Æ���E�/N�x�	C��sk���k����hr0�c�re���TѵaJ�I��/��)4*u���k���mw����E˛�D�8�g�~�k�A��i=&��J��TJRtU(�����o�~��b�y-��0�r*�c�3��d���Z�Y�+��Ob>��x:��]�:�[�٧)�+)���ҫ+�8��5f�YU�v�j�'�e0�'R���.��ƓG�QꠁZ �h�<���:Ԥ�I�J���/��I�V�rG�J��O-X۲$�K�{;��
2y��r.�>R��v�C\r؉נ1�;����?��V�Ɋ�]` ط�.�vh�����0<�����{A-MG y;��Rc=F�-8W�?�T	s.���M`c������o��n���GGj#�
A��Uƌ2�Vx�|�h�0���5F���f�ה,AbIN�4CE�}�v��`�Vk��B�`K�������i!�>�FĔ�I��j��S�a{��ѬT5�H�(�Q�EU^gD꽌{�^ȁ�i����Dc%,U�V�B�7�MmV��;r����070
W�-���	�<�?d��r���£��M�l7T��H��@
W�~��<\�ب�5��	�+�6D����c���w;M�4����O��)zZ���~M��w\��</Й9B�u#!YjU�lE?а݆�~6>3��~Ϋ�5�����i+��x��[y�$ɥ�yKQ/���ua�Ff)'ﶇ��v�+s��U�-��:]l�ȮDGn +x5*�	6��h��/-\OpdiS��S���>_��;`o�� �B����������8 �=��Jt�6t4��mMF�/q���:����8|���%i�r� ¼9���?�w�c�;�,E��f"��}v]E�$�J��mOCS�����q�9�ֶZ�4�O?z�\���N������=NZ�k ���{���i�)��}�(i�����K]�q
��\�0Z��;b�_����дUH'8�e��(���r��MjY2t�hP��~���Yg��	�huxg������S�D>�vu|�}4�V�a�U�թ8�	�ߔ�u�o��c�f{�q��&�9Y��2�~/!�Ke��Lp�gw���X}��X�3|��2�|�q�
{�lڒ�蟐��6�������>��� ��_[R� ŷ��9��۟�;)|�J4U�36S��BS�n���.}zh��#k6����j���ށ��9���?Cg���#���
bU �*K6'�GT�k��aE�_���~�� (��k��F��6cr�|X?7nl�+�Tn�hF�I�@� ��c���@��5�<za �Ȋ��G�Ǩ�Բ��3�j����E�6�tr���f�Q����ԌN�=��R.rPn���k9迪,N�n��j������K��:`)Ѫ����o�O>�2�����b�ŋG�^���zj���8�G���[n`,{HE�r��1U:׿ĳ�ʶ"�6���]��f�����)�V�x���8��`�n1ˏُ��*�8j��|Ԇ�y���`��98fK?*yr�pM�^����N �8-��G���d��|^��%|X5�^߃�e@�c��"���a�x�p?@��W_�CE�׫cccx�ϲ �y�)���l���2�L8M��a��_|V�Tc����̖q���Km5f~,_�V�w�?Uql�u�U�5_y�*e��c=�Fz�7��e�}�ϔ΀|?��{��g���]����ۃ��Z;�9V�X���N������\��+����,�w_v�<V?r�����4����AZ2�}�N�./�X=�����+	���S֍�m��V�[��p�18��=���BS���z ]�'nC�k�pX���]mc�6�ͼ��K�e�5+ŭ��j��Ǡ�K>p����K���#ϤS-�d۹��^i=��$�^�[ 5|_}�	�����a/��}�g�?�"���>fu���V� �u�;@�-���C�4r��uT�:8����ѣ��<Ӿ}���Iڄ�&*m�5��*	f �h��6�-P?�½ �52/ᢻÿˆ����8��~Z��#~�L�����η�y� :��65y�1�'9���r������\�����Ҝ7�q��n��{W ��\����� �+���:#Y��s�/>�k);�!C&��`��s��,jmq�W�3��PS�	Ǳ�ͪk����3SOd#߉�s&��:�:�!�F!��x(4E�����M��f�P�f��i�=��BE�����
ZLM�Ay�(�k�I���}C4���y�(�c��zx"�T�e�؉!���'i��?���p���HRA@��l��C�h��/;��#��U<`�C+�J9~_��a�^��Ж��7���n#Ƨ>wYЌoVn�
�De8��'1Th;<.ޙX���4_������	r�8�o�"����~�l�X�RI���k�{��G���"�PQ�E(�'C�E��.�Ϩ UN�:���jr����ȘL�K5��+����,�s�"s��N�`�1�x�x����Q����tV8殃}�;8�V���	4H�}VP�v��d��\C�z1�����r��m�\y{�Y3�+Kw���?�3���̫��U���~+SUf�#j������U���V]�iN&�����8YumTx���i�_=�+���#n�B�x��4{�%N(|��8	p�&	R����X��U�W�:ڧT
�Q�l%PF)BA�#�S�eB9��4%;f��0���`;0�}�*?���E�H��hy���y�l�d��5����&�q=z��qI5%j�h�]^�kl[�0���+<m��GW,��n����R���^~_�lqzK�0M����X�
���.$����T��-&�&�䐋��>R0W��$}��.t��vLA�Р�+k˰��d2���v�Y�^ ��?Z����ët�"}�����5 �a�?���_Л��+���+mͦp�[l�	�Dh﵆�غ�0�etP��������FYȟ�Da~�F���Z�{eM(�&�j��t�呸���`����F^���=��Z����@:�=(g��z���M�ܢ�Ky-�ɫ(��».�<mq�JD�����v1�v�6��~�h�I�M\�Q[����0�B?�������k|3f�o�a����ظR����g&z���"7^���"�,�<*B[�e{��)ka�䌫 E�-\<0(}�x����XƤ���(�)O�# 8��.<&	� ��S���є6��N��#7��2�������W}������L@���ː����,��+�e�6����1+z����[TMs��e	�B�~IP<v���<T,�+�x���0�E� �h�>�kA{1-2Z��l�r0�K�#�#��a2G�5�A�7A����1���pěS����ue��
�I4�*��U����6#�O�m�P�d�挛�a��Ø$-��1 �������<!���7���
W�L8*�|�9Wi���TxB_8�ԝ_���q��tC )��Q����t���S�|���3��R��q�<FD�S�"3J�#�Ka�ψ�X/';�##��R�D���s�6,J���Ǥ�5��Gd\��H��l>�z�]A�0��+��L��-��-��M��^mdp�G�7v@vg-�i�r��SK����ZZ�6���B�h-��v����v�,L
l���#)R8����!�3">�����C�������p�%�+k8DE�]0�Y��y�.M�Հ Z-V��e ��E�z
�v"���<z���{1ݤ��/w<,��p�|�royrLĐq���,���[�=��3�L,�SV&
pUK�
(#07v��=�Mw�!�@�i#�xTW�o��&,#]���v��3���M����9 
�#�ϱ��i�:pc�ǂ�$csBUU�)G��l�{�����֑*�B�^ܨ��<\Ģ��9�1��{.5��X���i�ހ��׵h"IjkAm�Ȁ���N-òˤb��e9095���{�-�Y�M��vc�aZ�3Z�1M�a.O��j4Tc�DH&�'.ų��|f�4��zLa�d��L�e+@��S�(��BCw�YN׸�YyS�	�&���b��j׆�hD�P0|�﹤�I��<e3K_�$cC�X��9����8�[��!C40�VE0WD�|�7�a����H �#`等gNt �£n�H!y��,��b<t�T��(���*���y���!�Mj)	I�F���	G-���D��}(��#�GD�t,a���J�}X��OW����r"���Ƥ����Oh�
[u�IZ{�)x�C��ך����t�P������N�Y�o+��D"��*$�0H���6���&�T��|>ma�$M���*�O-�sT�fe֚zC�W?�d���B֥��A��L��e�3~1f��Z�o�US]��xH�.�(kgK����g������hQ�7���m�u<zw[6��	'U�H�/����_���D���o��-�u�s��{�&��$�#b@vf�¸p�p�u&�"�5i���X�K�1������r��{�.¥����R���{�0F:�e�Pz�OTn[-����8Q��r��g<�htR�?A;[�������$�4�&T�[��qT`UQ`'�W��X��YL$����7w����B�ā.&�"�;#�����
x���S��/
���s#�gZ���z;Lpk���a*Z���=���eV�<$�}E��;_%�,�yCU�G���ZiU�W���pZ�	��`ba���A��*��5�����e����N�َ��\�}�¤�>�	�$t�;���мIhٔ�(���{A�2!|��T�q[ƛ��l����u>~�#�h7p��sQ����DJP��D>�+�E!��8�?Z���$�˞8�ӝ&Dp��i�(�L�c���Z�g(�<�V_�1�i��;�3����c6S/R�&ƹ<A�rfM ��ݕ��H灂�������ζ��$n������ڙ_�dNC��؋��*:'f�;���@[��~�ܠ�y��'{w��O�����1!)����}����s�h@���^b�$��S�|�;��1 1*�SF#�0�7����X��̀M҆f �aVE�_�4����#v�㎥Z�&�J�O���q�dh3�97SD-���$/S�m{Pdu�nv�b)�K)�����Vw�����I��g N�
��������vt.��}ϴ�{8�!�g�6D�����Q��+���wн�%BU7�mT�ڢ֯�W��g�/�X1ݡF����a7~9�9=(ѺТqF/^���c���4�E�5����1}�4�h:n�����8{��~Ho��=9�<VD�qGנꝹbߗ�d��W���"� 2dJS��W��d�ƹ�@̭F�7ѱiЗ:�"9�s�ha$�Lܦ0j~�'j!��!l��79D�~'�"�4w�-@�����pB�YZ�Fm�����%�����--�j�ߤ{�+ޡL�F��hq��Qf^��=�7P�Q!fv�Yq�àZ��ҬY� r�EG��{#��K���U|v��֙��g[e�]��z7ݾ%�7��0�[��ꂍ������~#̯��]�����6S��t����s�����f�t�Jخn.V�����>��x�<�����0���kf$�BJ��k�%д�����>I){��w0�5�!�l1�`W�L�Z�oY�-=�!�	ӳ�Z�S7W��-T	��[1�I�x%T%`��()Jj|"��~�{���;,�0<l�Q�m��o��#�����<e�M�LK���}�aGb�ԯ �2P�O��|�z��Yp:w����"ƈ�5Jy�S������r�����'���3�Xj��#fl�C�!��bvv�LFZ�/���� �O[+c�ѭ�u	�8z����{���D������/�d���-|�4P ȉG��E��E0D��^��Yϖn�����Ιۭ������I�l_\��pX��X\!Tv�2�������I���G�Ic�s�tE�ѷ�Qx�vD���, ��Rb�<i�����M*N����g1����� i�>1�(�gΞd�H4M$l���������J�Nǐ�Vzt�|
Ԉ	��eU˃�"���SG��l�&�A�fQL
��;}˨ ��+B�����>�P���Wۭ�^��+-Ü-&gk}EkuV����d���2�!l���I�}��dȶD�����	+]#;R���M���mm<����z����|�J���|�׻��{n��^K���G)��W傼͹cA��ҍ#�RA��w�SgJ��~N�*��,bl�����a^�&����%P�Ё����|\����x��;�z}Ve#��t�h�0BQ���"z=ټ>��<�_,��C>O{�%k����X�ѥra���gK�U	��{���#�yr�TR�S!�.���vҘd�"U��A��V���v^x,ߐS�Ҍ�45�Ҧ��%[�' ��@r9�����2���J�=S1Nj��:����Δ٘����� �5[|��`�C�ףek���"�ᩘEp�F����_�0@�X �	P�c��*M2�����mt�P߬G��N�|.';Je7)�H#kiʜ
�~5�|�_�̀�<K�\��Xnl�F0<�3vI����
w��օp�s��Q�Q�Kl��^Q�T�E8=�-;�
�KP�rho��:"�D����$"��w#`&$CF��6>���F\d����N*���^x�e�������w�9F[�E�յd#b�ʺ�VM���}.�����(��������k84��ʱ{y��U�!��Z�d�}|�+QБ�2m?<����B]᝕���^�@�%���"�v~���4�A�!���^y��:$[���T�F��Ҁ�If�L�������X���2r�o}C�^�1g����
7��/�)�5��g%P�ۢ��[U����Ⱦ�(�~V���'D�YHM����*s�����jk�Ƹ�s��L�w�svgf�ڧa{��;�+~���,���g�/��5�Жz�6��9D�s����5qDً����ֶ �?�g/��>f�K:༠��������xi5�8�f&m��0nSO���@t�뀹�˒��?�,>�k�_`޶�T@u�W�L�n�zn���SS���g'�#*v��vOU��}����	�un ����^�� �����=GI�(5xXV�R(�w455��o�(��VNV�t��������[4_=sּ]$�\�`�~�?�ᨱ�1D.K@c��?�G8�<��8ܠb1T��������c;�tI�h/�����xz3?0�4��S�&}w�)�v�����+	��L�CM�U�����p��1$j�|a:��\j��&+g�4�ՙ3�y�*���*��呱z���J��$�ݢ2����nT���ʼ�~ ]&�	�)�<%��AX�k7f
������K'ļ*�������ّb��ѵ��3B{���H=�l��	�e\���z3
��\���	�m�Wz�lfd-S�(L������	�:�XO�	��%��3a�Oプ2ޗ��\h!�a�2T�F��	��!/X�r������<�����0NJ� EJ�����ճ����N���]%,@0��!��#�	'�_%֓�apD�G�/:������:�J^�!s:�=%9Wz0zx���=���]e��3:,170:5и���7��=�X�m�����^I�gM��1�=,1�K𩨋�b� �_YJpr���^��A9�}�iT7���RԒ⺇��1g�˞�L/�>�Tm��늣3
�
�����a�W�8��𲻿����UEL��k��D���M��$����p)k��C��$3���	|�Ӣ�O�S�m�����Mr	�ҬR�_Y�O4�[�r)r�!���*P��n{����r>����O�ܡK:�Q{4Q2G���V�E�a菇)M�
�L������� V����mr~��eu�28�;`5�Z�E�� ��)v��V`��ؓ�n����e���e��r�c5y?\Ű?�c��|������L��� 7���4���l7�8���ٵ]�k3T�6��Ӧ��������PVE[COŪ8W���̕x��Z�1��|�?nT#�����$ݏB��3�M�����}�������ڹ��콆�~H4�>�m!0�K�/pȴ��]){�7s��1�i�:V� �G��*���%����t	���zq�lv�����VUt)�Q�M�2g˾��]��:UO�;��[�ڏ����\�ov9�Xd�$����I
i�9�ȭ���
���-4�
M�z�!r�U�, hЅ7dZ���	 ��9`�q1��}�+哧s�x�d����I��6�A�έS�HN>��5X�OW�?8�%^'�'�X��H���#�y���0�
cɒ^��ƅ?AR��z��E�Xq�W�aA+���I	r3�#�x���5��$A�Ӎ'��}I^ʸ�S����QA=kE�]��-�3�S��P��qJ4+�Qt���*쟯�6����=��0�3E���<��o����es�7�s�E}��aT�Eγ&��,�[�2��cY��j8���OCd�F��WU�|��{�&�(����]�p�A����6�mWoP���[||��[�����6�a�%��Հ.��B�s$��cRI:pq�l6�(��w��P[[��f)�PSNP�)�J�z�~;���/�zTC#�������U"G�L6A���-d�֞V�6@|�qN8r5�QQ��	Z@�:��Jm��� fk���S�/����YXJ7�T��jgt�A6���[Ս[���A�Ϳ@��>h�l��!k��y渘�!�~���s��3����;��y�E{I�9�����֏��7�҃bI�[\A�߱ t4*��Iֻ�y[���!�֨n�K�p��'��GM��#C:�/�w@��W�6�E�P����&���H7�.�s�n�̂)�;����T���6��,/��FY�N�*�f[^�u���4El��c���h�tb���D��E���\}5.�H����z%�gf�݁� �V%v��ه,{��	m/�8�N�6��ꀤ�>Wqi�<��~O�&��@V��m{�"9�5�^慴���n���@�8�ԢH$�.7c��k߰��b�տ>x�T]e֩r�c�"v�e�M�7�z���T�V��!7���@��h=Aa�I�į�%����xZ��_���S�T�~����M��4���/QK�G=��:��y��MvL�����d�����R��O���/^�X�S���KA (�R�NJ|��ʍht��O3���\I�j��@^��ꅘ�A�o�e�>���Z�Q�//ć/�/�Oڮ����*;$8�1��t�t�=]"Y��<Ѭ״��ͬ�gD�4��U�u92��5�����P�G3n$ȢM����h����;�<R�hQ�O˪����-_�%�T��K�������
���M|L*�ʫ��;K�`�Ǡ�	S�^�8XY���8&�)o�^N��Y��na׉��a�'{y���谠���N�/�K{��N�Z���
W��!��d@�v�>�WB�+�\�#�y�]�����ǙX�����^�@��;A�8�Z:qұb����4v���}����t��m}-�Kh�n��x��q���Ej�ַ	j�ux�����{%@�;��.��y��S|
M=��PW	���$dȐ���ϫV�v���m�zR
`�"i0[G�[;�ȕ����Y�rXr��Y�g�/3e���T��>��4 �������RPe���[�J�,��ᓦ���ϯ��!�/����Ȳ��:5�N�|#�	"�]��Ai�)[l=3�� �p��mX*�+e�@f@5�p���������Ç-բf�^H��(����U�oE}@�I��2h��z/�QN���e�<H0��,Xwl%�2�o�ԇ�"�ȫ*���U�Z4��0�����&F� &�iZz�\*����b�~|@hv��~�O��? d-F�gyz� �q��}1�ﭪ��E�6EgTTV���9��c{���k`*�b����[�IzL�Ғ���Y|��<�Ʀ�-�Z��!�3�;�$d�Q|o�t
���,�K@>�]��N%˭�@�5M]򘼅��3z,@Q��Ɋ4�T:6�EH.4=��x���㧳2��
�BB�{_+|�\�Lۭ]�'ͬ�k�\y�n�`����$h��'5jR�IX��Q|cp0�&����f͝��f���̓��]����-����\t��3Q�-]��_�V���e=�h
`������ӟ�l����d��� i)���0��B�-P�:��`/<� ���m���]�8-��S	��(��eD�v�F:bJc*��/�!���s#F�p��uvsZ�&����N4���o�~�����dq��<���V��h�}��,��{S�E��&ֵO0�<s�4��னe�"l��?RoS��1����=1_���'�y��(գ�"k8�Hyz[v&���4%�O~/���\�9��5��!���=�A���F�l
�b��f�
��Ĝ���S��Wt�Nҏ͉�h��������'����|u�"I5��jY�'��$��v�O���崒'�Ro�>�r,�6w}bXu.1�t��8?.����9^�ֲV吤����_,��Q���R+Sbn��_k� 切�����~?q�qQ��0�r���n���KB�Ĩq�u>�DD]W���va5���mEs.��zae^�0���Q���Ncm�%ҋ6�nT��p��v �]A�!`�,e�{�FҪ��""�q��%ǰX�^����m���!v�U��-��!%�_<�0��bJ/#{ɞce�X����G��{��}�;7���Nt0�w.}����=H�Lĭ�� 2q�[\���s�c��hs�=�wHQ;������q��Ade�������	?aMC����:AJ�jFNHA&4W�8��<�*�js	6�	y�ֲ8��A���ɊS+b�VK3��uP%=!��{�^���h����I����)u~1�<��q*H�xBsVa�z����E�W�r���[�h�py�гt�"p;��� �3�����q55�Lݒn��N��7v4l�D"�ٸ|���X�&)L�T��w��ɳ= �@�Ƃ�Ӓy�7����P�����(6��"o�H�W�M/����_�4�!�Q%��!�8]�Oǉ�}H�-PD�[�ֻ{�4���Eu��UA�2%�,^?é�`�1�,�2�a)ث��夕�{&gb��U�l>�~�X\w�Pw� :��G�x}���J�"�+��b��S��]�$X���*(���߸��\�Y��xUh:�� C5a�qUk�8��B�ղ��J�K/K7�w���Q�P�����U����e�m?�W �q�B�I���(]�QW/l�;�ۅ��oAlz��(���Zpu]�$$�U��=�A�Ռ:�`��B��j
�5C#��V��*��]�J�n�l�MY��9�ic���	�Y���my�� ���ϭ:��ծ�"�M����>��F��ٷ<���o���*]������D��/?-fO̮��w	��,�)y���cxFw�\ef �2병�c�����nu�?�N����MIX�w�?���*���da�O�n�f7w
Űm�S� ����\�{#�@�C�.ͤxz��m�%6�|ns����c�J�~�]��Ͼvmf�(��Y�Q��7���_����˂:������(9',�7�ȧ������v�D��4�H�÷�Rx:�r���Ӻc���j�F�����q�r,hPR�_�E3ˢ�ǐ����&c'��s�-^��+n�IQK � �|���ΰ�e1v	�[�U��+_�zܚwwH3�`
�9͞-�[�E�Ȏ1��b�Ӧ������%��jZ��!��i�qj3�h�����V�3A�jxd���R����T�N�������~�}�)1-Uv��da0v�݇��{�*h�e&�X�}��I<�<�	w�.�� �.�$�y�Q`��eȝ�%12���36�å�+��5����Lث�u���������%m�O�e�\k���b�!R��F�4L˿�~ν� ]M��u�Ż���>V������,���l�[�f�Έ��GA�J�J�s���z|vb\�����m(��? p�%m*~R�C�s���<�k����yXgn˔�>��j�_�g���[F�|p��@siG,fUR'iv�{@����fy�O<v�:�/�/�{r���o��3: �ݴ���G������m:%j�g�qv*{��+�qUMت%Aؽ�q�n�/��e�8%���4�L�)�v>�֢�w�����0�C��;�>�H�
�C�ӻ��𘔚���BD�����S�,��B�ja������Z�_�n�U��Բ���0�ˌ��9�0��@��S�0zx�a�V�Ԑ�S�^'
��"ο>�g� N�w�+�T8x��
���0a��!�za�^~�&���Vq�]2�r���҆B��,�:[��H��r͟��RK�
A��
�E���Cx���~VK��D�E��fx��D՟�XÝ\R���H�����4WE�|�t�Õ�4��+��Q��xZ1-C�"m�%:y0��ͮ:���{���ل��B�P�VC#�K�l���; _tƲ�J�y�$�\�F���u!1�"7���X_t��-�u�9���GI.����#��,F��zӞ{�#�<^
�̓Ƀ��(�]mۚ�A�`������_�o�E��Ẽ#Y ޺�O������W5�?�<癕�Oh\�s���M`H~�����(�����My�pX�����ʀ,ޕ�	u�I҈�P��+�e�����.R�:�xwy�+g��A'��)�O X������ac8=&��*�:�x:�XGQ��IN������4��4�ԡ�w2\�!#f�����^\���eN2K�ֺ#����F�^Pw2��v�eJ��',���0l�y����~��ۡu��^�&D�Hy�vK�6�Q�r���!��l�/��j�o�X"��$��(�ͱ�m䎹��cм����)�(��� �B���E�7����k�-���hxǌe��ݛV04q��$��v<�a�A�+�Z�4;꒲g[��ɱg*7�~o[<���iU�&>ׁS�<�rS��)�oo���<nXP`\U�߱��G.L���v����u��\��
��<�\uʿQ�<��:ajq\��,��
�E�?</Hʒ.~�e��o���]�>�(�ռ�uU������0��h���(�L�:��72W˲��֟k5�?�gs��A�*=�Z������e�=�����FO&td��&ȅ\D�2G�JGD��@g�E�`.�0+�U2��$�F���qiu�4��'�E���|c
|���Ka�;0Jg:2�w�)tp����?f�KK�v�h����e����^��`�FaL�=%X���/�u����0�PЛ^I��e���Z�K�f�ό+�\}>=�i2u}K2����~��f<!���|��C�c|� ���D��]�׉\HM��!b]��.�4�11�[*����O�ej��$��X!�Q�.��(��7����xb5;�(����W�#�b��>y�5��L��'�`>i��ς:"�� 0u��_s��������)�����q0��%a�g����W��S�Yc����gfG�� ᧵,"�b�����i�6~M�VS��'sM�V\����F���z[z��)���t�����JjW�1n���܇5�Gv
�ͯ�A�O"0����U��C=�Si��½�$���p5��b�a��n�6(ZRkXwHq]�fP�D�#�g��R���2�����&]Wv���a��,���)ك�I5;n7��@k ԇ���51�� =�鄼��f�84@_��?ͯU~"{�k\ea
��z�}�!���i��:�(ky
�~$,b��NO����T������2ia��f�u��逦�2(���͞Ǖ��F�LߒWf�����$��3����M[�N��9�!�����NX�uE՛e���1(�M�G��G�q����q}M�t��c�ZV��הO�E�����z�Lܰ�8sH[��;?��J	�Z�"~�p����cҦL�A���ж,��C_��u�9.�Q(9�C�n�o'g�-�:�����d)�V����'DI�E��t9�*�@�[ ���f�.���0a�o�	d���LR�0c7�&II��R�!��f��nX1�@3�HԹ�Jܱ�����/y�y
��j�)=��̷l:�@c�U"�"*9G��;��4Fa�]�0gVݓ�(�h�/w3��;[�g��d�ro�J	B�o�I��ґx�9R��0^�.�̖�e�hm��ȑ�X!��1�=q��3��-W�q'� �,���7�NB-�?�����$� y�'γ�<�m/�+��a���N��02頒������q��+V�6���C �w�%�'�Iǈa%a�\Ȭ��]�N-I	'Aٯx��"lFv�����Yй��,���Sk�nP��v�|o ���lf������aTN�q)x�6E ׹x�u �u��:�K�ն_f�9��|�#Wp+���#]v᝹��1�#���M�ʸ$�Ԁ4�b��"�:�pb�),�zPԖ����$=�'�+ZD��r�H3�9r�~���r_�Am����8�;�� A����vcn)����r��@�1vyHl�w�B�;Z�{�I7�U���xK������l4�Q0�[i�Vr�[e�5��a���9"�ϵ�����!eG�=�W�'�B_���^#58�'+kY�h����>��H���q����^�hOg�j��3��E�a�h>� ����Z9�f��������7���/�� ^�1jF�X��o�`�g��0��c�YOL%��q�f�Y����&���I˧��&+:���sld��6��;J�ݗ^W��^�䘎�L:v��� �Z���p[
\����03
��������`<`�V�Ĝ��j酈�ibX���_<Ԟ��Ǹ���}O;����8m�"G��Z���D� ;͛�(�&���-T���-���e,P�'!�x���QV|WW�vE��KA�`�?�W����T��/�N,��I���
7�>�*��NiJE}�L���S$���
c���UI)}��Јf+%� �8P*�f�,�gz��K��/VX�r��nO(z�K�4`�1�a�ؠF�.���U�é�j���[�+8��9[�0_՞��IDxa�anI!���0+��N��P��!����ɸS7{���`���ƹm}"��æ���t�.�vܲ��H�xБO�A��j�}��L���<��+E=��J/%w�iߙ�9�b7/+�qۻs-��5KIO�h��4���5���#���Р�����}SG��ၞ�Z�7gQ��i����}jO�6�sU�b�p�b>���̊��G`�W7����U�ڵ����R���'�.�A�1~�e�'����ps�,7���D�^��2�O�ťL�VT]�/�8�ب'{j4ΐL�wf^���Л�Ho�qJFY~���o�p�2��i���:qS[���L-�{N3j0Y�n�
�P�BD���Xǡ���;�u6@�#�]ĩ'9BkJ	�u9d�B�n�X��+aP ���}����]��c�;�!������`��qU�HV��{�?�]^��>[$��D#�uJ��n��=�w�f廴V	%''��Jbq���IB`���YezB�cU�7Ͱ�y�S�m���	�L�	�&)/N ��Gj�[��o=e4sC��8!M�.B��ǐ\�S��k�j�N�o�&��R�t�0���E���%�xI��"� �����a�Gfs����Zb�ߖ���Qu{"�P����3
k����ކδ��"���ň����sV�2T�Y^��0!��z=L2�I"uY�i}��ж���%&۽
*������=Y�t�+�c7�yG�ؚ"���7$8���!ozZ �#���ݚ�3����0RQDM�I0P�v��A2�	��,V�GVk�Vcs����OP�k݉(��Q��k������Qt&�{����[��v�x��t�@m����`3���#�Ӛ-*��"K��	n�d�n�F�Y�d����j}y�`�x}˞�n~&VcG���x�x�	��~��P9N�[�0�Uu�&N�_q��St]p��� ��P��0<߹�O��ƃ�hd�O����εb#Bmjx!fNi�pu*��E\�#H�n_��yK/��?����m�"�t%)	�R@��ObȊ� '\i���ȴ�B/*�t�^�c7�!���&O�����Zq~�%�P� /��j�J�#5���L����(���(�Bh4V��d�)�Ѕ��N���=v��4Ѫ<+�B�u��T��7H�!�����X�v����l`ߊA�����z)ݒ�e%���I����3��*3�,P��K�V��������J	erod�Z���\F��۳�b�ns�b���8�߽���� ��#.�Ʌ���&Zz�˓C���,�p�.cgU�2�Q�9����J���g�ł"g�WvZҴv�i�Q��	���T{o%�
ő��o�M,�y֫~{�AD��X�C�׵$���ƔZ*�.��X�c����_�p"�綒P���(���??RAↇ�s��I:4Z�zL���'��x����߶�	����+�~
|��.�J](O�U|;Gb�q��^D
�֖ao��.�]��Q�8D�ʹ�2���Qv!����a75�ќS���
��#�n+���i@hjb�Fc��V�g!.�
�@Ҿ`bu\����Պ	��� �3��$d���\m)��/����l&wԫ�X�2(��jB*�H��G�T�#��C�h��
R�r��4�}���A�K��-)�X�+�^�I"���x���Ӧ<��Zz:��%��1��l�ԩB���.�,N:�+q�V}��;LI��j-?!�M�?�,\�
����	���<ji>����)�-�[>JD��U���'aƆ �7�|9%���3mv��Li2���n >�ɨ�-�]�lr/�3?ƢI�@���;9�4h��s��Nd$�D��s8v�;�������ꕮ1�15����&�PD9�3�����f0��#���7�	�Z������[H��^r�"q3�iuj���_����ó�ŏG��7�L�j��vF�uy����Y��_m7[�
�lP��>��Jȕ�-�?z��S
S���^��1i����g�Q�Ѡ�|�{�9<��-��ز�m��Vhw�\�g�r*����t.�2��߱�k�����f n��̒$����3�h�+�+x͓n$��]����lIO%[B�{�;%\VC�tzuF�L�I�l�� �H�`���d�g�}�ڿ++?�KSZ?e�S�<^)���̻��g���Օx������7���ܡU(H�'b���1P9�+c/��YZ1@�9�4}�9K�O�>��Ƹ��M)ڨk�{�ƏD���ۢ^B.0�,մ��7'�?�jn�IT����f��I��kZ�CJ!
#P��uf�gΠࠜgq���3cO!��9���P�߶1���E���%��vo3���08��{C�$���J+���m��ā�$9��N��B?ʭN�B.M�gX�,`��g��9[M��\?�gh�Wx>n���wuCLS�@~v��g�p��ڝ���ۊ����x@���(s�h�[΅j֨�Ś�S��G�J���vTх����J�9�2@[!����E�?7���yc:ieU�\~�Q�µ�f[)��y���}�)K���V+�.�����]`���\�?�C
�N��& *����&�8[��8��g3ձ�P��~��W^gwUYt�����ͮ>�%�v2 X\����i��݈7�9^�6�����u�	GTs�Û&l5s�ӴvNrU8I�
)_�m�ڸ�p	t�-��X�,kO�`�0��Z:JE}`�h�IE���v��E���9lzE��
8|�U>�ϴ���#U#T���
ڱ0��Z>��H���q�2�&H,Jl��aѵ�I�R�U�ƍ���)Nc%V֫�9e��w�k�N�_�,��?
��?�|������5f�����k�X?|-�6��!� N��]Qѡr�Qp�~�d �ŷGUl5$�q����D?�j!�Րh\:K~�
^�/%�'�87b`�Ҧ��A
(�S�8�{lC���ř��ɞ�{ ����,�R����Ȭ�`�)������1h4�ء�ǡ�D�܈�a��8	#�S�:XO����a�BtQ����@r��9%�lŔ~������w��x��Ȑ�&L���˻��h�� �]3`V2`o3A� ��bI��~�ݣ���2�(P��&���S��@���(Y+8c!�����k���9l;f��	3z��J�?���aO�Yq4��T��.W�l�:@'�׷Z~���~^`��k���)����f���8]��_T����e��n�Ҳ�Щ���ȋ�\3-�I冤��x�Zc#c�����y2}���qzuy&�C� ��SA���J����Y� Q�6�d�wsȹxRs9u�=���S��la��utёy��5�b�ܻ,�r�!��Ժ���f���'�;g.�Q������	�߻��~t����<_0���;~ø�f�SWj<V~2A�u9Ձ�N.��1�7�CG$N+zd(�Q�)5���Lw��A��B<�/����	���&m�MA8�/�*N���aajY
Ǟ�]��Io���^��I�r����毇��7��3U>�6��˓&/n�Dux�_S?�?묶�(G��,�p}�ᅍ��m�:��<��q6�o�Ǣl4v>j�<�/4�6�a�93'�r6�br���>��ԅE���Hǧ�z�K�w����MwA�#ZL:e֑�v浢�s�K:`S!|�+D�Z>N��3��Z}F�,�ޡ�( ��K�z��6��ȶ6禋�D�L�'��T߈��Vi�N[Fu�����@��G��/�׌��5��M����� /�F�H"�7�ɪ=����'=�J���i���UAc�����u �5����yG${Ļ��-����80
�Hko�"��a�������_�'Ϧ�ܑ�xCaUX��X3�$p�>�凞�H�?G��fk|xF����1P�:��	��?��k��w-R�/�W°�K����/���x)���"2���X[��o�	�64{)Ɓ��rQ'�a���QV��p3{���Y1�P�ǚGv'��3.i�ܵT��N���7A��0�]�r.�O��<Ԓ\�;��{eD�N����K��E
î��Q���i��D���P=����|�^��n|�f�UL|�������<n��_�P)O�ÅFj5�zsW|,���q�a%=X�o����x\1�O=��j����2ڄM`�(s�;�s�U�$A�GfE饾{?-i�zߓ�x�Y��䁺��]����� �$�"5[���Ϩ�3�''ϯ;�=:݄�	l���6J�O�#�l��,�6$�R�0\w|-Y�h�\�q�4�^W���y!~��7��1�q��LrO�*.�Ț����Q���3w��]�L�֠�j�k^��}�s��H-;��9���Q3���̥��i�Jƾ�ŧf�q�9�GF����P<(���-%{F|�Y�'k
?�kNSNӘV tħ�C')�{��En|��6g�����+}�AX=��K� W��sE���t3;;���;�EOdz*�1�=���D�^�ޜ:�NX�e��g
W�hq�si��P�.tV^�0�����?��C���?s�r�v��Oq�Gb��m�^�RE��$A��tʟDzt�}8`\2�1P�j��Y*w�ޜ�a�Í�`P��@!�gbs/WW�G}Bҟ�)!�oA?��v4�v�z���7�L���u[K�uIT�Ԧi?@��IvU�ŦJcFi��C����
b�/9��A{�֤U<�[_s���3Z}y�.�pK�t��*	΢"-v�>w#1�g�|]�ځ�ąNT9� -�ꌒ�z�h��^.)$���m$��d>��vK����GL��)C�y�:Y6n�F��VCxjز�0���Ϻ���>s��i�j7�033	8����!v�'�d�UF%�A"�$�9��,ď���$���"1����a���LoT� =/m��������؜�xD�{�HOX�K��n:�yZ���A��'�9��:��#�Μ��ŷ{{��W[T�9A�ڶ��LN<{R]Yy�
�k�t�b��V���^G��_�f�d�*s�\��I(��_Mhۇd���t����{�O��J=Ŋ�$8��.gS�X�h�����ε�<�f�\������rh��@gp��ۚJ�	9E���$ikJ7:�@K�Y�E����N�p�� i�R'3p�jc�v���~��{��4q�;�f1 C��d�թ5��Z�$��-'I8<_� ����6W;pV\?�,j�.ZY$b�v^M��M���^{����^��|v33+�\B�H,_�ߊFܑ���V��xI���(�h]�Ws��+�l��k�>�2�����?d>G�"!ahMk$�3P�z���"�+�ISg�r?:�O$�I��ВqJ���q�!8g�P�<���j���U�!�0�6T�yf�;C�R��Y~�{��wP䍨(&!p��n�e�u�Ų8Cz7c��$���,���i��lh�d<x���י5F�_�Z�d-Y�ٵ�w���c+�@�ˎ��bޙ]$�>˝��'z�B�ψO3�_\irj�ZrhUؖ�H|���)��V��~��L��l��i�ˑ��H/��^��F�Zm˄�l�~��AV�oǑU�o[�eu)��&kޣ:UOY\T���$��qnf[�ëS���h�U�\��a��wRV�VX���-��r���Wy���^�]ɦ����$NtM&M� 8��4���-�Y�(�~�80�n�	�<t�Pr�f�"Q��Y]xǴ=G�~.��@��F{X-�Co����Șc �!#���������~k;�������8:N�CZP|yJ-ԝ �Y?]N��u�V�D'��<���)���U�)�"�`�OJ�i��r&3;h.x	+?��Ƹ�%0�|}�}���Ix��_������n�&��[�-m���:A��@��\��h�L�bK�[^g�<mGՉ}'`�ӕ��He�	��tu�F�"����V`Z�����l��l2���-2����x��9l)~�B�����|��s���&��X�h���IՓm6�v+X���3+������/���dO�vj%���ܥ��:Ë�/��y�&��fg��J� �,{NN��w_Am�'����%�(~��"�����r���'1�>+g�R��^��S3S2Z�Zv`� ��'w�O�Z�ˤ������|�ޑ<T·P�i2����(g͑�[=;��^Ǳڈ:X��x)�;�CA�dGs���T�����؆�k�������Ӛ ��E-���T_q��LU�'����P������Q�zbQ����뽔RIi���Io�p�x�r�7�}I�3�kG���7�n��Ny^�K��JtP�jE$O���3%k�'!�e�� ��������W?ed����P\��%dF��������*a�
緿@'�.�a��l䁀�p'E�����x���ܯ�������Ϯ�@���6xE�_����h�R���	)���8�y,�0�1ñR}�@�-�@�%��,���io u�j�{P�c!ɋ�^��M#d�Ei(0�p�]y@��x�)��9�r��O+��L,3Vv]��ëj����r���;��$�|�1b�N�G���ß��!ғv�,k�i�W˅���g"G�3��Ef��ǈ)?��۾�89M����ƻ�%��"v�`n5;�+v>VX����O&������;B�/x&�ʋ^�����$����5x�*߲J�lD��f�łlR����'η.1c��z�g�(���wӊ���U�>���b/��V#j	p����lO���2��Ix� �X\��o���.�� ��}k膁�`,��l��M�e�0�%�3Cɒ��x�(8t�J �z���G�H�&�*5��Dݾ7#m?/OĂvf��ir|�)�,�l�G�؟�xI��0H�s�w�ݤܯ4��"[X�����G�d5�G>JJ_/�p���N�9w��R�B8ӂ|�2ۅ��\�(�v�*���@�Af��3�]�T�Љ Co�['��[��b�pf��m1����Ԅkj_
)��$��!9�YE�e @�J;M
�~1'�	4!D�ERi
�Ӛ^/} ��򍴋�0�)�n�� sE�s37wޱ��b[��[�{kڽ���}^�m���K����o���5M�k�,)c��l".؍2�z������\ķ�g�:�|-,�)-���p?�������&�[��c�q3~�}d�͙�:�� ��
��%�V�@�����m����9YC���tİ�=�u#�£O����<P ��/��P ��g����A⼮O�����Cm��eR��\�U��4����(]a�i���O������WE$yG��"�s(:��K�]̰��5!�#��H��F,p������	�2�!�$�,R�A��0ɢ�/�Ez@	�p��a!g4ە5����c�L��?k`D�ޑ��(a}�;S{U/��`�^%E�C+}��-�4���a�ire����x�����!�}�d ��d�����9��+w�.�Z�͏�8GH���xپ���G��V~YD"�'�Q�y=���s��2 (���������[�ڶ>z�G/c���]A�
�R�h�*Զ;^T��ut:�t�h0&r�~�kdTꦭ�f=_�D2�#f��&1Mw�0��s�xJfΔ���g�z��3��4�@!�Y�qz�$Ÿï�X8��&1U&�Q��V�0&݀���^�;��~:rF���\�������	�44�&����$�Ơڴ[�y�)��qasF���\#�I���,��N�s�e�5�cPg�.���ZW5D��]3z0$�fd�����b��1j��(�lY�4�?3�
�P�[��Y���	^���UK"���� ���51��I<�{��3�	t��JG!�m�������LaZ(/��������)k�%LPKȗ<^���_�4~���ï
�	���od��T�7�my�vTA:A��r�(ȝ���,�Ӓ�)	���ѯGĺ��j�<�C	z�3�G�%�n۲eQ4K����@>[�8�|R��;�����|2ٟ�(�E����+��;q�ag�F?��9�\M�э/C-�VZ :���G�Z="����{�GkF�ZY�x��2�$fK��J��98��FF2��n<S�}�ȋ�1��=<��++�U晴�&mt/j@�Ȝw���yμ2\ �C �]�}aq���-+)����f�=�}$$)�-��"�jA�S{�y���V|����ݲ}Q�r�n�SF��f�����~���U�|_P����0e[T��/W1�xT1���x�뎱9���o�JiR[v��vtp��K#
E��F�>�Z��ƾ�\��MYȽ)W�{��iYa2'4�� �b�.����١U�͛Hx�}��&��k��&"*��Rk��ݚ��q�%[����|������BQog[�X�5aB�F?�!f�`%{�Y��|��� �}ĺ�{�w.ܾb�W���Il���X-T���ΈR;�)�� Ȉr�B1x�c�m�t\v�| �7�U ��DX����A�QL����@;`�,��b�[� ��`i�1�)����V�`A�єz����t��v��;��%�D
m��|��xa�P��zq��4��k@J��e̊�&ܽ��\��$����FZ�N��	�l�j�Jp8>����e<#�N���MD�ƧR�Lm�#\���`�j#`��2����>�>�0��:o�WJ���6U�@�Z,KeǭzN��M ���靀k�.�Ɩ�����љ;+�v�1� �X�J��NS��ӓ�̛�1�y��L����t�L�"/��]����<��C��soJ_8`C�Z���X@R3��s'���˚x'�c#?���׹^��D�W�r�7�ر�pYx��?ͦ|U��_����~��`Ձ��sg��ZO�-��P�B�����bP 3St�8���s�-��{�}��ȮrߤruI ](�Y�dhw��r��OVWp��e�-�1�T�R#��`*v/�-���fc��Y��Q���/TC�O�V������#��ա%Ǐ� d�� �����=�ug��l:Sb��^�tT�W7��bh������ID�2dX$��Z/d�5��� a��ܼ���JJ�Ja��W��њ���jP{��,�DO�B��.
+��4���Эo2��T���4q�k����9�G��ET�Q��Ŵ%��SJm����Z��U� �5JŨ���K�� T}�:8dB����Eϭ�5 �z�E��Da�	DT���D��ӷ�\�R�Ͽ^<����X����|�-P��	/�&��t���P�Y4�9���/��EWq�|��OYY�� ��U�l�~�uw��:��oo�
'�x��Z�a���M�c�9l>[��Pn������&B�+:��~�9�}�I��̏A9B�Dyg�0j�:0�b}����������0�t��o*�pQv��ה	��u��{��2ʈjƪ��S��X�D�T�~����\�aT��Ak�~�0#]�� QW�ԱJ�g���޽�m	����f���	otgO J�E��l��/�Z2�r��l@6��?����f�R��%8�PW�.E�FUA�g_	S����9\��FL�h���Bܼ�a�h]Σ���P���o~�s��T.����I-����Q �;�)�d���r?�O�f�I��k_<� ����'i��e#�=0�N����B���������`#Th�*�;,���	��%�%�Y]�=���W�
����Qt�2q���8讕+}�>-7���>"I�~un�p�N���M����`�V�(ICu(6��!��1_�O>"á;F[��s�۰��M�G1�rk��>�5����-tш.�1(a��@q
��X�s�?���;v0�!�~*�=�a,}�b��ߴ�A�l��2��zM��gԞ�|�C�R���!�^ZX��`�/w�;7@8Vg/����qc~���j��U���W����[�� 3�B|�o���U}eD�Y���(����T{� �l�׼�̩�c�vb����U�U;�wp�MN�s�K쑕B�a���14A�Va�IE,(��K���+�-_R
�v��3�W�;�A�Χ!>JЕ$��@�@f������u��whH��"#P/Q�@�s��,���M�WaP���l;���K_��:v>2��;���U�-O�>�~u����]*"^�z2W�n�$�mUnL�ۤ��1�&��z�o�f<��œa���A9�8�χ�]�2
F�6���R���_?��_5/��1s����5#��@ܪR ����7��������,(�M
�F�.�� ���U%��H��`>SF�cHqùw���٭���bm����X�DrcFr{�"��o���h�R�јHy�D��軚�J,/��~Q;2Ҏ�9�6H�P�	��1t�>��_IzO&K]�^�6HPv��3Ā�.X��I���V����.����,%t�xE� �s��C��e����_�q�q�4R��+=��&�V.A��3/V	>Ð���AD!e�l.�O�����(��	
�]��~�P-�h�S�Z����R�V��(eކQ�X-�1�� ���LȨ�.>��7��>y��? �=�����L���?;�hy/#�y���< ��Ey�����X�U�'��4��+�[QX��=�bĆ̦���ۛ���^�����=}A��!z"�0U�. ��9|*;���e,Hvp�am"��j�w�;8бK�� �)���}�:� 6ZHB�9i&<��$���$���r �Q���Jݣ��,�E���<���{\���-�F#w������j�UP�����T�}L�Lh�Wz�2+�r�"�j}�o��|���Ad�Cs:� mvSAn¬����*�_�qӆ9�{L����<�������!)
]��@`S����fچ��:k��Z9[�s-�0
�[�W��XT��{+�z��+�?܂����r�K�Lv�����fL��:w�MA�(�dQ�*5z�C�/{J������������pF?�d�_�b|�}��~]l�"+F=��1).�XHKju�P�b>G���3�������	�"������v��@���>~�$���=�"Ěob�ƞ������D�$a�h[�鍵
���K�&U鐯"�_~�j$�'��vs��r��t��ۜ**n*-�#���m��gύ��F��c�Ж�fݢk%�6���4��s���L�����O��t�2�E_�����ЯI@dw�8�+@��;��A��$����na�*<�����H��z�˷�Q����D
�����9�s ��>^��H�]8�<�P��g�@2&��g�M�3`�2�9�eq*�*����b)56�B��J �'=�Wp�%?��R�?���rx��XK�\O��BO�	0����j&�w:�oL�����)m�|�!��:C�o���ס��GQ�?y�}����t���r�KLok��x�z������;�v\S��3�D�{ f$�������_<̐�̋���$��~�9z�����E%B��c�q�&aE�3�R���`C�(3����y������P���Y�ǮTG��#��?XW�Tn��5��]�Q�)��+��K�TbD������:�8zN<[5�s��gt�i�V�x�EX�ܣ�w��g</�k�pl��jrBA��m�i�e��T?���4\�"�]�ֳ�e�#�ǈ��h0RB� �6�N�P\���0���'�f��w��T �e'���P��"@1��-k���p�$��7�(�G��uyA"�s� 9ޕ�z�G�O���T2'n��|d�_�8v�P�S�.�y�p�g��$�<�%��w!ٳƭ�ϟ���5 h7�y_��¯M�r�P���X�Kf)H={W�C_>^�>HD��C\8��i[B@6[#*$W5�V�90�X $�+qT6�T�RD�LW!������l��9=��
�2�o}��掣2;smq���<�p�3G��Ǒ��ℿ�vA�q	j#ȇ�-�n{ӆ��t3.��Y�|������L�t�U��w��4�p�hkQ{O{�Y��T��^n��q�ё�jfA�]P�mI�(�)�P�B�����J7t&��h���EO�#W��]�!�:�W\<���Lk��bt:�[���3M���c��Pz6ד�����^���\LQ
B�������F-Dr� ��B��H�6�?�"��B�5��n<D,�R ���n��z�^��ŭ8?���\V��I�G��JC�`N���7?�KiX�Oٱrᘄ�{����œ��F��%*UP�#2'GY#��fMJ��C݅{\��nYr���^p�=7-^i�3�ޤZ��:�i^�jQ��n���\Su�ߊ-;����_x\%�y�C�B��4�n����7HI��``�.�&{��j������� H��"G���:w�!t���e��0d��Ү��?��b�l�P��dI��#�{a�@�o��y��<.�nP�����	��?M"gTL�"��4 �(e�5��%2��9`X^vG��/^r�H����Swzg�y`���*��%=(=v�h��\���_�l�>���'�=���!��bv����BR�֛��;�@�G���,����+�bҮ+3��:.33�o2�1�R �2��I�����-&���jMg�7k�%@���u)��:C��g��k���8R@u�e��^�m�DR,�l��ɸ�~6�I��G�D��qtuwD�4��?��3�໹�5�h�Dٙ�r��ֻK��螈���C�^gx�,�$z+D�~̡�"�NB9����崋�ʝ�D�m	�	��~K���('e�ԕ�:�C�/���jcn�r{Eʇ_^��AD��.�;�	j�����`��Ml�c����<�oi S@��@lG{�C)LN�L��ڿ��C� ����Z�F7*���=j���
 -�6x����I%ܟ���X� �JO�	�E�_����g۰n�ڴ߆��!���YJd�ƯŏH�Xv�x3M`iHC���c�L��������|W�RH�,41%�r�sS��l"c�h	9�Ԇ3�=dP�����[-ԑ��h&�$��Jc�&�Z>�.a��f��HL�����0��=X���������nbyJ��.�^�Ģ��G;ځ"�?؉��W�Z�Zn�-�t���s����tG�wN�{V�W���bOH��5�x��I�ˑ�6�6��QS7��N���~��&��8���d�V��7����:�f}��-muGY����˳|R_��f���� �T�SNo�${v�Uʍٿ��0!�;6CW��'�b/,�������UH�*�F�^��O�;Hn��fWE�"g�r|_HǑҹ����N� wJW^ze������}�(��bA-������&~��G����C9��|�UP�Z�<g�J<)��U��r/�T���0Bg�*��N�>�;�&e�F �X���ûj���GP<�$21������IC,��:zj�l:-ܠ��If��]��U����j2ؚ�K���ܚ~��X�Ň:��Pl06�h�u���d��\��콙���nH��Q�3�]���ޔ,i
�IZ�u(��r�(�ڣw-9n��r��j&%���0� l f��d��cm&X����@cԚ�Z%�$��o���FM2.�U!��+�����%����q�O�*v�sBl�ȜI�i��^0� �aLйl`wy�� �9�xG��}��c�I�3c��p/-�E�u�J� �8}~ANKiٔR!�H� 1���#e~EIa��ܓ�Rs�4��m�`Iu��]�{tg@mg��U��i�Of���#�(L����/T������U9��fȈ�yTr�
Y�bc L��$	1l-!0�i���W��X�ڔX��W��Mh���L*���|��NSiuo�a�|F=�����/vO���(�pߜ�<]|{�SYrCj	��/&���	\ɳʝ�Z�9�.+Hm�<�4R�]r�Cp]U"?~2k0��U ��]^��l�͙�D�\�a/�iz�e�1 7A���+�Jι,ϳw�}�u��ʐ���oO�ʫ��o��ɨ��^h�7�SfJ�v�me'\Z���7��E\�ʐ��8O�%���8�s�$Ua�W���.�{��/���l���D]{2 c�ʥ����S�I�uFM���39Ȟ)�a�1��f<�-CL���S�A:�Kvw�{�~�Ҡ�h"�f�R-��ebrG�鬟n�}]�"���%�C�&c�F=T%�
˖W��4�ʐiTv�j�U���14|�ʇ�/E���{L�?���ιq��k"$���O��п���ƈ9qXڱ��9�X>�V�Z��#���e7C#�Dk��4����-�m�i%��g7��"kR;f�@�,��g��\u 8���5����RZ	��ך�T�u�vm-m�a�S�sƐ�>R��U�_���Cս�#��C�����iB
�'K�o���1$r����<D����G{N������Ь(�&$��"�e.[�*�����!E�R���-el-�p
-3*·C�/u�G0I��ޑ�n��Ԇ.� U/�_*OLz���?�S��eE�|k��˭��"Q~��VO�iI����VAt-˞�T���#�j�V�ږb>W�)ý>��E���C�޴��qM���30���;t���Βܾţ�9��e���&�u�
�ɿÄ��z�]Lk9��<�Y Yji�nCZ��
��p���_�T�ZJ�X.���*�J^�uW�<9ѡZ��ǲ	w.Y�~��%�*���bZ�D8�#�C��7���;��4�Kҟ��Hv�f�E�_�n�T�{u@��3�pa���$zR�$�c\�d�=\�qc�UAA�q~�&�N�����\e�����r�6�=�5NLx�FZx§� ��ϘiIm���<5V#r:�qJ�;=A�(���!�Ohv@�)��9��ѩ�^#p1)�H��+g�̳[�I�;���L�,��	��H����g$
/�{y�_��w�ȱ���?����9)RsL^�S���kh��_����|�;ٚ�MwS�Qg_��1H�$c������cxr�ģ@�HvX��p��;�\f ������X��\g]�*�5	���I���Y��~�Q6qHFN O������$�D*,C��/����϶8U,�)A�G~�add��q��JL�6L-��� �n�&2�ه�������tf�.������Kv>���>�*�g�v����_�N[fۑ�D}����ܭ}����2`fw�N����S[��)�I*D�uF.�pX���=J��ۑ�c����
�f�'�RD>$�ɲ9�w����_�1��� 7�����;���s~�Z���`L\_��bj���#1o�<�ȧ�p2�!%���54"S;�EZ۳Z�U��Q�_�k��!g�.X)��i0Q��� ���"K�	&4�S����e2�wu�̘k�puxA�|Z[��jyN�i*B0S$;|��w^	O�;��ch�1�k�\=��?����O��"���=��W�� y��Xw�N9�ђ���T�`�_W�W�q�B����G�\�^�r���?2���^����y*��8�q���RA1_�ټ޳�N������4�d�!��Cl�]Y�&�!�w�Q�
U�)�e�R vX���u)�@����|�iG��.w �N�Vܑ3A���֐G��lZ�SӜ�O�`�u��vX�8�̕G�����yo��=8 ��6�IU[��IRL��ƒ�s��gˀ#���F���_����w��L�@"����"B�S��c	��Z�t�m�Kء�\	tk�*Юh�n�d��4/O��z���<�O�W�����[�is�_-HY�N�C=��q�,	 /���\����-k����!\����mV�_����^�b�xE#��zp�2cͨ�Eؑp�j�pL�%Ӄ�|�X����F�6��`
i����o��&yO�_�5��/��qh#Gf\�B�"&���
+O��+y�v��B�l����@��=P4QE_0�E�K7��߃ȉΑ}�ɵS��ɵj.So�95�t�rp  �87�@�IM��|�b�aT�K7&�ۊ�eA�VB�J��Ʀe�ic�<�6m3��o�Eߊ��
�i+�
��a4{���-?�N���E����ff�w'Q�R'��UT��
HSg��?Dq9%%�����
_}UG��6�㈴9+��F���,$OlCw�UD�(#�F��Ie[˫P�m��#+��( l�����#���7�J��ɻ5�% ��g�x��2K+ZH�iq�&�3��u��6|���Ob�=��7%`���۱�^������t�E��"�r��yB.(�O��9�s)C�5�Z��[X3��� ��Ge�~ N��2�)1���c�mČ	�c(��_ͤ�KO���R���U��w�BQ�"�:�hܢ�"�%q��&���Ӕq�ʦ��)�R}�UX��Kp���5 �*qU����V�B�vd�4)�	4��A\��'������O�O���CҾ�} �~f����̡V���P���+�s`����
��U��9E�4M����]2�E3���vem�q�m��
 �{�5#����m�rJ�fW�s�oiu�wA������:1��*6A�L�Iτ�a5�������@�~�����/@|�6�\C��`��=�(����$�a�IG� ��	;a�_$��V	��[����:<�G�����!�c���
�	[���]�ҫ:�s��MQ"�5�������&;���7�/��kw��ZB���3_z?^|�\26��59{�>�5�MT�u��B��s��Փ��+��Nm��|�g����/&g�4۸�K-��mR�3���-#�?�Ǧ?��.�8��ݲ((�9Pr.��Y��5k�\�4.�U ��i�՟Z6��e���
u���IJ��>�xz%��+�ZRX���DK��Ⳟ���!DM�NLN�����_kC#?>T�E�j�����r����e�����#��'��d�Vo��l���Ԫ:���ug˶qWO�o�B@9�'�N&����]0���*��c}Y��CG��e>p��[����*�Ciey��G����G��u$��4ـ�]�@���Wy��|����қS޺iD3��Q\3[/d�k�2�6	���f{�m���;a��R'5���@���<���5���M�	Զ�'N�l6ʢL%��	���Gq�(w��Vi��X�)@	��վ��m$�}�п��Ǟ��ѥ*GL�Hv�"��-�,�@���E_v3�f�8MPs���_V�b�&[^�4/� �ĵ������<y�2�XGp�Mc\L��j08��A)�^2�.W���Al
@/N��������&S�7V�X��"�/��K�9)bXg��lDz���,ѱK�Q���L{���\��r�!�HR���M[;��j��K�(�Iċ���G�Y�i��3k���N�
�˪+��Q�~�¶7��xrp�]X���Z/���S�%����gM�5�KM{������	�Dݗ��*>(@����R��׉�!���5���t���>�q�p�����\hoS�M+"��}��(�tj��(��ESi��مU�;�,�Tx�%�t!��!@�Q�L$�[�j���f�2�̸E֑�����O��;��*UP � ��`O�Is��W'S.�*w�Ǯ�S�#�XT[� }�s�1�@�&��N�4���s�V�O���/�/�D�ZL�g��^>��&k�>�:��	1?&��3�U���(Ï���w��vwj��-�B�v�:�iZTp@�G�@*5'�;~Uh��%�Z�%��z�33Rd�r�O�b��8���%� ӟY��Py0Ĥ��R�Q����: v��į�1�@#G���9 ANz����Xae2�k�`��u�gI~� ���tX>��C���f`�y�f9z>�o�Ui0D�>�����&?�,��[�HC�C'!�qD����xX�(?0�Kt�}G�d��9C���%U�Ԥ�3#�@~ �����eO�b4��V`x�M ��Zhܔ^.�����Pʫ��	�ஈ*��[^�t�����tĶe�n9�n�q�5��Q�����B���0�s"T����%���kƚ�mZ�9��b�ț��j������3EW����Z�s�mh)ˌ�O��U�ݠ�n��D�m7=E�J�����x��L�Tp	�|��m�N���濜�,�����т(2;��d� 鞽S�� /�6�=��'�Q4+;	1�f1]Õ�L��)e	��Sá�`3��`B�|�Fo����Pb��������z8-�a��a`K��<�2P�m�\O+*��\�Go�!���н��'�ɥ�}[�Ÿ}@�4�bZ���u�q�{ ���Ŕ0�CO�{%K�����	�fH��[�[��wĖ�{��pQ��h�F��G�1i�C� ��{��Ku�ZH~B=K��ZW6�?<9ÿ&�%�]�o�	X��`n=N�5n�{���$@�+�ɤ	Gm��e�.Ԡ�����͢�u����X��1R�ؐ����^?]EmႧ�FΜ���9�����O�c�M��#0��D�< �w4����_`øz��f>nx�8�1�]��mmG<����	����f���(�N��7�zH.�@~x�x� =����d_���z`�tbן%�c/�z�ڗK3��y���n��U�:5���kηی���q�(�A��)��{��0�]1�ۨ(�F���Ԫb��\@y�P؆�M�/��L�z8oR	�#�����ғ�$L_(5M�VZ��Y<���;L�4{���a�1j���|�~8�ڽ�
#��K[1{@JY����l�����!��̨�$�f_��ҫ�	�'�W�Fj^n���SB��ߛ�	1�6�������G_�o�nL��Xen�Ħ�5��s ��վ��H}.H�·�
�O�Cx�e�'��r�3h�@a�6��`���J0LqR���}(�ڃOM�o%���>�h�4���_�DlF`���
���r�=)�lF�ԇ1�}��x��K�N;��S�&�<ntI>or[�s3�_�,&Yx����K�\�n#v�o7�h1�$�j�c��6�¡U i��1��m^A�ǵ�s��?O��Xc�-�$���(a�ք1@+��4[p���e��hڣ�'�B�u�c�}�D�ߦ�h1��C��%ΐ�L�x��f=����n������q���X&
k�=y'M:e��YA�lv{��z�	8oׁ\�
̉.�b�z���5�zB��#�3��L5�8e��:��@J<#+�pH�A���ޑ:ؑ�s5���Pow��zG�����O��A��c�]�  �6��ܨ_[,:���M�8x�����V�~�� ���TP�X��������x� �����!��F[�vc���O3Ћ�$ΟS�F)�F�4����B��c����4JW�h�����9zR��{�HՇ���������Pt���#T�>.bi�f�e�
/��qqPSX����7Q5���06B�%$$�L����r�e(3֮�p6�L��x�������i���l��
��ye��5�4ݗg�d+}�/��(}L�9��2���R��Q�j/ҽ(�1�d'��tQH+��N[�A
�] T�SA]s?Ҁ/�g!�w�A4í8�M2	a_�D�MZ�x��{�>!��J[��ڳ���j��˴.Md_9<�`g-�:��~��L� ��B�;+�����ǱZ�����⫦^X�ɌF�"�%{ K腚�v��A��(Z�K�ij�y�Mx<^.\�i��+l8eb�s��3s��[-vJa<I��c���#��]rF#�#���$��g!Ǯ��-S��63'X*�A�x���:&>Ԉѯ��S���Z���j��_�g�Y~,�r	E�� ���DI�ǀ�?e����h�q��1hT��B���4�����6��V�� �*���l�@�/���o�<�����5kg�����?f��9fUz����p��h�)2)Zg�?�\e �Z4p(�oc]�_�|����;&U�ɳ?C��?�s1�h�`B����tv]�G���v
�7����(�h�Iq�=F���DG���D��`�{e�+�D���~ m���%�3�ƾkT^�<���џ?���M(�4c�4\�/w�˲���� �g�5��͕Mݯ��K���C�e��,�H<�q����WZeQ+�ʦ���.vCI+ ���f7�ۿJ���0��a�o���劊S�hH��n�qOy����� 0��^�4�E�j����H�ܾ��n�)�ax,�2)���=�q��a#�zҹ�e[��+�#�w��+tEm@�5:+�a�流�ʓ4������,�W+��C�/�@�=��
�R�����:�!�1�ܶQ��;�����c�<�+x؛mR�A �h02n�3�_��,�ڇ���v��wȞ���L2<<���բ�(#��w�Xг�}���"�p�?�����p�zQ1��V�[�qG�.��m������S^�:���:�K1f��h���:��N�K.߀!�9S67�R���+��s��'�Ee�H�i}���k�V����y�}d̊ө������,a)�F.l�
�oh1]���,@�J�%Q�x�h9��+�'�hl��6ŋ참_*�6|�+��"�����1�yF-�(z�ƃ����Ǹ�ZwGj�^<Hw��s�<}��[d?pgڕTFO�vD�i0����X���J�;�M^qǣ�r��W�oL��Ni�Ց�K�:��? �(���&ϊ���^��:�6�2�7]�R���1�{�\�3��ܷ��N�4H%�*�1|�y�ծr�-w5<�Bt��Z0�ؔ��~٘9�uR3�Hl�w�����E���$XĦ-��fs��uUX?�r\�w�G�c8wJ�4K7��YϵIխ|k�zK�S}Naͧ䚛��BoSx�&p�t:�Z)n'Hn!�gD�|{ 1'q������j̈́���k~M�o�<�v����.R���'�V��_Y:�	��[E�8�7n9RE���d�7P8�~�dq�Ua� R.4Ӱ�_���6}��&�z)��r���W7�V1�Vc�2���+��>v�ĵ0�э������_9�F$5yhO秼��,�iU���&�zÎ�;tT�K���Ǵ��7�꒤9���+��}����r�/L{���-ϊ�n��]
2W��B��g�������>ω�������t���Vy�!V�C]��,1�e"K��x��N�c|����ϙ�hss�����)���O� ^I��g@���{WřI���<L���e��w�Trk9�x���PWfx	:��&d{=��u�������.�g���N��/I{;�2AɈ�2{�L�;Ƙ�cCpm�;I[���N
3~�㜀|���Ս|���p�5nϗ�و�eDA�Gm�qT�G���Y��4��i�3�q�	�Hu����)��e�������;r�{� ���G�Q���j�x`�ٟ������Ѥ�?�<I��8w���qKV�Fp�剸o�$n/�z*��n�Kؼ��H�Y\�r�1Λp�qI�Xfx�+�v[��̐��C9��;Qu���t��o��JקN�׿n�4�u�kW�R`�M�𰟳�畑�0�jǋP��D�FV��� ����t�TN�[)����e.<C@< ;�_L�^�S����eO̅ ��KQ闌g��Ue����������_򱒖�:���F5<XrЮ�jH�V�
��d��b;��٣k�8�6_�p�������sW�|lZ����dBE���Ж!΍DZO�84��hC70�S�F�Y��K�,BD5=���˂'�u��/��+ ݯR��E��k���M����0����K�,��;�K:��>5[uW�㿖��Yp+�U��o�?Oٸ#OVa��B�uڳ��"�`�&-��S=#DN�?M̎�W �v��qN�.��bF��K˩,�(b�ܿd�'��*k
��H��2�l��ph7.��C���M��#!��QRi��ıW=h)�pnP=&I�+��\�\��S=�d�q@� £FY8r�R��9���hA�#�8a�Q���j�.3)'�t��ES�F��g��L��ޜx�����v��t;�EB+�$�����Ǻnla*��m���k��b�x��L�8�EܵE���u����VLn)W�,�J�~V��H$I�Z�m������t���ч��Dk<�TY�Ѫm��0�B�/{v��0C�SuTp���S�]���p��$05k2xe�p���`�ti��d�Qť��TP���λv�^�+�xhf��m�(���?J����y^65)�*���_F(�� �<Y�+��!���W8���\�Q�Ka�����S�8���Æ2��{j�%�z�9n��2%�~� ���!彩>7s7�k&_����pne��ۑq��	�|��hXc���g�K�خQ�\�����T'�e�d0u)e����P��V���Tъ��Z�g�%�x�L]��w����RYWp��� ��Ԙ��+��e�	CoҺy����Џ�X�	~��	���`V��U�����0�J�w�w �G�.�I5�K��e��ۖ5��F��v��H���JQ��Am��߯���Jd��+��G�3�����������<�W��Ü�fvL_���đXX[4�UW�61Ho"d�q��׾龍���EO!�M��!oD����M0e�J$|�y�x�ț���7.����	�m������ʦ� ���T���5�ā3�$��@Cc�y�:���*�k|"i��	Lu�1�gՂϲ� �h<u=.<��)��+�DY"�'��Ek 8Ez�!��{M�$�<X.a��9m��9"ÌQ�eo�Ja"�
�U]�&Bl��z����A�kW���T��
B��\��p�Y ��)�x/�r/�(ښ1���:��/>�����$`AZ���ñl6�⩍�T���FL�o'��M�n�5K��ι�k�'$�;�Ga��� �ؕ@B���U��p��ID�!��o���h�V9dEB��@��~9D :h���;�������55&(�-|`^nzd6P�N�� ��E)�%}�����*���u�!-���l�ĩ��9�6A�1i�.�J��w���v�T�m;ǆ����~<�ѻ�0�3��?^Wep��Čq'�⢧!I <��ʯKl��l���?�J^t��\��F��;�w�y6ݬ�Z��ut��jX`���90����wf�yl�ڕ"(T����M�V���i���J[8f�G����K� �B�I����k�� `s^�7�m��>bjp��^��=.�ȇ�e�2L�t����A���PHC��$��#�@m�┭�B7�j[���IA�A��)Ǣ�V<�Kʨw.S���r��B}}B�e�D^,�P�?��>�i�@ё��1yb�[�{�cϫ�����o#�Փ5��9��p<�����<v���Wf��8�n,gToi��}b�Jʲ�l�hng��q���̧;�a�m�L�X��(&n�-A���C{3/1�ʔ�`�_	_ٞk?���p�+b��O�a�&08`�_��? �E�T����b}6� �@x�BҀ�t���.��C.ahUn_I\oR�
Ԕ���J��c7+|����P��8��s�U=�1"��Ҫ#��j�C��;9�QH��O�*Z�w��O����~q/�foJ��C6�jAT�eOd�o����`N0#�AĜ��]c�
�V�NV&����8�8��B�� �q���5�t�Z�{yR�􀦘I1���B2��ūꕮ1��me����=�PGY��G����������O2�Aƛ���I�?�@���;��g2q߫�tL�XA�Sf��T$�	�gOo)�L��s%�_�3�d�߰hf��h�T��;yE�G5(�TT���a��Jfϰbq��p{_0�t� �B��SŎ���a8ɖhvi����ުƷ-�N<�"�6����,Jz�9���=PFe$D/����'� ^`eh�Z�d�4�!(�o�7t��u��\�B�h��'h����T%A����FE�<J��wG_�	m�G���s��D�D|�F����#����:&bAFkX��&9q�O�:^�2Ƽ�z;p�����c��|с���6�#���`SK�!�d9C�/� ��m�5>���q���2���/x�=k���)�&����[ڥ��6�o-3��|y]��CJ���̥���Y�'��'BѬ���#��>3jYsA6��]�M<sQ�ԾN�	��N�+mס��ex�����8���M� O��z�~���(�az�Y�_6�-��8*+3ϩ�!�=��j�	��<M��#*�-�5�9^]KN�c�=�3umt���l#�D^0�j��9�D`<I�^�ZO��jh�ң���*<�J��rg��^P��I@��84�ib"�#å�ƐK��*O|��2����4@}42[*э2�r���ݲ�R����0��q��k�3S-1f���̃+q�a�]!�^�` �e�� 1Kd8��{M�z7����,4���S�R��{�؈��S��"��~��u6���1g��C�lU��ʏ~��ڇ1�\����i��@.�ӧD�N����`�U������	���3"|�%�y�1m}���d��;�@X�Y�!���u�	S_跞�\�ǝx��
g���Y1T���PR��a�
��euʞ�q���{�O�����x:\D���W��|�����{f��*o29��J��� Bg����bg�Z+p�.���P�S���Dh���t/��#�?��}�8em��.YZ�����l0!�bt�����=����ެ��m���2'����H ���G*W	5�5Sv2�n�"����p��j�;#(.��Me�W�@ؓ�L�F/�<�UCu�RP�eĝ�˝���ɣ��Е����##�Ī�v�&�J���;+�֔����Qy�I*�=sk�)���SM���)��0�b.,ޫ���f�"?�Jsf�V����+���K(�#hԙI��<ӡ5�~�p��t[�PC~j %ያ��������r=+�-
�Z�y4X^{����/1+�+M!X�"Rd]O���\ߠ��� ҡ��/���m�[����he��-@�>����,R���3�?�h�����,o�~�)���&�6¯�RS��!��g2����~��U]�"p%xwW�y���a�
P�-9�l�W �
wk�+M��_��a�Uc0��Z�ZA5SE%*Z)g6N+���r��h�*o&z����W8�l��_a�l��R{�����ek���Zg8�>�<�vg�H��f��x��w&�]{�CuF�s먉l��96M3K���Ö�.�&�x���S�l�SLm�I�~0�ݙ,�cTf�9�73� 	Ȕ�fV�
������v�Rvf�):SM�篎j�쟓�\�`�4P��i%��hb �ʺ��C�|[�$?� "�@2QB�T�6���3@��B����k�1/�w5�v���>ίG��=��,���3 >���༎��QB������i��A<Q)�6��G�ӝ{���oc����5;~���2��$��$���~��W���\x� �4{J��y�A�4�4����%�r֓]H�F߹�6��I��,�ۂ�F�)�2B�����?X�s���( ����q���n�Wo:u�g:?� �Wh'�q�)�ΨT�.����?CA�x��ז�N@xx�ݶ�ty�9��'�� ��9-�����>b���NA����g4�8O��p�m����皈�߂H@=�߉b��ɬ�ܧ\"��/�y���p,4Yą!�,�|��]:{���>��*Ʋ����2,7����O�e�C��:�l2��wj������gt����lY��4�l��)G}��'H�y�`�@N7r��L�R�m�����q��o���\]���� ���>"WO:���GDIW�ӎ�����@3���m���O�s~�B�7�Vp.[Xd�mF���#��de��u��P�+�.J�<�M8H�֡���_�����&k`8��'*7
no|=����w����`?�T���ڈ�<�#����bў(>�(���"*ג.N�~RE>�sH�3~U��?J_�7��	�����D�5f�Jb�)S;RYfFo������1Zf����Xǯ��,F�Zܓ9B���N�-ppiK)��$8m� c���e��Zv��lx���=���$��)�>d�u�,��ln��bh�@٫+�:j�֢�>G�dȻ{�(�+��tG�S��>8��j��w���Ug*|pPpU#&]7�
��xQ��Q��$�Y�
z�[�K���1�r&Z����Ś#TK�p�BE�c
�KF.|L�������q��՝W蘎u��-5�1���t�c�"
I=��Ư�͎ϲ���Lg�Q�AW'<(T
A�=��1�y����R�`'�饼-�a-�:� 6��tm7��P�S5����q��Ȃ��	$�b��k�$��ZV;dݥ�l��{�v;\��ą��͛�`����Rx��+�/f�B���,�.;[ҩ���	Qj�V?���DwVhd��rEK!�q픜��g��KﴵW+�x����⬛���T
r��r��6��ܚ���?�b�[|�Ly�zr���p`�{��z�|,`�p�>��&TD�XAw+'�G��e�f���}X�R���v��q��&$�k��4�8�T�ٞ��ģ1�ryoR�֫������-�)R)�S��}�_ޱFm�R��܂�\��^e�C�GH�>����0Į�B���ſ�<�e�W�Go�N�i��i���)�k����4��3��'d۩3����`M`��"��c+p���_��dޮa5,�>���n�����x ��t��cs��F5�����kS��:�j�m�	�̉@4��T|�%�l���X5�t�MR!�M��m��?�^.�u�s��U�\�!4-� q�_�J)B���6���'&�\}�a�6+l��\�t�<� �%[��1��r/
����D��)��(L�b>�+��dƍ�v��mi��y�2��*�-��i>�4&/$�%;�X'��n0�Up�Sc�t��������������u$���Wm�u��y�S�b���RFb4P�b���5~�Y�/�+ ��u�JA�aD66U�S�e��n�N>-R��b�4d��eq��s��2]Bf�5�{��'`:�[|v��������lI�mc-}��
��
�+�2�πr�+�C8��>�����S|�R�7�[:��u�hA�e�=a���۞4U��@�p=������<���cZ_��"��?���O̦��܀�.��қ�.k�t�3a!�xE`s�a�)E��܆����#4ɺ���gs���q�u�]�rd,�P��[��X����V�L��q]���+_G/�˷N��l�q�7�������T����H�=,2= Jy���ʝ�u�'Θ)X����Ra�;��?��Vn����:y�һ�mK��r|H�v_���?����a�����,O{��߼����y�q��n0|��J�;�EԹ���q���<�1�S�Sao3�p�jﲄ~��]�R틥�}ڡ���� ��C��|^-�61��^��&[#8��˪�H�IR50�G]AnP�� S�*�����r��`�.�K�� f�b�����?,a}�}w�(.��C��!R��D���r�"|}���"�Ȁ8P��vBVB����+W�rɲZ���z�]=�d_��h��{�.ۯ=�@8�B �ھ���A�L/=��Ⱦ��7|-�KZ�6�Խ11�w��?A1m&������ț�%P��a7�v'S#��||&����ώ��HW��u=�ѧf.b��d׶F�������� vw���_n�{sr�m�ƨִ�>I��s#V��y��W��U�:�0T�K1��P��#����>�l�2�kӇ~,�E��gTM#�ԙ�h��t�A�r�kY'p��1��=R�iw�saM��1ۭ�������6X3>%[�I0���hZ-�~O�vQ��we�r#,�^:SE;f���H�)����Ƣ�%��`2���~UB6��J��3L��� ^���8P�6���*�^�Џ06�^�g脏bG&"7�\��8Y����Xb$EM�yk#������X�Ӄ\�X��"HQ9�9�ᦱmf){�(���:�{)�KA ]c,u���P�����SQ.�m�����#	`*�{\�~<<{W�Sπٟ�M5��e_f��,]��<�&�v�K����^C�|ǘ�[�������˾���u����U�p��L�TB{
�������3�^���\�����'Q���R��RV��pd�̣$�I�� אU'�T��gf�8�6+ubo�V>ݡ��������U�� �G֬�s�@�K8�<��ݨ��C+o8�_�m�"��d�O���]�.a�d�b�+���*��wޅ�Ԕ��;]9O���W���͈+�L!x�n=��HVj�6��'BlS~���`(!�2���@; ���I�����A�U6m�ޒ�n������y;�h\D��ځ5I�eiB�7W�B�Q���&s��xuyv,7^��Kdi ���1��L�R:��ƅ���*�to1e����'�ENr�����j�L�y��C�Y�)nʑ4:!�΢��Y�q���ϋ[裧�K����٩by/^{��Iqk����
��1�Q�X���(�5Ib)���w>�#]�$�Crt�ٜ{j2��oT�/ƭ�Y�B�+�K]��ã
���wAPb=
P���kq���E��-)���]_赒+�u�	������XA�am
�A���Yg��y�Z��H_��`2�d���8P��1��RH���`�`
�q���E�?��ӝ-�xμR�ZAF�!l���M���J2x�����Ӗ����î�su���k�1�(tz�߾{	3�bp�^+:�?$�@�Ua��rr�.��2�Ev�	�O߭{��d��$�2�Ჿ�C�<m9�Ɲ�����<n�[�֟p�d 8%��L葐\[�pS���.���4z�d�]Wˎ�Ǳ�F-r5�D���ϤH��pr9>�?��Y�,h�p~�����$gv��S�8Wk�����64p����
ۈ�D�A|��?+�~�A/QǪ�&���f��WH�c�*/�� C�ܛ��:��Ɯ<p�/��1��G�G�-�+{�-�L.�a�0��}P&��Ѻ�����;����9����_��(�o���?�f0I\�i²��Ax�'�O��k�pn;8%Cg�Je���0V���M�3������i�H���Q�P!�<QO����ol�V0[�2�ruݜ���D[��ˋ5�����{$��Bh�����}��.٘���,�:����!��SdA��ÝpD�A}w0/7��L���{ȳ��{`!��V7"�_y�P���򋥙� T�S!p"�2��Q��[�2d�	��{lj/�ܡ�����[����fH����N�"�����o �ؑ耗Q}柳�Q�`�ޮ��G�j	��v����G�%(�)9��_f���5X�ð�Kx��\�K���m��_�j�=ƣ� �?���g��ށ���llkgK�3�I$�4C�>�qdF ��r�����!�B�E�s�P��L}Få�L�'��F,��d�؞[�U�`jR��!D�G8=��?����OD�q��)n�F6�SK��Hg�Y^��}In�*���}�$�Q��c�춱�����9U	3������S��&�n�`2џ�γ�<@J�	,�r�~K�J ���Q0�{)|i���!'�T~I(sR>j)�L^)��c�!W<\R���s9��V��ϰ\#�~���I�)"e�G�}tCQs��/K]o0uMaK��EЫ�ha�d1�l���U� �O�OW����q	���W/�~�mD������?ې>�Ļ������ |�aJ