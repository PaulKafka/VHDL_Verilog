��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"�ԕ�!p0��A]2��X3�F/F��Z�`RVd?�lL+k;�E�(���U�ZvD����(�9�7��F�3�>Rd�v���"#�\�8X�����P�`p���k)W�1��z0Z���(v������.7OM8�2D��3�-�>�!�ռ��9�OTCb�ffR��SHpΜ�Y�������ve��fm�ߨ<K��v��x�5mz����1ǿ��ʀ+�t��.�����G=l#���H5��}^�y���t��$ٟ舯��*^�q:,1����l�SD[��{������C6���^TBS���n�s�ڝ�L�����2o5��t�R����0$�X�x�8ب��R=g�X��c[9�}�4�k��%R��_�S����Α�v��1�Q�S� �)\+�,�0�Hmʁ=O�<�����5�gtR@~�O�l��"�����檚S5��D�PBu�F?��CFn�X7 �w@�Pq9�Ɖ�]����E0�|I� ��q[��q4��N��y�7����IU���=��3e�R}��nM$V&]^i����.��9�#��Ѐ��]�T��rf95� �@�<�M}6���@)�m��#�1�y�6�\���g�~�����H[LA�`��L<�wB����чIz����Z���P������k�hN��N� '�j%�C���RPI�X�'ݬ5��ֆV����n�tG�F�K���4LE��0��U�It79e��{�V\Q��LȎ�P�S�d�Z,⁻�>���i&�Β��Ir�)��x�S�KE��$���û��L֜��5Ӱj���]pn�W�x+w�D. ��	�,u��xj�o�BW^1�/5��+f.P�;&�� ܔ���T$��>�h�v�_s7�MǼ^��`�i(����4��֡X��%+g+/��	��F�-�Hd�g�j)�>�L���hpy�+���mf����+��sJ.!Jԕ]PR�IK��(��^�Ǥї��X�*yih�����5^9_��	�Nbyb������K�^ H�R^�򨴉W9�b��Z��^C����߰	n��W'F�:��^���f�%-k�,-��l���sT���dTp�q�k7
�5~���S8�������15���h�P���=A4�=�I;���+���S��
��'���ʍ�.�AOC��5/Sy˰�x�iD���Ba��u�Hy����EM5�$U�5&�e����
�H���*	=/e��{����Co��&��1�v~=pQh
��AP���{#ތs�����ʠFW���o�\��*
�-+�A�죒NvA	�����V1[�A�}��C�UL���"�.�'#j�C�Su�j�T�z���Lp������6�)+���:�Y��u�qW"W�t=�a��!*�m��g�X ����t��W���.���F]����b�G���<��1]�G�c�AP�\�jڲ�����md[E��f�
,f��QXB�w�ΰܚ([?������f1ys	���(>�1���:�l��A-�IR;��G�\{�?����_��p�>V���ĳ+lC�)��b��G�	_(�U,�dV���Q�ŉ?�G��$P� ���(T�F��F������f�[ZT�92IQ����\��J��M�����k��0���uC��V��:�$Kb\�pݟz#=�6��wB�TdS�X�� �1w[���W�N��Fz~�����d����×YK��ǈ�H2p���U%;�A&J |��a�o��&�w#Rݲ=<�Y�{
2Ȕx�%a>
��<4֙1���s�r�s���A�.a��1�4�򂪕�����;q3������,��D�[�aɄU�{D�'ӫ�\�歘wa)��p���V�&���L��@�T�K�^��O���Qe�0e�K'�p)2w$��� s_Rr
�:�$���U�UF���ƽ)� �J�%�aJ'�˃`X}�n �^=ɃJ�U�^��3��9���;~NQ=0Մ�m��Q�m���*�ƭ �h%/�a<��䪑Q���r�2��o�p�<<&D[�O�h��������}A#Ot�� ��2+=�H�j�A���5�v6d����]Jr��'4"1�����w�ۏ��C�iRY�ʠ�����M�\k��_��j�{����
����P;}?�݋�Ș�7
W7�"�#웎��̤��"��\W��X��81�0�	#�J�����#^++O�S����y<�et�\!�C��9�ã���Tr2����H+@� *:'V��+��+��t�&( ީ;�H6�Tb�C~P�t��稜�]�_�n�F2WM�����X!��� ���f��t
���qajIu��; <p���D5aM!-m�8���]M'�ը	�"S��{С6>i` �$�ؑDxU�"����܁��y��hʶ}��Ph�?��ab�=mX{`�����§�M�L~�$�2dvݰ��WcQ��_��Df����Nx.�N��4��K����a��C�P��x�ŦՔrà�ۀf����+�l����2��^�d P�G���jE�m�a}7Em������\�!e̣Te?�6Ϙi-&���ãeｈ❻��24~��(�YN��Yݑ�=8���j,���e�Z�g+���x*��C��da{�����f"\�
	���V$u`K�[!�;��+��m��&�k���ySp��n ��J� �R��LMj��Vg|F���C\�y�(����w痒��_�7��>�r+���5����&����(�����m"��n7QN'I�6�.��[Aa���O��ҽzI�9� L qVl�MV�A�¶A.x��3j&����W�n�/��;?�C���#H�tʚa�4)�9�t��/��HH�{~6eu�5�l�S��|m�J�n�#Z�r ��6�s���^,u���eČ0Q[c.m,�RW��7FB�А�
�{Eg�[3+�%�Ҽ�W]5 �s��Yr�I�q��[i4��yv�!w��k)�oz������c�T��I50�ޅ2�N�g��I�\C���:)�����g�����P�U\�*�H~Kf!
�{Y�����͒�Ƹn�uPI��	ϱ�g�ѷ�}E�g/(+�ńO��{�Y�я� #?-W�(��v�#��0<-"�۪�V��A����Vwo�0�+�����V�<\���a=b�10B�c;O�A-�1u�^ެa�d[/��횟���ڮ��Q`ev,Ȃ�4��2<��)����=�Gl�O��z��]��D@<(�&�� j�)y�be���
���@:�t��x������.���H	x6���`{f`S���NH<L7;�1�!��H��>@�tJ�QnW��F�d���r!���{����l��U������	�˪ج�����qD$W��p�SaR�?��7��V8KI�(9 [w�\�5e�Y�V�R����<�f=n܃�)�i~�����O�������R�**��+�<Nq52�X|��ݰT7Fze./t�1^FrO��@�C�:����[�M%�V��d��x���c�"��g}~-��������ɣ2��|�߰�#t�4�/�h�?;j� 0�	dp,������5�W��R�!4%,lc����m�MM�˽�jІ�Y���˲��-�/5�&���rՇm�z�|�:ө�vה4 t~ !Bt֙jo��~h��X!y� 3���B�faIǢ�n��?Y&�W�@�q�s�<�'��˱@#o��-��{�/�1��9Z�X����y.2���N��;�e�톹��"բ��eQ������Ob�%'t[H��2=���֤�or������5�?f�3�u�镢c��hǫۏ��H`��]��,�-;|)'{Qhw�ɩ��m�*�V���P�8`�6"y�.�����B4ڰqbXIq��D��;%u8jD�&Ԡ�
��4i���$o�j�_W�:�a��"b� d�ra���6�Bu&���F�4����{�k/�����M�Y����ۓz��:�b
8��u|KB����p��:5�LW��}3&�$ӊ�E�R�-v�������9/ђ$�߉yj��|]/��r�.,:�& &IF+!]o�.�!�x�|I'Sw�f^.�v�5���m�Ք��e�V.�Ax�H�q�＄͙�"�*��oͤ��;7j�Ί��F�!L'�f��@ �q����è�j�^���Ҹiₖ|�_!;�r�"��Ɇ�A�z�����kg�V��6�BU/�" ���Q�,s�|����nآ��$���n��#IT�\�Wm/H��"gzo���(���]`)�Ν$]gX)6�S?Wzf����K�˷y��Y�mlfY�QZ	I}�#�)��W;��d�A�R6��ᄢ1�(�����,�x�7ͤ(�C"���Ye��,�O���"����yt+�4��@����n�/�-�8�0�%s�Ґ��y�{*�nF�E#���G��P���R¬Z�G���x��E�C"�L�Vo���P�����N��X��?�Gp���=��� ȋ�.�
����F ���J�O�:����X��/,1�!��v���� $�*AV���h�M�y�*+m�gr����4��s���g���|c�R�.u<Y���ԍ��+}E�$p{"���Ę�[����;D1e��v��o,AL]D��2�_u;njQ���MR<v:�3V�5�9�"����M@��6&wT�2���`z�d�&+�����'0��X��z�)�@ɾf���U�y� ��[�3��n��ջ��4{�,�Ov�D<҃�Ɩ��i��lϡ�����Ζ��?O%UA��Q��3���Dr����:*�Yn	za�x]S$_���Y�����n�t�+�;�ry�	��{��}����i�t_3�_5׏�9��ph��x)�мeI;a!?]��=��5U4
�D�f�
���k9�\;%�f̚~��v��3������l{�/�DXx̚��j�M����Q~��	�s	�d1��Hu魈Ov��[ 25���i�7�vВyy��V!��%�&WW�/r�,2�T7�Ur!�- lɎ��b����W"t���;?�1�>*f��bx��a�2�����F��$p+42�*v�����M�b_Bz�@-�Ag��#��BS<(�g���N�0���6��iʆ�jC+?���dۺ�!��������ܷ�!m=*NkztAp�ep���t�_�2�.����#Hv��t��Z�WS#�\�c0/ߨ��+�!�X�x����.�E�3�J��S@cxS�pB4�-vn��?��J`��F� O���mTUc�L\ ��I��#�w{u��«_�0[	�G��ծ�6����2r���*�xl~�����/����N�,$ўw���<����P��o4��k//��.�}SK]$�Q(H����8�	"W�2s��^�v	N��편�؃��c�LI�g#��D�)2����ڿ���g�<�]#�,�N�H�� ��#鱂T�kBS;^�_/�,Ǉ��qjQ�&��c|�Y��@L�İ���^^�=)E�vͥ����k�Ֆ)# c�Î��DҜ^݇�c� O��T��*j��7���)j%WKz�6�F�wJ�'��\�����̤Ԫ�C@����±G���}J���^��0T�{!
h5�E�v�R ǚ) 4�g��*Y�;x*�%2b[{��69�����:��:l�]�u %�\%z>�t.,��uY&�SL׳1�in�LK�f0��~%�����ޮ6
�_���b�����O��� F�,:��9���bѭK[��龦0�&�B�AY�&��m>��YIg��H�z>��¤��Yoo��GC�O�!0���ה|H�ە�&I�����"����=
�z���iRz
R����6�b��կ�w(0��$�X�n��}C�W�`j�Ld
Ce&t�Vϯ	�	U���y�Z���AQoGX���T��-��_�~�"jY/��)�f��0�7��.C4��:���_�����@�������F��A���q����5�*�lƌ}�iɀ�F�9�6�n�n��?e%��e�jlK��Z6����|j��.M>��B/�/u�����b}��:�<`o�6m!���.���6�\oT�8iX�7(�d�)��9y�!��_2�j��\�Vr�1�F'ؿV�+rG����وo6-������e��r��|�+y.���ab�=?B�u��+n3À	A8Uc�2k��![��-l�ܷ��s���q�%6l���6�BOr���K4�P�Hn��!߲`)����1�I�oNxL���Y4~u��e�e`�2����W{*�ߡ��n`~_j�6+慊uTA ���������d����9�}�TfT�T�D�.+G�-�ꙇ��&�'�W����BLm�_�(S�i!|�<�%��[	�;Q��1���&��]Ets�����s-�mT|�kj*> C��v���jh��c	1~�����H���C ���h� ͷ����P�����l�5�U�z3�þq��y��9;Aux�jz�w�m�'��'�q���m���(���c#ۯ�ɃY����s�kޙ�,H)Uڼ"�j_��o��&�������1�dk=`�u@d7G�N�r���<.��Zڿi�H��e��5�{�Sܻu*&�W<V���t��ٓ��r-ԍt��o�aXN4.����v͝�qQ��@q	zzi��ʴ�|-���om��Ղ���y�U#�zHs�¹�I櫇%�w�]+��-(0����ʌ�d�w���=j�>@Hߓ�����{�z8Y2>
m8#��1�Ƚ���Ѳ��~��̅ӣ�jG�����گ\��$6LD���7Ϗ��p˕� �k<���tWAeVE+/:\�C����L��]�]1�]���gn��>kZ�ZKj���'��7[P*1Y�@t�UX�.�_��jrt2l)�I@Ό��I�UHU[���[�'��#˺��r��)�-���ܔ"��3e�署�Wh0�|��b����B�l��B>4�h�����%�j�-� e+�m(;K��:�:ר���{��d���ac܃�q��&Jf���*7��{�2L6��s�[�w]���{�z�g�'�h��H .a�����FQJ����V�e&�j+:��~����:��@E�RQ���E��#b
�H�������eiａ`I�_���ᾫj���M�6	'��N�}Ӑ�Em�$DI�~.����퐖(y��s��BC���q�W���dQ��?
�kj�|e�oW���ǜ�q��s)�-Mh�P���r9�����*�|���k���{&[gE���7��|��fl�Oq9� �"M�Rؿ�ʽi�\Z����������`@���9n-#h���f�4��v��k��n�̊�Ԧ��rd��ьa�k��rc�LI2i�C]��K��Ɂ���B���+�RҎNwiy�J�����kHZ�8V_�.���t����]c�2��L��b�#(���}g���N�Y)�DcU���[t''>�j��
�A�I@7���«eƺ���x�xu�ߘ5kpG6�:��E��NtY��X��Jh�;��0�[�� ���o���0�@�s��d20|"���Å�C��#����cS�LTJ�u��N6�n�% �p��UFe�;��j?`21р$X���Cߺ��Q�f+Ѹ�#p1
���M�w-��9=\�k���xn���c�|�H �a>I5>��~�Y�>��Ԍ�gg�G�R���\�����h���X 5�"}� �V���S��R"��^ Z�
���|'F�Ns��KC6��Ue���K��,�;5E�d1Lj���]{p����m��.S�~�����Vo{�{>&uv�L�W*}d�ڳ� ��Y8������m�/�i�y�YXJ��L�M�2�3G���ʬ�kF�id�nd�6Bnq?,��\���>�j�������	�9e'G2yu�c{�[{!(5�U]�7���S�k����o]���Z�zg^
^��|��S\�<��y��(x?���S�[*~���c���2~��ihtnF�D�&�}����3���os��_�'='�1M��;3*�^�}}mZ��W�J'Q�f�TN�nc����'Xz ���d�۷��j����
72���7����'S��^�;��Iy��C�P���M(ˑءV��:F��pxjȷ �����gN2F3B���r��wZp/|Y�|�a�ш�ʰ�}i���d�L�Jv����x]���G���nL��P�5�#�%��`�c���� �7���8��l�E�H�
����{3�3h�a����!N� : &E���)9b��<I2mx�n�f'~"_%"�.��h��|w��piY�7���˵O�<�,��lW�w�r z�&*��˥Jy1���.��w�C��Bm�7h\RE����gs�JB� ��l�������_�;�|�RAJ,��ƹ.��qJ,)Nξzs ��!�H����`FZ�@(TZ�����B'�� Q��̫�AV*뮊�w۟�m��"Yz�^ASa���hu<��t�3�W�_;�سiçx�↟q�$WmD�Lv��k!r&�Y�=�L� O�1K�;�D��Obu{t���H�	� &I�����F��^�udt��tF>�����y'�"F�FnsF_��ɺIN̈�G�.+�}��<?���� �P�j*[���6���sh��wY�T�;G��Ft�j������Fu#,��81K���Q;γl	�K�i"�n�+���R̊U>` �	|��M0�2�	OEofz	B�Iܫ�/89&c�!|�!�x�A���F[���ēyM�D{�! ���QC�P1szE��(M\��%V�!1����]FWSz{( y\��$��6�S+�
�\k0eҥȐ�X佻;k�Z�1tat�}ɤ����R�g�-З���O�V7���'1����c�w�d	�������skt�ȧ�����v]� ��p�t�q�1�D�?ߐQ�D��#���Nc�t)��Ȋ6(� ���r���p/�1$5'�q���S����z�����b ����Y�l_$ `�<Z����<�]������$��n߈�L�'�E&dq�ȁ^B�.�,mŮKu�c��(��ڙ-.�CK����F�����v ����#��M�F7������}����J��G^���o^�H��R�|ζ,J���E�X���\�����3J�w��)�Iގ8h�G*�wm+j/�o4i~~�n�"��Wv'�Ζ8׻�pS`�YM����zv�jn �M�m��p.ι�y�l�M�%�n��)��% cl�0+���o��m��65�����*�#`��Ed�$���d�hf�=����×u�&�aSv�V?���_⇬�(�8��	���؇f��eև]�Z�e�I�xr�g�z{����ᩖ��zG��G�r}�g�5Fڭ�..H�؇z���L�� b�zJ����AG���጖����u��b~j�f��t��e-3�耑_E�����!����7L�U*lȞ� �lg
��nx�S�ڡ�n�<�h�a��?HLP9�xj{an�zEݨT�ҁc�B��yx���V��m޼�%Im.�"�9���ќ�O�*ck\u��<��,�\G�-#H�;3� �7��3�.��Ԋ���(-��Ȍ��<3�7�>Tu�z��'V�m�ɮ����GT#�Z�|+F���#ȧ�s��,��� �l|Q���Z�tm	��f9Xf��5�r\�祯��}�����!o���� ��5�YҤ^��1sQ+l{8[WJ��l�i�nR���˦����7��v�:%�I�#��4t�bq��#��%��c�u��A)N���f3*u|k��`lQ�8���E�  ��qam\��ohCu�4��	L�p�ڦ�i�������P��S8���D�\4�V:�2+_)u�ɫP,�V��}%O��ݘs��I���-��Sj�nc�>�g&�Ԍ��� q'��r�*�� �-���/����2���B�b�U��D��.�v� �8��D��'\Q��<����35
���,�U+ i#��(e�lQ:/�B���+�I<q{x+��p��ʙ���BJq�7"��ݽk�Z�[M��_6��/s̑�!�4�O�5��$�Z�>u�c=��������<էޣ���evrQ$�#.A�5�{�I�^B�;蔨�Ш���U�ds�Ɠ�}o��Ƞ����<���+�Տ�j�3n����d�Z�N"�����v^.�)!�l��w�V?���N�kĨV�	].D��w�1>,�J�w�=?�l��Յcc�lN�l��x�pj���kR���F|�a[�ӰD���s�
1������s13����>J4�x����5���kN]����>���FH�w�~�=o����I&�`�hf//)��+����D����鷤��H���nw��g�ފ<"�w�oј���G�x*-�������@���?���^5ziJߑ���P�����9M�1��f���O�*�&Ů�l5�/���X�z_}Q$c�$:Ѿ2(b�<���z���9�����ڑ�Pm"+��Ɋ"�X��xy;����o1�}*�PQ�>K��mg� �5eCGD�Ǎ��H�-.X���1,�bM��v���0���'��)*2�mM3b���{�Rbk�:�9���r�ح�kķJ�5H���m�x%L�X��b��^	��7����*r�x��B3���f�X����0Y�w5����C��*e�t��0:ÃUnQ�jD�i["������]�����"X���	7�X�Hg�U�JR�4�'\�1�/U&�`S�F�|ɉ�4w؀����N��9����>��\����; ����\��-dg{�5>}��4��A�x�ͱ�����$�U�-��J�yG���gd�#�+Y�77�Q���
ۧ09
�ܷ�
�E8���7�T��N�nۜJ{C�%1Y���J��#�ִ=�8�"�=d9�r���Kɝ�y�������B71��A�U!����& /P�2���)�`�$+�1�bxlm(j��jL�f�fIv�J�(k�W�:E�{5 ^�Zt{�5�55�B	y�-�Z�����u�%B{�2 ��n�b:�bȭ��_ªDƗ�L�|X�|-�TN\���"F{��?�q����گB��oue��]�|���4y�\�	VL��fዣ�7�uM\.Y��{��"�)n�S������r��ƅ�6�E�����j��E�r�+ڿF$D��OQQv�P�,�lHeR3y�1��+�f�r.�ɪ|��-
l��;Um��;�"����b����۰��� |�4��J/�>�����mV Y(���\���.�{x��d|7uZ�������Ě͈�`�L^&\���&ۃI�2�D��Ke�j��'O���0s怫41�,6T����V�}�3)
��͢7��T/�̀��pL���>����A5�]�-�Y���Ϸ��G����Ek2�
i� Մ�?����.)��ge�+���|�gT.�i�i���8��9oo&��e��-Ƒ' ��yQK7@��6���&M#�4e��U��"ͮ*�r���` ѝ3�ϭ���`L�۾w�J����+X~����'�Ed��Q�%�X��de�(�Ó�3�l����Q]���6�Pz���`�N�u��������P]Ț�~ߤxC��[i��t����԰��o��[����ɖ�KY�L�,�4��A1 XTM��!Pg��9�W��Ð��iC:ClG8���������ȗ&��/V�g$9�h]JX�u����m�_|16'W��d�������4�y�&rS�f^��D��݃\  }��h!Gu�-Gm�"2�?&
�KۺH'�m>_*�
������>�G���G�'1z���@}w��Gt�ɋV���t�!jX����J���	�Y��/ѭ�� ����唎ʙ���G~��k���U�n$~�#1��u�	}�T)�^�� ��A�ž�d(�QL�J���8���<�3!��{孪�����yZ<Kw�f<B����}��a݈�74���N:� � �w��G�+ ���y�^�V�	���.ɰ���i��d�t?�&�ҷ7�Fre�p��Ebbg�J��^S.7�i���o�`��>��B���4ǂ�'�pk[�e�>TY�_^m,���P���TRs��X�򡬅dW�K�3\�x�*��^܋���H��7�;�F���4JI��Ū��<J��A�F��<��Z���Y����Y<�R��6�|]_Ʒ�f��M++P-MN��[������)x@僢p� �{L�#��-W�e�j�4�����I��S���ۊ�.�Q������?`&Փ���}aj=Ȁ�
�����j-�9�M�Ȃ�8}�9���"��o�YA����*��[�c`�=�u<�/��#KDI_��';z�??���/�3fF���V��i��[*�P N�5ŵ������>��QMģ�����"ĺ%�F3�۰zB��/�yJ��-v1���႙��1�5���ǥ�f �F�#�v�r���D���uxpZ�3�"�Vk���@�!O~
�f��.���ڨ9�םu��3�m���� }c���/hPI]�,��z�ъ�f��;"�C��w#�S�6,������1�ʿ����jL��V��t�@J�k���m| �`e3�*H�N�i~�w�3�J��`�o�	���F�@���+��r��kj!�U�
����ڰ��q�1d [�h��D�+s�`?��C�/�xڛ�f_���˞7��!��3���֙�e���n�F�T7������	�4�넧�`��F�9��ɜ��Uo��f,�U�E�r��qm�N������sf����ZE�;�.����F����qE=�t����Ҹ��Xr;������4m���.�������ov�[�a���L��t6:*��(��D��h����8{@�ŇRU��6�����K�uAm���oq�� ���!� N±Á���c f�N�a�D�`����Ӯ�#�P:`̈N���#Ҟ��p�zÆ�* �T|Ģߒ�0��3�n����)��&✦��CfC�ėu�����]f��
��\�DIS�Ԭ��\�LD���hk&��i�,�cfh�Gd*f��f� �`���?��)[ό�Fڶ���F��2N�ʌ�CK���{Ϧ�=����\� �a^[�Uy��iLH�^�=������ţn&b�f��vm�[��XBZ���#�B�-©���낅���'K����֦�L��*�Qr�&�g���V��A��xs�V2���5ԍ~,e�)\1�z��GOJ�d�0�	f�yDtiw��z\F��e�M0~;촡WD�}2Z~~'y~X�AUZ�he�H� 9��>_�b�a�gh<L3dZ0N���5���Q�6Pcݓ�y|^�U�:���~ƿ�]S2�5�Pc��N���|:�W��a�s�)�`)�e������	A�E��DG�vf���,\�00�K,9-�@i����}��l��x��[/�I��֤(�|q�$ux-S�S&�����*����آ���Z
-�I���`+0@?@��1x����d�w*8��e��=��w=h'�&,q������c�f�\�,���������޼=SC�z"�N8�/�����nFgֲ��'U�{,��GJ��F�m��9C���FT�m:
3p����W��fY\Tt�r�H�#̛��,�	�R���ni�� �Ъ�
�[K��E�e�p��A�I'����$��2v-]f*mj�ҧ�,���a5�|����q}�I��Dk�.�*s���_�a�k��A\DzI4e��Ȣێ��M�5y��_�K�5̆����Jֹ��M#K�2c����{+}�#��n$��
���F�����7a8�GV�|$4��tG�w�'3
����j�7�3��~����,�WI�_��["���e��;�/�RN����"��F�΋�q�DP�.�=�ۼV؍�r����	<:%�LQ��?\WT���*�41���=���ݢ�/WRY�*,�b�bT����C�J��`��L���P�1�e���]��
�l$��X��zSXmj[�V� ��F��"ky~yS��o�x!�<Hs��\��ؗ��=bvW�+�D���+N�� ��b6��P�\�z�<j�ViO�#�G��/���j�br���@[�{�e���7�aL�H	�}J���� 	8�i+;	`�K���.b�z�x':۱$/����ŉ���!K�*Z#X +\rq3�im�/��������.��烺���K��r�]�>���r��~b["��.�ӳ!P�8�\O��E��G�
���X��:�.�A�00�����cv�,c`�׷�4�)ܚ���/�?�kA%+�_z�����2���Ⱦ~L��m�����U��7n�T<�-[�����aN�RY�ɷr�t�~��,�Q�ԅ\�y����T�&OqS�>d$ٶ�B����b��L��÷���J��������팆�ˆ�GA^_�ᨉXY��6-����-�� �\�!�ԛ"C[9�����KA,���Vy̔�2(3��ec���)�MD)={*�W!峻�S�����=n�;|��e��_����ԣ���K���-�Ԫ�����(��}�b�����K���n��غ��Wy �fY}
-5������xzѹ��N�I+���Y��S���[���Fy�`���gi���L�oE^8[^���ow����Q��7��F�O��X�6���-�lj���$^#�kf�/�*7~?���Zr]x�48v:.=��iX��b�<��&<Cȣ��H��1�����|s�U�x���.��;ќb��`%��dL�k�h@0xD���Z��HW]2?�z�0>>������\?�jԉ���{	�6�1l���l=���e��N��N�߮ �����|Y#I�_��:��9����?��و�`WU�t����^���2���E�?��Ն_�שG���u�m�K{��QRy�h�w�¡[_�����`X��f�>R��su(����\�e�kX��0���߾�te�]��F�䤿L����jiR����Y
|��G�@*�Bt&R.K~Ϻ��t��5�8��TV���"��)��ĥ�Vd�$1޻z!��Տ�l��AE ��{�\��P���i�EUﬄ����	�ۜ���"��e���l��t	C��.A�4�r��0��W,��y�rf� ���N��c��ۀ�ڵ�;<R$ vmuFQ'T�n��q[��������ڳH��G�H�S�t�Qdf�
���`i,-��a8C>t�R|�`F��_�Ci�C9�p��~4�&w�=xG ]$���{wz5%��!9оAʓ_����l�ȱ��N|u>��ø�Q�_�\-@�>�*8nz�eW�ɽu�W�J}�U���r۸h�D������dϜ�T�\h�����m�`�N�A�d�W����4���-��M�<��{�e���W�z�����ȫߠ�r|����G����'�M�1�3�5�V��`��|C��?WŔ��Io�\�Q��v���v�Iu�����R��E�ź���W���]
hV����M���04 D�G�t�>V�+R�R@嘃Ǝ�����#"�<(�N�bb5}��|J��E�t.�
����, ��@�Up�\�T�\ۗ2��`�p]���Ooiڕ�ܼ����H�H����u��G��[��85Gl��Ce�~�\�1[�`�Ŀ���^�`r���jmz�օ2zRdw@�
���
@�d
,�W�9��o}�XM��Z��c�R�njm��PR��C��kL٣��̠u��%��t�̈C���T���I�����/d��R��۟C����\W�)X�fU��^�@�*LY���W?1�жAs�Z�s��a���	���
+g��.�! (�;� V�	����ړ0��%�Y�=㡰ŢpJ�G��N�e�9����{�p�
f|��k�i<�(J�vB�?J���P�-��8�űȉpۃ5x�c��-���s�30�Ѥ��T:Ntp�*,,��ߨ��f9�]B����)8�+b�|�Ĥ�J|7���#�<��Q�j������t���֔Ѩ��F|�R�2�ug�2��\gGȋ0'���������_�]/���S��wK�/�JR�Yʟ���M�B���Gs�T��H�
��6�@l}�=�JeB}v1l_<n���M��r���,ϪI���xMXS�Q�ʘ:�G�Z���#ai��P(��;�WH��n;�\��:5���ZU����p�	�e�����)/��s�+^����V�J��V6�����O �h��#�f��}��@�^�{8�H�6w��cd�<�=_�1ڭe�2V�e�++�����$�@*�xg �5m�Uo�=�s�N��W�TB�Ɩ��eVg��w�%3|1��3c�<s 2��K��C�Mp��zF�EBJy����&C�'.f�ϳ�+��_����q��R��_%W���}n,<�fhҖ��"o,����� |{�F:{�j]����X��T+9`�>��g��_�l�[�����V�nɟ�|r=eտ�ʺP����(���~P��XS>�����跲/�ī8�w/_�JF&D�	A��ڠ�AxS��9	�%���ŧu\m��1Q]b�UQ n�	[m3RO�Y�!���+�$Ǹn@@f�f���Ǳ�."��x�1&`TR�1QR��!Y�sC\N�4w�ju�e5�;_��W�e�8����0�tQӚu���`Dr�H�4_u�K�~�X�s���/ٖ]���͆�E9�������!;��ug�Y�H-��Ώ��6���5��UB�B}a"�p�����FD�6��MiF+D�8����X�k��aB}�|�-)O熢0M����:��L�ķ���/8p�9�d��(1�ʏK�|���$	��#�Ͻ�u^�ڳ����,�~TNlg�q8h�NȆ�����&8t:�0��UJ�taz�>�K8OQ)q$^{ ^���G��Q�0�� �5�˸�2p��U��`���&��͘^��D0�TS�\�u��N��L
�_���mCEs�!gAm�'ǫL �B�~�Z�
�����2���5C��==ո[o�}M��m:s:<�?�ir#�f�S=
}�z�Q�B��i��PԹ��"LO'.tc�3K}�f�,o�($x�ɿ����k�dݡ8֯��џ@�I�� ��]��Pҳ~����ş�P�Lt��hi�h���?�>*����,U��ԏHa�֭�,hu�.��C�[�r�,71���ɀ6�m����f��Q��MO���BI��y�3[��9&;�$�vn�ىQI�H���_:G��g{
�fH=�G�����[co��-�Aj�4.��7��q�-޶`���;D�
"}��L܀0?��'�XՔ�в3�]���(�k���oq�Y��K����d��!rz���<P/y��ZN ��E<�i��]RbE��F���=�e�
���7	p�@�d��k]���2�>���� 뙝$,ӝ/���\!��܌L���.�`��=cˆ�h�,R�E�bS1���Ӿ�,�
�[`���3y���U��Y�Ó8@�WOȿ�ѷ�q���M��"��2�D؁�0[���.!8�@���K������/�w�����끵�\��{4M�[�D�����d�%{q��DJ$�lݴi]���
�[R%%���Z����$�vI@+%���.���л�1,��2ށ�3t�%�&}	)Mt���g���6@��_9���xr���r��cx$5mH�:9����ƾx��={�Y���LK�M{|4��G[N�r	4��2-�A�nJ��@���QH���t��o�����
T�8��NT2vW.�0D@��ə�T���&i졃�GH�l@0�q^���0O3j��;��^�ԯ���vꢿ����8~��bd;t���čS<>�IsQ�Y�����I~E�e�L��ؐ#� '���: -p]���xe��#����g��l�1���Q�6�6��]ו 7$j*l�U����=|��	��6�X���U�EXc�Ӌ�,�g?�+�ڴs��.Yi��y�)�AGTrM��E�d7��\7�9ȁ����O%�g�K���[e��yX���a��&>�\���P�VԔj� �N�E6�3Z	�Q`K^�ڱ�н�bARk��>��%eS�����Y���*�Rx��~�0�hUn��<�T�~|��1@!��`��p�*Jl��'�C�]waH����{��9���F
�B�2�R�M>5EK�ʬ:5��i1��6/��j+��7�}��dYd��x&��>M��>�����^��5`���+809����g ����6�W�x�623�}��:ڌ!W��"	�i���r�ί.d�b[ �E�������5Jf��Q�`����F�:K�i���� ���'��k�Ŷ��<�ZG�L�Ҹ���l��O���Q&a��TN%@�ߴ�n�;�9�H)��6׳��Lf3 ��!�ي�?��)m���Y�Y�m��]Z:Y��\9&�V�$�+[r��0{|���C2_$����&u�����1�N\)<���q����.��A8`UA��Vex.���(�$�>	,�!H=���$�C�s�9%Q_���;�fU*���x��-�ؗ	�)�7y�&�i`����Nx ~�̋�lrZ�ZE����o���s���P�H�D�����f����>�ߑ����;3��HP%K�zI#F;o��)Z�-C}��T���e�URzm�H��mx�A[Up�|��n��,ѿ۳�֓��t���gS�c殛-�J���V����Uo(x�I/��<�O���e����/~c�w�љUn�V�&*W������W
:$���/B�����"k߈2<۴��f�8��/Gk�H�$i�8;��m� ������zD ���y��E!)p �7����r�
܀�ݓ�'��Ӈ�� u��Gￄ���٫�����?�.���������}J��א��i��!!�~{%���aDDi�8��4���6���05\^���HHa`[;^o�~Gl��{���,{�	�If��ή�
���BM8h�Q�P'�}���nܣσ�z���G��@Ktz,7Bf��!����{�Z�tX�4:�z�fdA��(�B�K��+w'�ky���(������QP���5��U��YR��m��
2��w�<��A$��m��f|���8�G엿:q�^���}9�F�2����(���ʵ�~����L�3K=GD(3��N�.%�1���,�K�� �0��g(�u��fA�6�)]���J�c���i�m��u��E'��y&n1��<ҎR�1e��}�<������<�B�0)��#T�4�
ly/�U?"�}Hػ�y:?���^YW��٦D���F.̏�-�oY�I��)�U�W����ס[!����1��Wj�؃���g�Ԁrs�zq��� �|���?��F'�r��rU�w�7�!W �)� ,����y�HH��R�a�B�OY�4�@l`�)*�c�kZ��V,���A_:Γ�u\�7��8z:���K�]!�~�"���e��1��	�=���]�9���	5�mg��{k9lZ�E5��0/R��|����Zu[n��I������K�AB^x*��~tH�@e��P�?,�;0[/���ECO�N��r�.��	���&�G��$|�@��J��y����}"��(�n��T7n�Xt���0'#$d��|Z(G�������ӑbt�ų`��Qט.�P.1t�Q�i������v�=��P�U��mx$�p��%��MɜF�����_�'Ֆ?L�4�ʂG{���'�!�|��{!�.�.:d*����Yaboe �;E�|���1���>'�:�`�F��ٳ���=��So
�{�*��=\P?�@��ڄQiBE�����0�VV�.E�+6������ɢDI5��T���E����"<�0�S7�Y0�*��L�x�4�2�H˞�ǜ�I��;#?tw�v���������w�g�e!>W�9S�fE�X��L��"E�Ku���^�z�Y�]���M�]�t}�y�X���Fq�Ԁ��z�7܌Wm�5���o�/�����H�B�n��Onè|]�췁Ғ�F���d",
v��mtY��AG����}y��Qʵ�Ɋ>����j�rQ5@�G�R�W
�&�(�ʠ���O�j���:�R���D�^Zs�ޑ=�s�P�utl�"�3|�Q5�d#+�Z��sa`�����Q����
]{Ҽ����$�?��Q�]F���1c&H�{E,Q�0Km#��>� 9q״�2"o*�I�>&��G��sJ���(�R	5���,�z�����h�L�R��.�~{rk�	'���Yq�*�:��BF;5J���R̪X��7�����Ԙr�<��CM|��{ڭ���9�C8P�Q�;-��Oڥ�&sa�9Z��Ȳ2�d"�N�ne;)<U��J�?�]�4[ڴ�9v"[�E��bi�Ā��@hxU\��K���3|lȩ����P���!o7ʿ���H��]/bШ�؎�R}�����h����͎�g�.�i��R %@鏚�9 %�*I|,5^��7���%vq}�K ���-U(�~U�,���g��I6w�� J���F�����+�7)�O$��kWsQ��P����o����d�$���_b2��:ݘ�R���9kZ
�XjT���2@Ը�Qkd��v �ע���(zԦ��}�9����(vGu��ILp�q£ep;خy`�z��.!���b��X��\�<�w��au;�k�e."�+�"��'����Q����5��w��<��7$�������v	}]�6i�
�dt��ye������� Dy5���g���6V	|���;	��=dsPΐ�����9���1$3��m<!�J@&�km���$]������r4�u�A���O�GS�֊r,�D��Lp��'��Z��b��'a�����0ݠ�`[�e�x2l����?|C�"wO�'^�3*�QN��UKS#�P����Խ�����)X�70��������ɡ�����.J��` �~M�C9z��:g�v��͵M��;�j9ņE�\�k���.�����@&��& �%Xw���M�P�@�GX�D��e]̦�Y�4��}\��g[�1|��*����"Q]M`�z6'���VH0
O�/�(��) �P v���T�MDp��6v-�����ls�bDM�����5�/S;X:��5	��j��i�;Suy��sϩDz�0^�
��<v�I���~|�����3���J(rK���4Q���4�c��nܳ�p���ɥ�d�R�`Z'�ayln�
H@q�^�,S�-f���8��&��9xoƴ�F2n�����C.vi�k	�#m��"�KD�'8m�6ZhŦZ�$�u�Z*��*;����ū��.b��o�M_���S/��LR �j�(S���*��`�G�m8+�V�yw����f6y�6�i�Me�+>����l� -*Ef^2���*!)U 5��FCﾻ�퀶D�i&<e.})I�ypt���f)
F�P����(`͡}g�̆�_�Ez����K�EB��4=�O�Ȍ
\���c�]�FcƄ�-Z)�'�r�}\��~�`���A�t��X����$��&/Vd=I�kR�c�G��T@rc�$'Ag�vau)��
� �&���X2���fdpE��|��ƞ�}�&
}����Ą��γ��/����k��@�E8�:Nq��S\�1~��"�T� ���z���"��cJ;ٺHa��4>-����W��rl*`R\����%�!mcbE����^$v�@�����Y�`��
����%���������@	y�����䋊9�{3���]/՗�6�ˡ��[:�a�"u�dl����i-zRY9�]%�Pӿx�y��r�AX��T=�ۡ������EFɩ=R�f����ipvB�V�;�T1_-`$����,��ܾ8T�9�7��tl�~v��gI������m���p.��˥n�	���jwh�h��T��kQo��~+զ���t��l��R6 =|�p�]D<�����Jr��L��g����&�o^}1������N˶�d��-����|�|=�Ae�]����*�{/s�Z2&����R:Rki���Qfw���c�䃭jϡ��'�se���K2�F�-Vd�=y�5`�8�!��1U�)^R�Z����9�nb�O����w��#�,p)�#�Y$y�P��Fg[��C�c�4 Wʷg��r��v0Րsd�r�:ܦz1��VbY?�%_O�2�42�a��5�1`�@m�l*^ 	'�7�Q��1�+Y
���;z���ɳu�Z���Jni�jS�M"��f�S8�:D�I9�������Z� j힊<��Q��0w��㕀�7]�i�6�eS�
)�\lw�O���]/��ʀ��M��j���尾Iu?a��Đg��nqvG�[ݪ�a't!�]C���D�{�k��Pp���JJ샌"�
�	�TK�q}�A�Bv�))��R\���[�b�m7�V��v; dY��eFR����MZ\K��U�]�DX������ ����P�'����ESfik|R)���c�i���)��!\H�}r��k�KC�NW9��h��NC�����5�j�<G�0F�,�D3���8�QLZ�/en���P�������rO������Hj��N���-,I�{�JS_u�I
��G��Cʷ!O�b8X�f�d���v��ۇDO	\D��n����-�v��G�.M���X!?L
:�6i�eu��.H��+��Du'[�P���D�ձD��ss@$�	c�m@���@f��=����ΗNe.L�$�]M��^�	Q'���_����`d2��a�2K(-����/�O3QԸ`���\�g��5k�G�7�����p��n+OJpBܔ�6���ߘ�ĶR�́g�7j_!�N�P����2�P<懀��������M�DЪ�K`]��Q�jL�$7��q��4�]��Y�NT�!�/(�RU�F�w����Иէa�6Q��j�z&[�6:, �?�6��"O�LW.���#�����H���ϪHW�H��gO��]V��y�.�h���ݝ�&��P��V�Vü�2h3E��Y�@����p�]��s/B���d���/��X�c��_���<j�`h�0/]7����ٓ&Tr�I��%�;t��ﱴ�Tg��k�:�S��G;�Tsu�1/�����UtI��B��]U9�"]�Z�ȡ�� ]��b���ՙ1*�򯵌t;�+R��M�j�|�9����QM5ة�K��9D����"H�+��l�~��6w�Q�|���d�v�(�u�3��Ř��WzU����؉L��r��郿k!!u��N�9��r��ҳKX�W��� ����^�
xD9�4�������8<L���O��s6�=G>��9�w�e�3�G����|@��pB"��%>���8�X�fE�`�ל9�'Yx�����*�̫��)��(�Ҵ�R�1��!�	#�C�&^��8LH8�n���(쒐N����a��G�##�X^,)@;��:)e��굞;=��gjA'�`���i^���K�S�:��'�� ��?���'��z�̟�_�J�oE�X��ؗ�.�:�a�'򢋈a��������2�rkiQ�i��/0�}:���G�)8��[����u>�K�8� 2K��4K�JRj;߄)���	r��BsٹI�%m2��q�.Q����jF�.�~�7�)��c|_�E�w��&*/0H���X�-��2y�B���xigZ�� UU�Iv"�l���[�����v�y����-GG�����"hO�By+c�Iq�V����~��Vm��l͏6�?��nW�1�����_"�5�D���Q�l/+t�Tn	.�R�H�J�X'�rO�SBdP�7k��ѡ�� �ū����Fٴ�ͪC���Zn�Q0��;'4=��rL�SO��x	u$BH���h�Ȃ�7��щЌ���-TR���5�%�M|\I�{r!���ɗ��E�H�J��6�&5�����j������-G\SYB��n%�T..M��+����䜀��1�����_U;r����4ibԚ���h_�o�-Ac�1�_f�w�[t-j��}�{�}��k�� A�%Rm�U�Ƈ�K�TS#��ι��Nue~��/�˼@gEL@�U�Lؓ���q���,X��}9.o��� l�EƦ��v���<�/�f@�������ذl�3L��o���\?ޙ���)&���U��@�ŋ�B�Wm�^� �É��T@�ۑg{�lN=G�{R�V��T�5���{9�����*֨�9S/�qZ��n�7Iqc��{�,j� ��{����d�7���&�1��rb(*�.�&���^o��#�X���y��ܕ�d����,�>jK��N�1���в'}�1^�uN��z�T��q�|`�\�`:���mZ={͝1k���V )<��O�Pnp�wk�
h�,cC�f���^sK�s��g�*Q&ia�U���_��r�_!.��REK�J�>�u�3>��"���LhO�f���8=(��1�|�&J���f���\��w�N��y��f1�4�\���:ON|��k�(R#��X��g���_�r��7[p�S\��>;������<�S.�6YK�Ff�Bfc���*����᝘����S��'$��-�w��wf�M�D�o�ز���FeuA���; `T%�Xۿ(�{���!���̇�!گ_��#���34�X���
|:0���B%vR_N����F��K���WJ��f�,���!�mxVU��J�mrm�ה(�?������^�����);&]��n��?��%N�0d/&L��rS�=Q���-�Z X��W�ԌK���
���h��!Ѳ$��ƪ�%��*X�t�u�d3jw:����,��w#�;egG��R}������f��P�u�N���YFX�^��'��i������8\���X��!c/�͜�7\�x�t�'I�\����31���ޟ����wn��[�O�?V�U@9?>a!�kXo�B�`������C�li�����Ǡ��y�痡ER����:�� 	M ��H �������8�4ƮTec`��2�=�i��(������˲��?�uk��<�,b�;�6쾯�(#�ȝ�P&Z/	���E@d�� 0BH�y�S!�`��(3֧$<Y��O@&��=ڊ�'��+���%����l���.�~�<��� 8X^��T��a]/�� /\IF��n_��o �[,ɖ������cO������p�{�}X���K�t��/�t���vc2�,��M�]�i5.�bMbb�$�&WTv��	Ci�q<ʍ9���'�l�Zv�=�y�XS���#K�f��2`�b`u7�`�S� 2�cC�r��T���S�v��&�>�"E�`/��0��`�~Un�g��
��4���9m�:]̾h�����ُ[����3��_5}���VB]]`�;�	.�z7ng%��*�F>_��� ���T�U�o�mP3Prm�nٖ��R����D���f�eTC�̐���a�7�?N�0:�4�by��N���i�?(��U7��xڋG��^g��i4T��,1��,�R�L-�_J�L�ِ��T�����v�X�'�je|%U�3��O��>�|O�f*C�����N3K���t.��҉����D�<�׽����<8��1bOX|E��yp��p.t���E>�?����M~���,?@�x/E��+����vӔ�
w�b�V��_�ӀH ৥�r�:o<OɝDi��Y�%�DW!�i��
�п�؀�冩��@�E��@��S�v��<m����=J�;�J������HR���Dԏ���>�V[�-���?���͗�3\���������h�}�x/�Mʶ��T#��j]��E�z ��t����v����Md��p��r)W� yH�E���p��\#�5d�yU���\_���c��j��J�m�f'���� ��E6u{T����轠K����, U4������O�� 5�@|���&��$@�l������D�n������te��F|whA^�.��Z��á��ǭ|
�ʛ͇�/�0�c~ER���yׅ��M���T�*f�.aXN��4Lİl��$��2�oW+~S��Ag�>�d+x��o�u+�\����/����Ɇ��P�W��۲Y�M��I��l��]U��B�]Z��q��v����ϲ4׹h��Լ~h�S$o��|���T���ܕ�8�>|4ȜIQ��?"Z/�Y�S���Wz]#�ϰr�S�s3�� �׿�9��9>���C㾮DN|B'U�+8��7�er�4F�G(�wQ �����]�עC{� @�DOU2��*k��nS��p��3���E��6Ay���(�< f�� �U�p�����I��Fc����iԲ^���O[��	�9�R�?��2� Ῠ���V|�nsS:�����0�$=?o{.��<��м��<���e���`��?�"� ^A4����Y>����W>˩�Л��s��i�:�Aa�3��Ò�JX{>���OX�^U����~�x�x�%��(1�#��s�m��q*k`D��������<.��IA�����Ol���^�0;��o�È\�enG"�rI�I�)Ê���lv�acn�p��}�^.=���F���u��3��:G����s����7��>�S�4�1T�	��;_[{��(è�׸�Y��%�����Ԅc�&��N0��8�^	��r�.�Kp�t��׀ i�`�+��zVE�,�2Ҡ'��j��c�8(���K���_8Kj(y}IG��WΕ��x�L��L�9�������c���|�a�����|�&aux���m�O���#W���~*t4I}#���bZ&�'<�+����Ӊ���JИZs�S9՘�;Ҋ�ִ�!d��1J%�sɯ5�=�k)m7���s�y�+~#(b(���H�D�D=�A$��~��6�H�A��cR�W��C���􁍥��#�u�H;��5�BGQݲ���cn�C'��u +�B�iҰ�3k"��>���3$5�߫M���`�]���J�?�F�e
ޜ��f�ꉱ����`��CQ��aM�����b*�߰�3��)[ ��K��g�%�mf����(��Z�@�� ����6�%��T>:S����ς�V��l�T���,(�d'��G�����r��w��[H{���-�7X�ΣR�E������f�,��>�pzdx�׾v<os(^̈�7D�<+$������Ѵ�{i��]^)���K��o����:@s�~4�(A_�Aiey��j�_��b�PQBԔCEb�!���!�Bp���7�-���3�LK�������6[E�b^Ȅ>��`�����!*e��V�;�����ce�)�V� ��_%�L6���v�w&>��[���v��z8�ҼV��a�N�[<���/��;O�Ʌ�4D_<���)h�Z^uR!���g�d��)��<N�BT�06�3(�RC����-�A�1�Z+�O��[�G&�N�_h"\�H3 wN���?T��d̵;W��&��4߂��Y�K�1�\3���"n��_�qP�xjn�w�7~�i�f�zmyxv_�R�3NN�0^��cY��<��e04^�ZaL�k4z��ض��$�jD?E��7�"Tb�Gg�'��v�}��$����ǌ?ƪt���܆,�с?un,
aO�v욘Y`:�X̀�bncɶ_C�fٿ�(�q�G!��� VqxS5�Пw���#��[�Z�£�=��!X�b��X{���7�V�_� *w�3o�>�af驼��㾍U4sh�&:�T���j���c��� 5���@	��X���ceq��q}��sU��8��ܖV��������&5�}+�W%�ܮ�H���+��'�@9 jT���������:��s�ь]-Ij�gJ�h6�Hx��`v��UlOh;�-3��S��_���3��{�y�q��+5^W�{X�}?ץ�!��")�|�l���*4�	¨HJ?8����!�p��,x�1��1�����z���R����֍1rz|��MQw�]j��t���>7z�9�+6=���ś]�����V ����}�f��}ZKCyYWwQSo�e�W�$nR�+���m��f��n����4��J܈�����X"_6��h>n���lEPb�>V����/��ln���o�T��@����z�%���D��q�H���=�;�*+	#�B��xv�sN	�[���[I�7���<]qJ��@y�t
�}�����G����'pTJ�Py�!�B���:��*=yH�n��#���=��٦�n�o��9�Q��k�J/��z߷����\li�V�6��j��҈�z�G'ժs� �Sυ�v��(.��4QUy�?�Y�9)R�&-�}������6
�*�쇩�'����c؜2��Q��UO���?�G�8�i�,�ᒌɕ#�R��2li�W���A0O"��o|:�rMO��k��<�6e8�@s{搳.��u��^�5�CK��� �H�ͫb%ik$��q\�T2/��)�Vң��fh hd��q����\�m��"�c��}50�)��O��+=8��Wh�|4뺥�xr�@h�7N$z��Mbڕ��.��<8�K��ԍ��U`�R�;|�e�,�x��Ī/�C���'�p�=�`��hF��m2�Q� �2��o��zu�PX�o���G�O����
\M`�����7}W�d�+˼L��ަ�+><�n�I�֛�R�r�mo\=J�ZGf�_�NU;��CM��H_���+����J� Z6�~��{G(l��}�� �����cm�mL�)�.ꔉ�/��+A��2�l��z@Vs�AF�?k�q���{�sf�h7�n��q���d���ko�?n�ּ����c��s{���p���J�#�0�Q^����x$�#&�[�
HVHنu�������.m��F)*����)O����X{�I�T��"�eh�J&����*t�����%�uC��5_��N5L	�6�� 9F���> � ��[L�G��k8��a���d������m��>����
�Y��G��]�^�U6�2��\�� ǁ7�d��ۨ� ���a�Z)���J䠀A�H��K��3�7��@fx�M1��o��.�Er�������[��d^��e>���-�/�����\�����7�����Sg¦�^�јs��k�^�;{۽E�6.���R�~��z.a�������VhDP4� dCny�=s���c��+5�"c���q�_7�i�o����m�激����JM�"���N:g��Nrq,oo��4�9J%�ƅ\��8в� �*:���w���&��߄�|�~5j�Z�5��_�M����m�����-dF�A|�Uh~/OJ��u�����{�:�ذ'ǿ
�m/Oht�����)'i �ǳ��y0�A�o�y�z~��ݧ�9o�XV� /�;a�4�1+5�����j�����	_;��B�5��kԲ �^0^N��Z�6��Ԗ�1r���]�� b����5�³��#5 )&Rw��HP�G˧GSY��E(/{� �0ǖ�`9s
Io�#�4�������g�N%\
N$��*ʑ$PDG��2T���Aeb �H�Vah���D�g)����\�G�<�;I��z)N���@�F�u�1�ʿ2�ۑcN��By��zC��l�{�[��HC�a=1ݽ�u�rzT*/�������P�6���ڝ����1Ea%��ͧb9�f�)�-D��gu�cߤ��Kǋ~��d�K���Wi;{�H�N����x�j>4���P)����!|��ݺd.��M`1WD�*�b1� +�"�L�kP���D�����!�K�w�o�Ѐ��f�HP��gHO=ud�Ŧ�
���'B���H����z�]k$Z u��|�`q�x�d���a��_�$*������k#��N����?��u�,U�J!�2��^�g��<�!=#$1���y�gi1�ٸ54����&4͚��Jէ|";�r���lL��Pi$�lVҵ��L�z��7*���#(i\f�(��5ܶ���������3���6P���l�쁅X�Ǳ0}��/�8�Y�Oyu��@�>!���L�/�����b�T��ΌNc,�/ޖ�̝]6k~�}���_��>ubI����ܹ]mK4^�ӡ}�k��z��e4�e_����o��H����a�[0TE�8T�##D�;dy��c�_�{��W6ZE��w�dUz"���-�*��\V�i��>��߯���� �3�zg���]�>�mU�E���I�eԠ������o�_��ZU�flܐ�(ǅ�3��CL��w�-SS�
%\�-QSz8 �ו�%�0���]@��fQ�g��8�<[q�)l;�O[pK���t�YJ��Pxoi�N9G[����Xt~��'�R��c���n#=�0�!��L!#[�T�m	��h����X�31_!^�w��<x�nk]�i��V���O���sg�Y����F�kp�2e��P��>�9�rtB4[%2��I�Z(�J��.�S��L�T����Hg�7��ƫ;���MĖ�� mxcæ��itij	����� Z�g�0�D;�޶O+�t :�;	�a����2�D�����h�-��Q��=�t�W�|Y���\�W�a���b�)	�Hx��;��x�So'U�����E8��f����t[�Ol�M�=���N�s��B�.�:9\��C��ܺ�
�8Rjɸ��&�2!:^d��g?�(�g�5쳁�y��F'M�M{U��Bzw@��z[X�iDu�9dn<~� ���+��[�AH��w�W%ق_�q�*��%���|ڐ�&��Ͱ�ac,%X����iK!����
��.q|5vxo�p7��?&�y���[?!�3���*5x��H��LA�P����	B��?@Ieo���|��Ş�_sX#�:��8�+�GB�b'�f�V� m���2ZP�(�yX��XzI);�2^�ّ�5e�$���M���f��g�	������VEך� �I]���D��ط5ъ��L,qi�;�*Ƥ`��y60a<K���3���c�:�&h�����b4wʽ{>�ܮU�j�BUf1�%5�FC��� ���#�%���M�:?	��tC�n�؛���F��N�gϧ��-1�d"j�h�S��f	d颈�i��4���&�C��е��qٜZ�aBꧢ^�}K�_\�XA����K��<����m9x%����R�m&P{�������b-�G1�1m����;�>��@*���D�Y`	s��\{����4Vn�\f���y�=Զm���e \+�����Z���?ĜuE�]��+L> �&V:��,�kK!w��O�9���fA`T@j�g�N�Y���A΃A�`={�_�Ƙ�63`$�ٞ�qIE�����@g��h[(� ��N�S��{�V����Bve��cN��8�&w�� Xush�t��U����s�(-c��'��u"���gXW��ҷpH#�m�k1T��Ô&s�y �� 7V6��$c%��g�W��Ƥ��Vm\ڦ�1@�\=)����EIؾ��"#"~���P� �1�.������r�j@d�V��RYܢSy��Jw�_�*��?Gu�Ö�d�W�����hmt���u*�\:ј�s8��H0������+1]���س!#3��W��2��Y�.���=�v�RS��'2�����{���ox_~�
����-�d�0�nP"WM�ƼOXi��%TO����k�:��j�|���A~|��AEZ,ٱ-+��vx�v:"�:��(J�~\�4̟���[��N�7s��0�y|�"��!�@߃�8�v���:�ހ/ߪV�ӭ��Qd`b����N]���k=��Ye��5h&e��ʹ�f@w+�7���5W��W|-PDw'��\�q�#p�������z�� �xfx;���!��^�ηH���xN�ۙ���.������$�>��B�PM��7j
C�.�,���h��������CCQv6��}���g�qjD(�Za�	>�L-u��D4Ɠ��h3�����=#�Г.k����r:�1B 1�ӀÕ�Ωԃ��xϟg廡~��"h�ǡ�N���^�0.�p�ם߯��o���>ֳG���)����=_��SM��3��t+�)�oVr�+�H3&�f\X��b]�b���xU4��;aг�ą��h�F�q66`e��Oz��W&a���nI��V��/7*a�w~�c��)�y������c�EnΑ$&�Ŭ֡����}��������QZWl�&^�n��L�P���<qiC4�P=�6�-
�����=;�e5,V���Pk���D�ӀZhC'���A5��V1���_)�`��S_$�cݡ���m�R=���]���0�OJq�()W�m�����r�ȍ���D�>Q��܄	�"Υ���S0�CN��b(�^�@�+M��:�ӎ ��O���ׯt���%uA�g���NK��P�'gDj�F���x����Xr�|�N@���N2"�Zl`�a��(���m!��H��\��ҍ�MV�q9�}��?8�v��H��:zIvV���>�j;�=U��֐۝�M2���]$]y�
��פ=��߃����8�����<�LԂ�qK�\��l�gD����Hf1�69�|��쨶�ow���#g�I�������)���U�ĥ�	�@����pl�8������B,�%��$.� �Hz��17�%?��7CI����
d}��jw�P�	Q#ax<)�ۯކ�������2��	@��y$p��*Z�Z�W���PzC�#&�ݷ�V�*I�� g&�P=ћ�@�w�S5�_xV�̒��=-�g���X.��R��W��G|��?AB���3֪��	(b��[sx��c�l�	��xa����3˔FI`�e��x3[ڰ��N٩�W��?���V)�ۭ�@�����PF �4�wrR�z��#�5��V������͐�
��rj��r����LزL�l�im���l�V_�fY��$��y:����(��0 ��9}߭�M؏\���?S��U�E-h���i:	u;�ص���c@���3^�"�g�����wX$6?�,�F'9)�/��>����@�u��p�|�h��ܙ�,Y}q\(K�a���O��b�P�w �G��� ��1f�)�[ߥBl/�K�l���B�ěY�����dCmHr��zҿʢ����2Q�R\�9-�\�7*d[ή�}�>S
�!��taА�i���J=祟X�|����Wc�6z7aC ��ښ�tGчղ LH�P8-��L��(w�n��2mω�;źb�>�\2c�Y��!��l&5�Yȸ�Aq�m�D}���R�.��.|��]����}r������y\ը
h��R|Nv�Z�����B�V�:
~U�j`���M�R
�(�*
i�3�=��R���g�0��\�N؁QI�f��7��5�kP����X��(��A�封~cN����<���&`B�i�κ�L�,j'����*H��p���[��Z˪`��a/�D#��^��ut�`�o��w���U���hخ��oC3E�{��Z��j�j��%ı�=`&dJM����p֠��Y-�*ղ� �����e&_!�o4$3�0uT�a��v�g�ij;gX�A�,���'��ɘ��r����O��"�IM��Ӟ�D?�}����A�х|dL����4�M:���5I��+Y#[E��4��T�B�ѐ}>�X�H�!�&��C/ؘ,��
��j�NU���HT����TT�}A���Q-p.)vl0�����.4�� ��'�E����]����F@`���Ɖ�l��դ����>���V�?�r�� ek�Ps��]l�.��P�ʋ;��̇+�n�_���d�}��[��J��/�Z�X�[qv�d;3�5���Ʊ]���^Ͷ^Y��ñy�1$ߣmBL1	�V��`e6��]���*����,�0��ѷ�^Tu����{��O�Ց�6��J)]zk��5 @BWB��x�-�~h3r�C���c�M�pD O��.b���'�`]�L�������:�/y������b��Luމz���_/����n>Z�)�d�iN�zyt1��f��y�R	������
��c�^f[ͪ3w�E��7Gt-oտM���6ɑ���:��*S$ٻ�����V%υ�{��ʂ*�]�2�̋��[&���&�p8���8��aB��֛ͫ&6b�\�[ǉ:��B�Z"�z�W���~|���xRe2*�>Up
.�\0��.G?^�_&u61�W�H��_�� tj���u-���+�BSOS�۲^1Q�*��l���{i�����)	*b���j�<���-ٯ�-=�O���5��]��������'.��5W>��vm�&Z����^���ٖ0T����75clHS@J�G_���*���`�훍�m�������ʪbm��6�F��v�U���:|��HS��j �?!X���f&��(*W���N0{!����B��v��:Ble��� �G]t�}����,߬�6���s�p��U����x/7^&�c�a�r�^�b_ܭC�/��g�e�p�/��ѤP�y��q��<[􁺴��V�?mBs�D8����j�90`�x�Qv�+s�V$f�S��G�fl�y^�������#4T�L^�[h9�6{�b	d	&`�(r����TX��Z�95�\�I�@.���e9����A�vdp��xʓz��*d�?j,gy?*e	`-� �*�)�i4]���/�0��5$�0y����I7�������&6U�
PP�� �}�3W2�p����m�J��%�_l�=2��~��)kÖ��kr��JeWq�\. b����QK�>��+�ZM�ץ�y>I�`b� '�ia�r��C������{X�s�r����a+wi�/�f�����>�Z�c����ͮU� �M���$�2�(�VF�y���w�d(�[L>t�R"��9�zs�U7�2sv�& k`����]�P`�x�sQ��?���K�!��?���>� U�Ub)7*#SQa�_J¯ɥd�8)d+�c��f3�H�g>Y����C�܈����q��YȒ>��!2ai��h��$4�C��pu��=0����CE�h%�*�����j^��Ek��j7*@�Z98������)J�ֺ�(zȫ���W:�R�/�E26��re�EC���1V 5����H�tFϨS#S��w7M�.[R�9�p��TrQ�͈gh�V.�2���9-_����T�`'r����x�+=	��w^J�3�.T_��
N8D�!~谒��� v�����[�H�δ�9JŸ"~�L,�s?�  �>o�
�y7����F]wE�m�6�y�<��\����a�<�dp��At�����k�6������Lt`� ���x�WS|R����7�"Kg �]6��������y�o��O�[��iJ�8�FOD̀�u��9���f�㬤\������݈��e"�����'WAA�R�=�K^����1����%�/�c�#CbHa&�{	�L�jA����\��f�-W��J{v�5��^qDd��1H[���Nm$1����\#F�E�l�)5(�?���ߞp�j�9�m%�L�G'=��u��H
̼�5�b	ng/�+����4p�˃|�a��lv
a��4>�M:!t8�ef���Y ������^����� �KZS�<?�l�������})���2�����G�p��'3�`�L�o���?R�ߋ����w�����{��c������y.����
����})f�]�#�H�'H���.D׻��>�c׈1����e��z�ݔ�-���������gM:��<�$���MV�ey��0��̅8�5�Z�i�S��e��X�Kr~"e�̨�1��@���k��NH�4���� �+Ip�~�‿X��<�u|��px�gcw9q
IY���p���ח��_�����N7�4z���x (O~x U��k��( W�C��ݧ"�gM�m���B�W�拮��<�>���U����F�#�|ػ���l��Ma���6���6�o�#u:�B�HS���A�X����.<)G_�4�Yg(�<�b�&�,j��{��Y��{�B��f�t�W���tTT�(��_)xxi�?v�\��l8�k��j��+*����`��l��j^�:�x��._C�9yC���P�6q�m�U_,�PI4� ��5Oި\4�� �O���#�=k
����V�-_56���~��OmJ��Gb��q ����%2jI�YM'��R~G�vߤZͽ/�X�k���UA�mKi�w	�����du�k�*���h4sZ2w��(��+�I�� ^Β��v�4g9��9������Mp��.&�C��j�Jz�^́�����o�������t��K��	������0�֭
��ҭk3�1�^����xQBq�|o�(��O0�����S1;����}^q�vZ��KB�dc���+%�	���p���y�0�D�W�:p�ͭ2o����pzˏ�y{��>�(5�R���ؕR�s�ڹ7���<����j��p�VE	~<����n��ڍ�zW!Y^�҇ܟ�7$�v�i��k�B��^�M>/�y�g��U S�����l�ƉԂ�'ͨ7��֕��SG�h�j쾡��JEj<d#��]3wA���<���}�ʫ��h��LD��^����v���Ah�+�E�sf_q�t\t;��&=�gU��{0~^��tȄ�V�W�um-9�I`�'��`^�i��~S��A �^�%z�%*,�X�w����\ Qz���-y��DQސV�,�(e����+�2���M3����&Qu��i<e>x|o�CeqD�[p��\�4����)u��|>,'-���{�~��U
?{�.x������)�7�`>.C�r���� ����_L���(A�Ε��J�/n�(�-φ�'��1�VT��8���?` 6�&�$�^����p�a�}z�|Y�j?WW�1��:Ng®����@ ծ�hEs�e�w�-�T=J����]f�4ZN$Ј��>!(bU�$u�Օ^���R���'�5O�zf�[��<
K# 3W��j�_�2��RR~��D��zV�6��Z��Q͖��%"��x>�L��� �t"�ජ#HE��s�,��-S�co�w�V�g/�Sa���,\9f�h����-��&q�Y�6z8A>�Z��o��?��=xn�ݗt	�����XD�.� A�ط�)�.�=4X�`# &�\;7�<戙����o'������0����{/��̸d�ݧH6�_o���IP?ZŇ�V��Q��|�IY��(�#I�.�Y��u�Ҥ�LSm�buB���u�bPj�H�����ޏ��<�./���(O�c�7���_В�����#�RɈ�KW\õyX�ޥ�����%}纯Z�Vytp��4O���g������>�����`��>�I
&i������F�Rdћ�D9��aЗE���;S��U�!M�|J�gL�o��;W�܍2mS�P\�C����o�d2m��MD�Ϯ����́YK�k��}�\(��e �o.�\%&��ssn!c7��%enV�f˼� �_��t�m|��l����ۣ���?l���1���~��Ԡ���c��	Vlw2��7v�8�����-�RJ8�M�����)O)b�T��+����{�w�x�>����6��Ⱥ8�W�W���F�AVn��������'C�\s�;65������Z��K!��t���2l�M?L*?Yc1ZB��|��@09� �J��X	�f��(>�m�j�;^�=�+����9�.$ǂV�����s��N�𻸻�@�$^��|oxEK).؞n/���*?���D+�����2���C�#���Ni�Z!� ��5UkO�M(�6�O�T�N�~�}4�7��b�.�x�zz���������ǕA�к|� /�Xc˙B��Vw�iG`<���Er�����K;� ��ۛ��2 cX�%��#H����ү-{~z
�Nj���K&QT�+�@P�x��N>¿��Y塿
7��:XҰ�L�Hk�9Egl4��@�Sk_6������'�J6���(k��O��]��aRO��>)��1t�w.�?�FJ�Q��+>I��N~yi˴�˲������kl��F�6
�t��|���7M���xѯ���J��|��@�A�v��e}-�����f�a�*^��L�$ms��� p}/Uv'Q���(�6�K��q��Z��	8��p��"2>�ZT M���W�FC³m��~�.^U�.p�!a��Y�
�����	,[�L&�g���.�s�}{}�a`k��D?J�^Mwqz�v�Vb�־�����f ��\0��"�����o��5zR��7 �\�.���
�����HPbP�J��B�D���6ܝ�I�ʳG8��)�~岍�ԻyR�<�!Hœ(���ؘ�6яj��NǬ~�Xf0����Z�v�Zڄb���y��f=M\�-�?9I*���-0�t"Ғ҉��(�b_U�'2�G���4�����a�1�?.J�c�L�J�'�g��-�a�b$��:�!�.u��ą�xϰ�re���x�Z���&����Ǿ:��)rXo��2[��_ ��Ty|U���G.�w����
�R��aWQ�d���hRdj����H�%{0�mE��^�ښ��غ��م�(Ž�ei����@d.|�u�K�v�t �g��Ě�t&f�m��Q���Pjo���\��Q��.�ڕ��8~aR���!H�`��r�$H���0s;��2g�Lip�~���&_:oOu揫MC���(�X\�ݦ�k��+���X��ãeI�r=qC���^��Q�1ɬĊ��EF#Y��
mO��%���W�S����}���[z=f�兗]��P�%���=diVRwO�' 0;K)���yl��vo("Fn�ǋ��l����Fn��R����F�5��`skC����ʭ�� ꔥ��tO�TXf��׈-A�&��@+�``;�[���)�b�Qu����V_<f�&�พ�.~�E�*y:�xo������o�'#�۟C6�[���a|� ��UJ���?��&�D;� �� lcj"�+�#\չ����@�LQ6�;D�ܾxt%Xe�Er��*.�SB5/Fm!Q�C���3�8_�".{�^0;�di
ב
�7,rTz��D*�W���s��()�S�>�JP�xt�l�|Ze}}A��'�Ɂ�[s3��������z�u��Dk/��-�e���1�p�NXI�%����>x�G�@��(�g��d�D)br_���J�ۨ�I�̢�@�j���b}���0��m��S96�$Fw���,������[��[�}&d���[m��d���˫Y���P��~�^"���M�����b��(�߽������IF�9+��M����%>�l�3��|�~�{��Ὃ��û�EYQA �g"���x��P4�tƪ��C�i��eFuc�EA3�OK�2so� `#���Oʗ$���p�i�,�Y`��I ����;��Ȯ ���B�'Ņc~=�1}����.��I�߫���孪�׃b�a*��?3o� ��X�{;~N�ce�7+����V?�al�s6�($1j�!�˫ `/���'�{�x�=^��{�ҍ�)�����?&(Z�%P�9_�E)���q��)��7z>mr[%�����j9�e�;�]1�J��/{g�[�<D�����)"��R!�V�N��3����lN 97s1s��?	"C=�.u��AT���Wc������MB��q��z��
�Y��"���n����g ��i
v�>�&<C��@�=��]MӉ&?�b)�X�7�\�<4�}='��4�1
0�q����UU8u�t�Ҏ�U?5B%}��5Fmi��*rc�	�B�p3D�se�ʏ�@'��);�)L�<Th2j��j��Z�u�9�O��Sx~� ��\/��X)	ށ��Ȱ_��|��[��ddٍ�����O*.��]l�-�8�����:�
P{&�XC?��$X��і��M0
G�W�0;��w5���	��c�
2%����t��KX�ǩ3��wa�K��7����{,%��C��V���W��3q�h�U�V�5���`���0!?H��р+�0ׄޤQ"q�q�4��sR꫺*�)�Y�G�^a}��<����˾�AM!I��m�F�gP��oZ�Z���F�\�uJ:V��`Jyp�[�Go�	�����4�.1��֣�{�&=Y������ͺ�V3l��ӑ��� ��	��6Ng�5|?�Y��L�#�g����dm�wjf:��Y�<��o�v Ԡ]Ȝ̪_�V �'�H�l"�����
R���+���GS"�b�OM�!4�h��Y�E���[�$N�Pu&����L�̆��6ԕCt�訅]��d<����#4��"���v���!n�0��������T$���V�l�~\�:����UPR��S%��f �<�-�����D��	��m�f{�j}�gZ���s��~yS�g��?��	xz��x�D$�c��{''w�~���+CL6}bZފ�A6�ֲF�l��j��������Q.WȦ��H&�L_ٛ�^aA�I�o� �ӳ�S�N�yL֎s����\?�W|��>>�����r �ed.�	�r��3:��F]��\�Se
"�e+��ʜ����'9����L
6!��7�	4I;�n�:U�@�J铖�ظVN�2m }4�÷մ����FT�# v�������f*a�+=3��H&���s:Z�Zh���+7��Խ����0�҉)�82*)��ol�;V���B�s���W�~Y�y�7ϗ�o@Ԥ����F<&~��y]�3,	Yv�Ȫm\�6�h�#_���%
�C�<'�g]��V=� � ߘh�^_��_��v&B(cC�D��hV뷝�~>���>���v(��ka��㟞�K�7���:\�C
�-	FTr����:��iz�Ќl�`��4`�N�*�oM���Y�	�lp�fo_�0W�m�O�E�������W�}�-��nR]��2P���3����^�e��A�yXQ��e�%�n�`���QU5(��k�UKE/�0/�K�@?b��Xt��Q# ^H��Z���::L����
�)�h^t|I��T�")=�h�<_ȷۖ왩�{���X�1��\�$�K��E�,���i��Pӏ�%Qk�g 2� ��B[-�/�$�i�(@�,�R��}R���{Y����ή��,uZ�ueO狡�w�0щ��z�f���v����+��t^�g��|��f퓜���6|(��m��I.+�e��s �؎���T�$�E�#[�����;��2�����!5 �FY�LEq��~`�N�`qIfe|q�u��PZ�kkIķ�P,Y)�%��G�*i��?�b2���5�+�"�&U���0��I�z�����A�3�:am��2�ӯu�[�/И�H�,�Q��g��q�����gW�=��}��Cɑ�9�o/�a�-[�F�&�iM�/-�`�9b���	��#����I��T<0�����]�R���Xo4+T�)�X)�/�9�|r�M~��f�L����e�>8�Zֆ������Y�x��������_c�W{���F�;4�<y�����o�[���o�TY�����-�1@�|��՗1y�s��k�ۢ�����4A�im>�~�qQ�z��i"������:��:��6w2�f2�EU�0�Gs�k)G�Z�H�6w�66y��Ө��d����MH p+��.�+a�M�/?b	��1뚕� �O���rg��x���ɢf�����	K�Iw��	�e�����5aN���K���8��/�i��:wD��������T>7�ub���d�r �/��0h�WiC�V�^�W�?u�o^}�lw�١p��|��|K�8	�K���������D�w���Acpa@Z��첸���!ZĻ^��T�����H��$ۚ�K�v��V~���׸jR���
��F���zX�cu�l��	���F������1t�ZBt�Ĭ�?��Eux�Y�&8>�-�#n6�p\�,o�\�z�
�p��깗�/9��	�x9�:*���J!3
&6���Y�i��7V�����θ�4Ml'���\���(�=i=��O��1����O��ѬР^jl���dY5�IG+��8���z���'��W8EW sۆ-?!{y�xnOId��d���[<�Tz���D!���E6ȍ���*��l�����~/dq�����f�MF���K�zLDSguS����i��%���������r�]kX��Z`c�x��$��ա��?"�� �t_���� q
���|�'�[V�����C��%��y5MH8�I*�4ӓ�}˸������q�9���	�=�nU�w>~4���{	7�c�^�N�e0���pߣ�ߋ�.x�kB��ʓ곔X�<���)U��w�Ht{\����ՈǻN��V�~��v�7:��z��Un����4�J;]h8�"Xc��]di�~u�%�Z)>��	c�m�((����Dh�5���-�<�v.ι�_:��$ߗ%���g(�9G���J9Be����bE�d������6���m��H��.�T*����"�O�R�������#vx!�TKq)�)��&)�q|�6U�X��s(���a��%��ǥ�@�r}�t�F��}L ���0�P��L^mpB#
�"'�γ��N҉k*��A>�U5?L��.<K���Y��L
�2�%���|��O?�~�_+�P�8�NnRQ��Ǆ8 ��;U v_D;zC~��i߯l(�G6p�\��~��|�2���{*���T�Zq�h��4�����q��
���zh����߉Ñ�<��=��UyX{�q=S��{nľ4���X�r^���n�Ad�TWӟ���4���/����8��9�����teld���F�R�V;Τ�?y@\�фT;���k�ͦN���������j��̙Kn&�>)h_X��n
4 ׿�q������������	`����y�Kl���*��2�j�J��: �茠f��R�&��fمk>����L�_Ɛ8��^��N5�X���خ
	쭺X�b.����Pv��#�mŐ�dQk8^!�^eQ $k�}P��Ph�0�Ϟg��ү5<����XIE䋶�+��ݨ��QyA��w�tc�ӊ!���\�}��Pk�O�#�9�#�OM���,���XڅIoߙ{�����8�h��IP��Ԋ�v\��P�s�l������� 5��aK/�wl�
�@���x�ѷ褈�vF�#��VK�S=��9W�����oº�����LZcL _�O�9��;�/J���q����Ӷ-d�w�4q�<�]���O
I�A��G�wH��G[B��8�^���Ɩ:[�H>��/��-����uս�ὮD���ꘕ3>9b��bPٸ�y�FL�x��u�C��T2�ok�d�&�E�]8��G>(jۘ���R9���U`K]g��o�D�Ҵ'K*3l�jt���A��%���읍S�׮�j�e��:�Q�u��o��U@p<��-�)�.�-.�e�,��_��Rdۢ�3 
<@rBDr����~4�D�67@����j�R��pR�Y_�1�J�o�2�}��2 �牦����X�o����5�3l�)�qFG~�9R$�5����Jh�3�CRxNZ28��?N:���t�F�T��>��6(�ؤ��t��q�bCฉ���B�x���1�ZWG��\o\�w.��ܲD`F8����ֈ�%��8�<���� ����B���Ba~��J��q�/Ȩ�M���ժ��957 ]��E���#�vM�F�v��6�V}zD�+k��dzKy���Zv�"��V^�師E���R�����cT�&O$�w��.<	�^&��?��o�0�I;u��DV����1���1�rEl6=Eſ�Gt,�ʔm#�)��"!��s�0�m:�?�A:e&�y�h�Wv��1��;� n�����W6��r��ms֊D���MUa�wj�]?�Hrj��Т�P99�N{�1�D�ѲH�����s�^$Y����ta��������G��^�IǲZ��5��_�<�-�+:2q�3�����"�M�3��b�L����H؎��K��VZ��Mnl+�ɔܦ}�
���	�y
��R���6��!i��1�)��a..5�*��@$���C�q�c7|A�h�N����\àw���E#V�}*a�~��H� �8ވjtUk|з~9�'�S�1��I�G&���ّ��pxq�c,CK,޾88&�v,���L�G�{��8�=����o�)q��g��8��MI�+��"������4�:F(��ϳ��)��0܀"��������K���^G�2�hI���D�^����x"�J�׃���V�@�'g�s#�����3��cQ��*�j��4�P[���	��\�\
@6��ؔ��rG
�ڝ���H�%W�z��}�����:}]��.�'���@ `"���H�[�ނ�5��9�> ��s�Õ� �ne�1��q���Y_�L�Y���en�,�{��R*>x�<���A��soT�s{�7�ڷ��)��d���Ru��>O�!{II��M{�|;Kej��݉Ҕ�RH��G���u"sg�ȣ�à��J��v�^�E��!?�|ۊT~C"��%�I��;����ՖA�?�G7���%+��~��z���ư[�Ѫ|?�4��k���X2��m����ퟨ���/,VZϸ˷j�5�ZF:#��l�����-�̰�v��<�|�����{�4<SF�m&�����&|����?4��Ԗ���$����+I�W��<��v�2'GԾ��p�0q����rN��K�� 0ds6,�S�T�@<*0�`���`��測�y���p��� �F�)C|%�a�PY�L��#	�u��w����y�!�����C�Zۢȁ4�*� y2����	h#���4�a\����鿷.��ҵz���@�4d�f�2P����T2�GZ3Ж�+��2��9f8\�F�j^tq3��~)2r��:��{�8��S]3挚wն��فے��Mm��(����G��`Ti��$�(��tw�!�eH|�M���O$c��͚LJ��׮��A+*�HkR���>(�ʤ}~O���B�	V����i���;~WJ9t��P�_��"��]R�z��{і��J���E^���y��~���W����O��\����'r
�3F�,Fﱐ<U��*����DwO���c"�x�>��A%8J_t����~u�g<�����8{�9ƐՄ�yIo���5�nh�\���D�-�l��ehwNe�K�X�\>ܱ����~+��,����w�m����^V.h�.�FN��U��3��Y��  �nU���[�	�IlT{��o63��kt��߆����Z�G�y�ӟ�cX�l�U�p�G}��,<�I��Z ��d����5L������ʋ��ݲ-I8�p�&�[��V��E:q�{ c�r����x����u��+0�V��:���zm�{v u��>� m�h����`�n�%���(�6P�:���j�����+,CN�τ�sf���Z?�� O�9མA�M8!��JD��.5lw�����R�#��䞦|"<9�LO�;��Ū�|Ex�~���i�Y�v� �h*b��^yE���{r%�6�r�"\�-��C�S8��6�P�ir����~�S`k����,����RyJ�v����P�(pR���k�65l�2�)�ĆJ�j��Of��1D'��]�<��\�[�N��_��s�����=�7�GR�"iW��{;y���r��V,D��,!���@���f�pR���j��D}�;�������c_Ѝ������K5]W��7�'��osa1�z� �H��M��]����#�^�K�;f}^���|�/vw�}�����Ŏ���\����;���D��DX�n&{����O��;}mU8G�e
�p�i��o�re�B�s�Q�I+�f)(c4R>��`�꟣y��#'��L��*��S�S���`�l�kMv'�x{?Y���g^.�9�"8��El�l�����p�꺜C���Ӻ������ac��%FY�z���	���)W�Ms��	øߏ�J�9uN��\��d�K���|^�nį�rڼ��������c�.p����:.=�"Q0�k�D�+���y��A�f�u8T�ϡ7��\gM&�X�_�K0Z<WY��	�㙱���t��35 Y(](I��S�KܛSEw=Z�"sL��>xhi�"~u+J��o8t82�r�*�m�h&W��[Qu���X�C��f���n�7Pa?V1�(
p�U'Hd�� ��HV��?'��m�t6����e�[17sH�h>�xs�3}g�	��{@�	��ޭ`�2b�����] T&�/CaF������=������"�/]Z���/�
	�C]��w@1 k+�L�I���)�̘�@EË�^��WS��棾 m�IA.��@o3xl��8cꖃ_��ob�D_���)I��s�0s��B�t�H�ۺ~�X��� �qH{	�\�@B��1�Mեe�H���I�=���lO��o1B���<��gq��U�NzN(���^��"��~��OhS��O�m@J5ќ}a�l3�DDϨ㫿Vj�w1�;���S��`��
Y��[�!�����iu�*m:�`��j!p��le����k�5�CVB�I�">�%旘����,���?�G�����Q�T-$�<���T��I�/꬘�h���E @TD��o�c�K��vaV5�]<8~$�Nն�H�r.��IxAɝ���s͊<�)V	�\r��r��B�*����P��IGF���*���=�4��^b��X�/�9�wQ\�{j��F}-�Eh7% L���FT@��e���>#��������eq�xsF,C�B���s�{Yg�d�ў$�l�*�@��i��&,p�<�˜ 1�;��{)�@k�w�c�-f�QA�����!|�A������gMs��s]��e�6��%����O��7J��v��_�\O�"��H\���ֻ���gw�-Md�����T�ոcm�rW��W� #�s�� �4�	�c�@վ����}U�Q���
�/!p^�E$"�����S[s"8bV}	��Չ>r��5�n��̿��>��nLV��`f+F^��y�?�(;h���l�L�F��־F���%�2�,����k����A�ˠmM� <� ٕ��R!l��� 
��!�� O՘{�O���鲋���"����QA2Vh��w�/(�)SC��� $m���|jA�Տ.�����$�Y���$�{Tx��b�ۭ��Od��B�Zf~%�Yʠ�E�v���Ahmo��T)'�EH����������cH�@~5�*����bHfB�:��KTlrw�n�>O�nt:�S�	\1����q&�<	B��횩����K���,�n)������]�(�&3���YE��Ս��X��h��T��ݿ[;�
�Ȗj�V�T�%+,�N�oxYT�d��G�&��4jJQ��n��Ҵ�ֳ8j|jiQ��X�ڄ���4T��k��\�ك��]pK�ZȲ���YI��ּ���r�������u����Cܖ����\������]��iu�i#x����b�Jͻ;�A���(��Di9C�)�p���sGyȴ?�$b[:�$p��ۇ$��B���Iɥ�s��n����{�y����2����1] ��=Qވ��)�]��esw�-�
0��
��;�w��wԶ�%��uJaR9��.�y�7���{!�e� c�^jsͬ}�6�����fTF�V:��U��E�6�E�.���H����=���g$��\έU�8T�(���8��F���M�lG�1ԡ5ΜL\��"���&��]Pu��AE
�C�t�sq=2�Ei������0G?-���Z��$�oԧSZg�7ba�a_I+g����t3'����;[�B�n��R�&�;��@�����%@��!�w��hZZfO���$���E�i���~���h�-��P2�!rt��.@�{MB���I(��%�VQ���]��f�"&�r�=����������������:�]�����̼o�0}����>	Ϫb�����nli
�in�0�d�{���gR����9T�-෶����xs*`�&�Y�+CC`��q�ٮe��)[N���r5��V0=���øo��q��Y����6���qng�[i�LO�)���h��+'�FPe������,�ͭM���}�,#�Xw`��"(Q%��kZD�^$����qݺa���=�ְ\���bÏ��T�C<���OS���q4L
�t���̣U+�.k������=�.Sr 泾�-Rl��H��tI�}g�h�2����CQ��Cn���WɤX[�w���9���&c���%�W�I��'撧l�,�i�M!��j�cר�uՇgH ��~�� 1������Y��U/��yX���R|o��D!�
�(Y	��T�-ؙr#:R�����W�L�1��i�u��P���/��9�����A�h{�u���Hv4�+�^ci&���`��Ѹ�K���iEkJ&\��� Khc�{"u]���� ��qI�IZUЌ����	\�G x�_؞3Sʴ�,�f��ό�����v�P6��X�3_� #���� ���њmWٱ>|ѰK���L�A��"$~y��5Ap���Uw?"�^UԨw'�?E�֤z���_��ȿE���X���х��9��X�ā�S��E�F^��@RԐ4�pC3��%��g@���x%��Kh��4��_���HzJn��K�b�]�����-��	E�l[�����L�w�.��	��[<Tہ�Mci 	����8����%c�^�R���Jyކ�;�7�*P��$�_Y���p����q"Bi��U����Ԥt��DeI�_���5$�W�b�a�?��#�xy���լ������b���3�(�@҂�l��8�g-�@T���{K%n5�h�#E?�Ͻz̺��9���mz<ت�� Q����&Ms�k���m����o$H��'�{�����à���˾��a�TnR��h�v���lc�`ڂ�~=�g�o�M.J�7�U��b�ڱ�gm�X��̒��n8~p4�>e����q�59ɗ+��J�^7�t&k�^ ��	O b��B��~���+ ʹ����Q�m~�"�J��QV�'ux�\6E�~��Ap�c��t�ӹ#n�
Q�+�J��F��K'���a�H��#OA�(v�FA��S���Sƪ:ʾ ���TO��AO��e��T.̣�+���ǣ�3��C��� I�Tٶ6��b�s�p�$��bU5[?��
�Nz�t-4&�[���Cu=��1��r�z��v[lG��r��b6ܥ��Us�_�?J��)��^��c �.�ŎHԍ�/�p�N^�F_G0��>B�p��'2��D�R�~1 *9^��V%���|l���;<�|�]����`��(qCse���#^��c���91qXI�z�!3k#��h���&D���Q�/ة^k+�~�	w���.m�t��B�gݕ0j�R�Rw2ט�4ҮKdU9К�	��^s0-��W`+l�֓
�A2͟�NO>g���:/�&�Q�u"�,���&�>�g�X��K#��)v���
|�8�FF��[Ռ�4�T���/dXy�K˝x�|�d�yi���'s�F�nv76]Y����_���-�3K�j`�xLL�O�����䬏�Yf*��� +�|NIx����� �56�ɖ=}~�p�l\� C��'҃s/���^Z�R�7�Z��:�v��������_R����<8�� ւ۸��4kja�ܷ��k�*��oUѠ�b�#����<���P�
�NM���h耉�[%�,حm���w��OV���\7.�
^��)�WA�Э)��2E����$
p�y�B]��d$D����>�(GQ�O� ��w��1�ؖb~U�/Y���g�Ծ�#W�Zf̟��iE�C�m:�D����M����	�0��ߨ��N�ڴ1�@&m�_22u�̗y>ۦ�^Ӿ#,ݦ�[C�z��A�\y��DT��;�O��Z��H����TN(o�Y5H]�8#�5>T�O�f<��}�$,�Z��`�~��#IMy>�,R$��u��]؞�����G0�7�'�����l;�@���A.�{���?��/�_], �DQI�PF�!�	39b2��QV�hq��;�Нe�?a6�%�C��4<�\_*�Ic��+tҽ�:9�Z1�j��z��h��ƾ
��6_d
^�z��kU�͌D�R�rQ�HP��w��c�ԕr�IH�g�z���daNb�R��CohI�iZ�UA�AS�k�:�h5��(��!Ϸ9�P�S1ѽ��/qt~�`IB`���,k������pؠ(0S��er;��b
�y6�l�-) a���]����i�5�(��<r���Uz���,*$P��$����pl�mb�2��?�n�Z&ʀF@Wv�h7mݯV��C�3������a���L�Y�W�b�y��%��풶��DUi��B�0.����;�����u��10p�'�ަ"!���C՚R�Vm}���l�� vA����t��2�/�D-��&�푙���4����C�c[��E�!��Zk/�5
Q�;�z���o����J�Dw�Z�����b�~������0k��*>�*����F��3?y�A��ԋ+�w��&�n7ʂ~�g$l=zhaf+ {�o]c݇�i}[��浍��@Vy%����F�
�Q�1Ǭ@����#@)9��DF��ʬcT��87V*��%�	?� <u������C_ǁVY�Gc�	f­��׀�JJb�~�d˘���Æ�w�(��m���9/�0����W���Ù��ʉp��%�&Ք�1��+Fꦍ ���#$!g�g�m���k@�"�cR��>��H��S8	m".�E��!��į��C�ގm6��:a�*�Ą���/�7�h��kE��Ą^mv���u6�!������Ȁ�^�2͡{��ʂ��|<�]���U]b�?�õ�;�̩�*�ߑ��9�~+Q�1k��y0�s�~�)�\������1��`�����\�/��:��T^1%	��!O���	��Ƕ��1k1[�Vb,`"���y�~lԨE��b�C��� ��+��I��u����7_�@H�`c�l������be��`%c�~2�;4vG4�Jp�����1��e	�f�4�GFtO��ķ�I��g��@�& 	�x��h�|`f�
�4�F��J�{W����x�W4��O���w ��*�%ȇ۸�\V̲��ȳ�!x����0�1��U�U�#���C����w�y�jB�kV��'/F���X����SR�gW]\&灄�<��^�.Ud0k�'���mANH���Mk���&&t��?F�hSn^�ܚC�bZ��xٰ6�����=D�k��ƥ�f��&��b�o蛤��z�i�$f0d^��@S!��{M#�dl��!5Je�̕�~�3I���J'�-����*Jw��$������ߏ�h�[֜A�(����͂����_���8 �I�J���Fc�G���+�t�l�S����9�9E�9C��ӌ<q㒝����y�	��j^�q�,�/FgP��6f�;V�OЏ��<0�Ɩp=5:j@+7�\�d_M�tB��F��@�.�H�D���jWsu�{�D���y��Bo�B޹'����-���}T��f�b���[ݽ%s>3[K������?mQZZ�&�Ɯ���4�� ����H���̲���a�����d[�iޖ�]݆�e��*���9§�m����M��:�<� �u$j���9;�_>f�jofG�uƃpϘ�'��,�-��n�YE��윉C�t�A5Q�)�F���f�9Z�ST`[�/�����`�"W�r��dp���Qx1�vJG´�
�5��)	�<R�J� !,�6�ڕ��'z6�a� ��OK��pd��7e�!�2u�@�1�}P~��iP���!Azن���A꼗�.��p.Hbp:���}Р��c��S�`��J���.�֐��K�j��� 2�'%x��j?�W��{ԑ	�K�Q&S'��+u�2����9��M�J���שׁ�t�������O;� >ÛM�Z�ߩ�z��*��1�S9;;X1�Y����K+P{]���em;��Pt.d�5��1������� �����74<��*H���	���vi���q��a����d}^�S�,���W7�Ԁ�3��O�Y��~�æ˨�ې@)��B�|u�Ɯ�c7�N��O�x_Ǒ�-�(�/:&�?\���U�bTu@�����A�V1�uf�h�wf6��3%���m�b�[/��f� ��r�8򐶽
�J����g������"���;�<.�z���{�N�\�r�`"%Dª�(A�`��,J��(��h��GD�+G��z�̎ŝ�G��#�S �^0��݈N3	�Fu��|��L�TA��k"�\�E��GkUJ=cXj�ե�`&U�U�x��)(Щ<�p��(s�Э��)Kdԍ=t2�Ym;��C��Q�8��ӈMʜ�+���P��e��sg�&��&��)8z0�ͳ,)���sh&׻r|�`�@�p�g��c�T�<��W��������O��$��.��e����wZ-��D�j�W��b>�g��M��3��fZ���4�M��]�x>ކ�_<U��~�o����>�(]�4�/4�FD&��{%pl���X>�&�ސk�
:�8�&
�5��~z��鎻���r)r�ʅ��^*���:`�C��[&e����"T�hpQ��Lg�
}tw+��vUa�Pa4>)�(��W3'%�刁l��4@� �����}՜�#���}r�#?��	����B�N��N
��-���Ky:Ӝ=0&���FT�jqos)bb�����FNN��:�V�PO�#0��J73, �3�Ŭ���P܁�̮��d��(zI����>�7ʸ��aHu.��J���h��z�_�zsPl�Vξl�0����7��ǵӑ�a��R�$��v'πVH��	�4�\,4%���ڝ��J���$7�b/�G閜��l*Լ�}����"����r,[�+UpE&Ok���N�H='�+��1��ß��-�����G'OR���^F���)���7L���^}��ô�n�bh%d]���KS>`�4mݾ1���?du�C��t"��qR3iK8!�w Q��X?Sxd���}"`ת�7Xt'�;��üٕ͘vj��#R,c��ʃD���hks�`�;�iZ#F35s�%�烞�z��o���dv�;������5tS@�ȿ̏p��!My��Tl����ͳ^�v�9��vM������ ?�U �-S7 o�	�qk��?���lx2��g��Z���هd��ө�j�,1�J�F�0�j8�^�3��dj���t�>l�J|�M�IY 
(�룫�_�N�S�,���_T2e	X�ѵ���T����ۼ+2�z��d�w*I�t��F��Q��)�g��k��H����`n�Pl����1؅=���p+�Kt�F*@��w��}##p,�?�Հo�E@�r�J�;��o,�N+�G|�v����ȅ��S����q����m�� ��lމ��@�?p>�J�k*st.��e%}�`�iX�E�?�[0�'�ɷ%��X�.�5��4�1]����qN*���i��	ʢy,�\��#g8��g��f�$η?�K[-f�Z�v)1��F�cZ�*M���b�Q#K����}��5����� �v��y)>S�r\�HkTN6[6�&w��+�MYC��D�.2��z��P��	<���h�[u�lY�
%�1�(��˳�S�Fǫ������!��~w�#��Hnp.R��% eC�D��
�Ƨ����_2��u8�����q�_���x��&n����v�=��jx%7}V�t�UIM���1,�Ñk�푛l���0���W̼�uw:��[m��3���2\|�ɨ�;|�و�Ws{����)=��H��2c��5�A��`���Ñ#F������L�:��)C.��|$-t
��'��p����>��^*�������A���25�raä!(��������|-��Q	��=��F�Bw(�+W9�́SЖLt�ӠJ�̩���[G�����ϋ�h'J$Ij�MT`Da7��ȗ}�q��q�G!/|�9 ӝ��`���DL��9���"æj>�O	�x�f�(��UkLu*��𵫤�	�I���4x��|����bK_���N{B�l?�6/mN�����������]�Z�@?��]��5��o��$����9�@�l��Pm4�R����8�Cpu?�.���{�)�oƯL�B1�+f%�<����S�n��/Z�le���db"���zk�`��C�m���؃R&S�H��z[�/�\|��ix��-����d7;�C7��i�혣�lA)����ɵ�n:��a2�A{��S#4�������4��q@&��rBI�U2@6(���B���NJ�F�%_���ǝ��}	�LH��i|����_pj�Ӳv�#�v���`�	"���T�"��lZf�x ��S1Ժ��o�m���.��*�nόqz�UqAL������icFFde)腽�2�t����zW�j�p�
C����j�ҳ����m\TB�' =�С@:��`�'x:�%�����S� ���x��j�R3���c�����8g�m�������3��P�D����B~I� N��2�D�yQ�+ B�J����w��]oELл���
1*���a<@S!�G7�]M�c{n+J�j��J����V=���j�d�F:�����B���n:dĮ�^�v(7"��7F�����.�-xVG(B�/�h �E��:���� ��HZ/��Jh�;�&p�R�>��.���Af�t�����Y�0�y�m|R�D�}:��qgV�u!{匉+"�Q���ٯ�j�5�4�k`*&���1��iڣ����f,L�b���#Ul�鼮�޹����K8��`��+CX��U˫����O�ˏ��=�1� �t9�������}��)z��M-�w�}1�Y�
�����I	��~�1�	�m�
S�N� ��T��+����O��ri����Am�(�/���Vi{E��\RՉG���P����=ZF���8�H��Bq��~�E9@����Z3�Z�jH���ǘ���Y)z�s��y�!}�T�0Mn� -�����)��ߺ���nY�/5K|U������'���U冁�A	�r`xN�r.� ǀϜq,�a"#�W�$^63]ûl��1��1$��.������[�Mp���W��],0��&�����q+E���e=�+�Ja���D�z�Tͪ���n�)k�Z��fD����H"[�[����k�G��uW���N��i�ߚ����|����R�H+��S���S�NS��L�b+�eS��'>C&V�Qk��_w�T��o�z���b�p�*x^��n)ku�s?L�M���\!�o �����T�=���P;9���� a�+�z���b4��,j��qṓTW�"���u�
���8�d�^ʦ��OR��0�d��:ً��X��Ϯ�&~|��I�?����v�e�����
��EU��/�Z^u
{x.~��� �BC!�`%MK�-���S�.�� o�i��� ��H��_k�%��~S�́F��JZ)rY�_%�x�R6�"����e3b�Q;�2��^`�4
霐��u����Uģ{�������"�C���|٬�3�20�?X���m��a)k(&�c�����ȍ�:.4� �I����C���(�Q)�{8-�խ1�;a4���c��5��aH��6��6u���0�i���k
��.��h�d֊��݅���R�S0Yva�{�Ԩ_t.�����g% G��K��b99��]�{AD������}�G�NA��@1(\����Q���h��c8>
��]�f��B1�f��� KOU���#\��U�/��yAӛ��>��_��70�r��u�5��y�z�B�o�eJ�C`n�����LG4׹"dz�s�����Uþ@���r�`i>ـk�(���ͯr�fl�ݬ��&��ň9�$_r/Lk��^��T�,%�31�8��:m�pGIsF/lv���s{r~�"�Mq49�;��B6^���kv�xcZ{�`!�6CZ
	Y_�}�����]�J�1�H&7����0@+�e��Y��߬���"m6|f�=�@���~N%�>��T��AY��8�#`ǧ<�c��/8�0-<�sF��o����=m���1t'+���;۾	������1U���w��s�Y�m5jS1}h~������4;�W\�ē����T/�G�_\P[�7m�\U�_�;��e%����;?���*SE�������'���C(f���+]Y� KIKҀl
߉�2�������=�����+�o���T�
Iݻ H�9L�u
'��d�"E��tM�w*�9��� 3�/�%����0g���%�� ą�:���Oҩa���8�{
C���3(�����s&�c���/��������U����Lv��P��\n���v����!%��A�_���2^�4�Ym<!���V�>�����1���7�iʇ�7��F��8���9��µ���Q��{~�~�ވ#"�j�b�4�����$N���͆�3d~�h���
������r�c,�v@M3l��p��5k�\O�2�7-S�R�{�[	��bD2����$��wI���ΰ4'$�o���5��!�ѫ��ݺ�u�א<�4�|��OZ//�������tK��9m@E�r�o�"��6���7D]��J���c&���iTi��1r�2XN-p�l��JU����z� 2ǀx�o��;�)�q�b�C����p-����*�|3L��;�[�ڥ^��e�h�Ɇ�v�V��Q��~3�r��ɇ ŕ�;6ኧ�F�L����|�����4���gfyQ:����Cƌ��E������@�!���/p�6�[l�S�lӺ�I�*��
7de�m�����x�ޘ9`FhQ�b�I� <���G��>}���m��t�Ð��႙DZ�i��l5�hH�f�d��g�p�G&�$�f�T��k���`�O�����r|����ӓ�o�ir��OJO*g�����3@�@��Xa�O^f;������o�n�*�R�� 7����j�/6��"f9��^��#���K��l�zg�T-�O�$4��g��ڔ�>�c)*P>?y#��J	[���ϷK��/��y��t��0IX7��CC�O� �;�h��ye�Y�e�"�چx$�t�gѶ	�S�kj�ZK�t���[���?IH��A�Zo�hg)1��y���>@O���	����ބ��f�����XA�l�!ѻSg^� dI>�6�u+��<��[�w�^�W>�����N@Em�t���I������!�t#wb?`�; ���_p�c�tƚ�� 8�w�&0
�]��&}��a�0����/?�Q��x=��G56e��n�M��-�����ΔB�-�8�N�{��t��2�t쾋d�C��۾�9"P.��6���K�̼z�+.C�P�8F�b���t����ȍK/LX&z1��L�w�Z�6�d�7�.u�CY�+��]r3��p-�cmV���8�H��%ܷJ�
9��(7����ѝp�	��N�קR^�ɗ� ��3QqQ��t͙�m��t=�a/�-A���
7}�ɰ�,@[>'�.�Xq�AΏ?G��)Gz:�n4>Aex3�֠m���u"�xފ������n>���jg����*�|6K�(�r��h_/����<����K�˾D������.�cU@a`^�@Y�b3j��P��s�y7"�P$]ysB|��ώ �m�:��U� D%�t����N�)�sJ�z��l�]��?�G�/lwj�@xw�L��1� |�IZ�yp��"��o���%��Y�;��,�w�cV�)G/� t������<|0N��|S)��%&@q�X텓�Ե{��|'�:��w0�V!���=x=KI2z},��`#r�|���i�U�v [��y�JĢ|��z��
w��c�j��r��8*����ۓ��>9܈'��#EN�t��:u9e !6!p�9�G�2��2��˝7������G�������Y7�њZ@��ϔ�>����@a�p6ھ�.E�"�,���˘s�s:3$$m��v)E��_�=N�fa��<�~�'L�׋���B_Q(�O- ü�D6���]3��'=LcZ�37" B"�@A�Ц�*�Y��,ȫLhDT������'b���\\�Ͼd�s���S��6���uE)؈�EJv�O?�Q��1i2��%�:��9�~6��#�24���*$	�!�Y�����a�g�ѓ��Y�}�#"2P�_��3�/��mp��8NPi�n�����0>�?��Ƹ���v`:-Ӝb:�b'�$R}L�lIAe1Wl���'^����Tn�~��I�p�!$Zƚ(NW�h����suPm$�%/AĤ�i��Ń.��=�yZ���яZ�, 
�����@�~2�����]:��l����q��E�)���FߣɴN�)����BNHy�%��`���)5�WI�OS����H9}�"��ķ �pM~]� 1#��g��E�ŧ4�Xdg
&���?�ٻV���h�&�>�8� b\��"�3 ���;�Wi.��͸m6ы>��0k�x9O2�[�܁ӏ�|-^+a%QBj��:��(�c|� ���{3(ŷ��_Q�-�W���ƒj�C2sz@�
�]���D��9�C��͖��!Pŝd͎��7���g ����G��Íi;E�K5e�G�;s��$X���t�c���ƼLg��<�Ʈi�E�&�rD5I�����nX�Tѐ.�#��%HD����P�g'�d򰭰`�V����!�w
�[FAZ��>.r"��u���(��vO퓻؉c�x ����`.z�&B�ϋ����ꏁ���j�yY���M����gi�V! �p��uu��6,|�-�F+l=}���([�f�k{pS����Y��X�]�>�C�@7�娞1r54?�Ш��-�(�S9mSqY��QX��Tb�-�"�c�w�Q�͌F`�>��l]���i�t$x�-PQ�F2v7���Ѻ�d���%�zM6"޸�L���J�>J:�2J!\ \e`�$i�¢A+\�a�������5��(�m+w��9�^�z�f��$��x�bԸ�(��]��ϧ3�5n/����cd^I�����F���i��M�T"5�²�!h��wˏZPk�:|��Z1���-VVn%��I�n�iW��I �(2<0��`h^N�ҵ j�d���mף����-$�Bp:T��Ǳ��L{ş�a��u����<���ʖ���G(��A�̃���(`SN���q���	���1�]��o�#L��� �����l�g�W��+��BJU=���x$� �3ء%s����Qڍ�*1X,��~�,B����j���<:�j��0��V9���|S6��Q0}N�$3��Mp�2����z�޼4Iǯ�2��v_�l����1�>P�t�y�8c��(�� z�ֆ����p��O�i.�~�y�r�W�%�8��A�l�̩������H<�뽳���})�]�.w�;X-�|�Z�V^�:v�?o�z��?��I�.c� z|��8�F"�]B��9�6� D�
[��؟��މ����D����ڕ�i3�5�ɮ��]�"���A�^f��AZ��2oL��b9���l��ʛRI��V�y"����ȓC��C����n���٦�	oԠ��_�%S�2������3X�� 9ȵf�%�`��wZE2��K$ŀ���Ĭn����yh���h�x�l�;�f||� ��lƘ˚$��y���(���4�l�q�Δ��j�¼c�.�KK_!�������^�0�{�m������͟֠�<��ᡰ�U���baF���m�5��wH7_pEJ2�v�Z����N����`l�Z���b{�A�%�Pk���ݑ�o��g^���#��PYݵ�D�5���{�Y]❚ŧ�q���P�3(�17�t�L<*I�xZ�oR�:�]v`��@Lr��#><�?/mX�ٮ�Px�]�ǕIP��T�� K+��A2kY�"�� n.z�9��!H�)y
|�=�y_a�mn��^�4%�'�*�t-�aM�Znn�`'$@c�Ĥܯ�ψ�{���_��q���gΗv� ��8��hǃt\+���& Qc?x��c�|N� �>��P]�o|�Ő��l;�|X6I��E��'bK&�zhJ�ά��v�����mhU��h��:�Կ�k����-�C��:���Ľ�4d)<^�C�V� ���[����޸�d�rgr:��~>�uz�^-�R�^�7����q�-ǽ �k�4�s�%�c��'�e�*��I�~x���96iZ�ޫS�է����h����o:@�?f���r5r���<�R�����ڃ=S�x�a� Ў"|��]���	�9���p� M�B�����QW���ˎ��x�N�_��l�j�D����~(?��2@��6�+�q��}M�x����H�[�L2:��Ѹ� ׽�
F������DxJ��8�ԑ�S�˕=��;_���Z��i�^��R�{Zx�C�ue%ܭV6���(�ɺ�`{-6�:�.���*?�d*D�q�������w�b\)o2�\���)�X��^�'�5���*_<���*	[�5��M��/>e���v�,�ç~��;�4�؛P��`�2�����/ǏS��Uuy��w-�%$���#��V&*��Թ�v7��Q�[-q>7�u�
�G�3t�)��qCf���� }c��-t�7����,ݙ�0��Y��%���gh�0�q�;|�b��.#H}���px�#��v�����LJ+��*�S<E\sw���_VHD/'�IsS�y%nUOg���� G_�=���ox�_܍��{�O�k�c,�U��U��n��7SC�υ�?x���@�|��.��;���<�d����Ή�� {660(e�����{��E5;<Ox"5O6D�]�#�n���u�*֭;J�ExZ�{rb&��]	���"�]E0$��R��&a�ھ4|��0#G���x:&���C���g�i	�zN�k�+	��8-���Y&9��I�M^��S�{�KWr0��dN����0�zN׺U[cԔ��D�A���T�E�\POf>�P�_h2t��D�z&�V�DN �y�.^lPK7�����p�x��L�|�}=�(U��Y���zG����������^�������Z���i�4~�ۂ}?�M�!:�ޟ��Z<��}g4�g��si|*��[�	k��I���P��ߓ�­�#=�z�ZC!��8�'���Av��zJY�^@�BUv5�[Bk'��<<r�s���52��W�3�0�r�j�j9t�_�I���z�Qpl���Υ\�����v�b���j����]Qsj��L�5��{�Wc����C���eo9���|�Ƥ(�:85��X�i����TSǟݸ�Q?�[���r�~��x�ֺX�u
�g 8�b�.�	�M6$(��[O�<�����X����^Dha�e��:P���!Ӌ�ϰ�u�R�DG�7E�n�k�RLk��lFm�r����&)`��G��i4�	�G��tZ�C0��~-F�>�/�D�?�iY��z���kA���d�3��x7��.�#��C��V~>JqЛ΍ r���4��� 
�55���f�7����R��S�U`�;��l�g
8���{@�R?�&�7@Q��B.t�!�ƻ"��e7Y�?�H�Dt �&�:�~t��x��#
ND5�`B������3&��7��(��F��z����0�U� ��A�/����??+ۥ^��{�ro:�I4��?�kK�����~�b�bSY��H�s��Eۭ��;������U�qdty,bD{*��%��I��� R�Ln��]~$5��Ed� ۦ�.���ߧ]�_~J�p�&#3A�;c҄ɹ"E���޾y�~�����6y��P	:�Bg��
�
i�(�u9�O�G�s�
#�ů9\�-ĤHN�)>a�M��� j]���H��ƌ�,+�s��61���W�Ü�M�#'s��R��p��o[nv\�W�8�1�gT�����Q :_dn�'��~o�*ַڞ�p��ޛd��`)]<�c��&��zǝ�6j6��L��F��C�A�*�Oh���ER$K��ˢ (Ƌ�~�U�kkd	�V3gU?�q�����ګ����R-�P�����ם�i�4'�ݒlK�����s�ۃ�I7C�QN���	�͈� ,)��CJA~�#�$�e��HZ�f��I�l�cS7v7�w�ٕ>�#Dc���ET�/����W֯��u
�L�j��T1{-���~�K� �!3��U�Ona�[F�Gh�F�ih*�Xc��I�I����6�����0�C�X9d�U:���dX�j���{�3���B!H|�Ǐ��8ڴ����U�J➂����p��,�b��sF-bTq��'R!�)4��ױ��2���F���(��Đ���T�xk��^�c��d�r�s����缽����Φ�@�����94�^	��l�� �TG巺+�6�,1�cm)�g_���q�V�W�|T���/OP����yJšb*`�Z��s��D��6ľ3�eq�� `���ᆞS���S^A���a��U�\�v�2!�����ϑ�.���زzC^p�J�#}ӕr��@�V�Qf[��藁��q��d�%()%��"�#��i,�X`�C��Ez2����c��� �!1񀇆m��')�=��?�J2k�6��bh���{�/u="���/��
w�"�#�d�"��ą!·P��� ����BҠ����Cr���?++�J&��/)!�!ݍQ�w���"i���#���H�5��� ��� Hy)Rf����·cNPWDc;uA�JE��K>���D6"Xۈ'%s2i;*U�r�����8�K:���Ȧ_�{ӏ�E=<����	��P�Ӕ;��Th���iԗygԩ*�~�������������[��\|�B��t_��dk8.t�L�O������dnZ����GrG�Ր�m��t�@�윤�p.W7{wk)d�5F|���ȗ �n;�)܊�q�dW�X�˥�ت\v(�����ߡ��0�'�{~Y� L���N�k����?�#��fݐ`�3#�����lR�N)��(�K�eCRэQ���ON�S.k��"�7���b-�˼��4#�ʣC�OV�5j��bM��R ��G�S�,�6Ck��m _p� �|$��~W4��G��q��zV��}g�����C�swg�Y�IX���Ps�`�&�����
�(#�u��=���n[%�X�!G 
��;��UAO�N������=Ut&m�� ~��ZNG�ז[P`k&��W}�L˒���CѱE0����v�����V.mt}���X�5���6���Z��t�EM�qI 5Ť��+�]oz��v}�����v\]��B�7C�P�c'�4np�Ƌ������;�0���Gmͺ�~�s�,Fb|k�K;Z]7aA�(�6�9�d�⹎$�H�I	�}إ4���c�ε_D�=��J`�����k:C\��0�s
������D٥)b(#����WǙ�Fe�u�[�v�O�2����yS�V�0���"v�� ����Q���b�H�Y�5r��w� �y.
��&����nsH�*+ӏnH:�H�=�Q�7�*b���:�9=v�&��Y)l-"�w��ڟto.��r�T(nФ���p�8i(�(���-#��`jZ)�r=C�޵�ip������E|��l�#Pbp��%3_��+�7w��l� '�t������F%V���7��9�~G(�@"��L�~��V�OU9�eVЇ��������>�����	�1i�@A:�B��)�i'Pc��ƪ�ry�ՇD2%���a��� ������8ŧ��r*�m��T!2�����w����`��G\ۜ�)$ׄ<�k��ň ��I���)��׽�,$��^֫ ��ds�^;��9ַq2��@�d�E���(|_hdx��L����^�%i�{�����lx}�U4B�GAd������o�0>�X���,ߕ?4°��|�36��a/�;�9;B�ED�&m��S����_R����n�%Q�&��}[���l�Q/k�d^5�}+6;�S�~!���/A&4�EF�5�7)J����Ƃ.��SE���Ax*�W�2��8A4}u43+(kd:�������}::�t�R���]�6�qm���E9���"峏��fS)D�Ã�x4�v{΢3��@�kix=�� \� ���<%�#Z� ���u� �T���yt�6#� n�H�MH�>g�+
\�k��V�.D%�7MOC�f]H��E���u R��6gW�s�N<��jZ�F�d��q����hu��Zhn?C7��� l�7�u��@8g��(֨��.	F]s)Y԰�I���'��`�Z�ܧ�M�G]	-�r�k���T^:�X��I8WRS���.��6���.�</�lgaV&wLh�V�[��Q��pLmK�H"���zK��� K�qc�����1�2T��Zw̊��.������� ��vW@�70ǂ��"�W����}�R�EK�}�(�5��Qu��`���C��,�/�pDc���k����m�Ju��
u"?��@��;�m�y��l'�wR_�7bp���C;��6A�J���4���
��/��UV#���i���d��^E��`ڵ5�聼��A��#�^�e"�l5?�iԨ-uU���]"��F]6'�,!�	��5� ^�k���roN���X��$Ӛ˪C�s���B�U�MX7���SWf�궢�m�Q^y����C���6x��x 3�_;�Au@���Dt����Ls�	��O��D�sK�����S�6�����4�1]����X��yUWR�kMj�/E��p�+�b[�ПI�*
$�=��pȭX�啷���u|G����{�p|�"(�;u�!�,�y�)&o����]��F�``Ÿ:e#Gsț�[�L
�S��I,_S���� �PTLN~�OcTTƍ�nM)7�RV���b'���":�Yq@���H�%0�C�T����{�O�6�R�� ����3�o9���i*è�Yc���ڤm�.k�'ޱ��65U�O��O$Z~�|iKj�"w�,ǳ��:�g6��X�c͟u�`�q���\�kH���~�D�՗]���:�^�~�/�c��S%ϱ�'��er[��勶��)^�֕��y�Y麍�h�˖����9nMW�����w���/	3Z�-�6ϝ?�pֆ�⏰���wޣ�U�ȃ�~Xm�-���l�z����u��U�P� �<�۔�1Я���T��w?x�ۓ8>0b�x�Y�?Q;������%'��k����νɍ��lDM-�I�Ғ� �1EX��x������I��ïRA�f�X�����C��s�w9Dz ��HW�I�R\eP�ן���v)��~�ˌZ�n�cx� }�lh�	�����I���0�bq����8CP�9Z�k
��	�;�A�AU�'��6=Fnۏ��2���˶"�s�˻v�"vk��]�����.��Ao���~�Rs͍�%C��]B��q�-�$->M�(�>2�v�ǌ\��gn�x�&j�-�#��z h:w�u/�A��<.��t�����P�_d�UvY�ݳ����+���)�9�k�5��G�,��le�/���7���B��6����O���*��&�n�ް�TM�����nw�Ȅ�@�r03�1koU�{	(����I�XZĴS%2��^Z��f��,;԰X���'��lf��1y���Uy�Y�Y^�&��hi��_��O�:ޡ�m"�|d3���+ǖ
�ɑ��"s�H�
�K!�t�6�*�n�'�c稢9(fqw��U�ic���b̴�Ǻ~������S&���^��\�[�����sg,��\������F��uDY�߾�ER'ya=�Q���D��}�X<Q��l�~D$z�˝G^�+8Δ��t�|ݬ���ȋ_zH��  a����N9���$?����e�F���Ш�8�
}@5�p΂�glag^jL�@%w���!f|(���GE��E�ֺW�@B��������v��D8b�ph�R6<�h�X��m$�R��|��D�o�eהj1--	��&[�Y�lǹ!~�ƿ)�����7�*B�L�h�ۿw�srnv9yD���1�9��*�L��͊�a�(1ee6
�$������p`f�A�F�P�ƀ�F�k�$��N�]�~A3P�H-#ށ�b���P�
%lRCy�=()!�^��
|�^�_��� �����K1��h@�����-t�V�of�u�wt��۫ךC)��Y��+ ��# ab�j�}w)���q��T��:x/�,�꘠�j�Xu�E�q��k�C#bI�^˓��Gc�Kq��u��.OTɹ0�h>���4���C��b������Z�*������~�!����_젶��X�O�J/�����ܟ=
������>ޔ怨����S��U��~M�y���8zo�Ad$�K�AHp_H��g���p�b�;���1�L�Z��'�Q�}��!S�(n�K�i�SH;-|�B;=D0fOJX�}R��k��I��1�o�C�lo r.����Y	]��3�B$�����\{�w�9@��^o��L�b�6�xgy��v�gy[�s����ip�ص�yA����X��Ưn�4G
`�q9*��y%ڇ��WMNM����}24����iu� a��	�� )�����O�֏�[����u��R(��B�xZ���}o�+�i/���l��F��T�.�f�v=}��}�`"_���Kf���w?gz���4�gocȉD����i]�҄#G���.G�b��W����[����I�Yצ����p�ilW�X�ޚ�b"+�-E#{>p��p�qG��z�Ebt�J~r���a�˔�ï0�`�"�-�w��q�=}p�狗q�8�"�0�������ki���x0�;�8BDNĴO��)�?�Ų�9��~
8����w��iR��-�n�c,ȟ�hƻ��lT��X���kZy�G��Ŧs���g�	��8�Pݢ�x��1)���^?1��B�Ģ�;|����B�)q���#��i/�2a=I0w��Hg
����N1�4e�aIs������������mH�"p�GU�K��o۟�U�X<���כ]��3�*K��q�ۻ���ݪ.��A��s�&�l�D�_p�·��-�w��cձ����(�Iؔ���a�n!��98u�E�k0�ې������������f(|�֧ �ɝ���@�'���Ji��F��^��@��@����L�*�GYE\�0�0,GSO�P=:��Ge7	_��|4ro2a%�$�u�!Z�W�P�'vh�A�"P�	��<Ss��d�������Ki:�������U^G��K��$^�B���d�M���ÿ���#hl���r���E�>�$D��W"��bM�AXn|b��̶4����_?H�vh6+�j�%�r���
^��m��e�/R��oڵ��4L4%��a�����K�'���?���0�2���jYy%iΠ��[)P4�:_I�P7��03�p���y�I��5�$G�b��.:҅D�ҷ�$Bem�SV�_�<�������%�z��f����t�-�m�^��_�� &��,	�CG�Ĉ��X���I�HTOE��;�:0ܿZ_�P]ȋr烎x� �:Ľ�?��W��<U�qk��¶A���^���^!h�m$�gm�V�{�w����z{����.h�`��!*O��*����� �5y�Yx�Hc���kLղ�Q�^��?�O�����E[����)8�	�V���a^3�I^��~�t����0���5�tU�Q�Ye-��S-G�,�u��5�`(oz������i��X�+9��=]�Y�z,�E�c8��l�Z�C��8U��<��r��i
"���	�(>=	�xZ���I��T)���I$R�E�7�'� ��2.��y3^H�����E	$ԗ�)�$Xd�l��@����q��T��C)s�٫�m#��q�M�٬p}��Z��TH�3��υkH�6�Z. l&j��ح���8��+��%���KE�ʸ�봑YAa:c���byk�x%Y7�6O�:��I�:������+���w�'̙�����gc��.�8�Ȕ��	Peݾ����p��$�p�)z&1���K
Uș��c��ĐL�ZL�*� ��nZ��#U���XB��=���[�#�B7o�\��7%�D<,�2��6��n5b����m�o5����W8S�}��$6eJg�}�����jw�V�p���Xv��)�\��TQ�6��|E���]s��0+�M{���Z��L�(�k5h|+<\T�yu��,�<S��j��+1��Iy��U�of�zp�!�ꓳH :�(�b�Y�:�Z�W��Ý���9mi�_��2�G��5�ە���<"�\�����
k3Dt8j�tNy0�c�]��_'���ҧ�" �D�1�Q��1�o�cl7��~3٣�F���2��Fy&"���v lͬ��(��� ��Ao����e��3��u���|����o1rkh?��){�NX�|�ԡ���"w�����l%a�)ah a'4K$.��UW�aܒe�gqe/߳���Zq�V���;�*��\���^!Y��%v�fО�ˢ�Z��oݺX�*��o�ɏ1Pl�잔�F�Ɛ�mD/5�+��߇���?LJ�Zw6�A����zC��VS�ú�2��&��QLCbMD���G��g��?.{�v�HP�j�w
���"�(�,��g�S�7�Ω�%��H	���A���er&�9�+���*b�t&�pX��p˖⥣�x�3n!��CMF>p��7��s�ϫ,ϑ���*��} �P�o]67�9zX�VਨF��)��X���մ�>Ez�y�(�"D�x;��m��J����衡�C��$N ��1Ώ�ɒ�~<sc�3�"}d���K3��K�w�jAY��s�9yV��%�œ�����Snۑk��xI���.X�^g7�f1(u�� eEӆT"z���e�e,'窙�B�d(�ʘ��߶zLe��u��T�ө�0g�����d���"�ژ�{�'F����
-?�%+zҊ�7����B� �q�Y�L�@��*Y�Y;
5ц�@��|��б%Ǔ~�����G?�6��Lq,9� #�	W�-:Ε���M��i����J&�<��� C"�pш5̠��P�P����7{��Q/��\�c�H�u1��d6�l8�����V���Ň7������˄�VC�J�D!Hܳ0�4�K�D4��ݺ�NT�'jwR���}P&RZG�t���=��[H�Xv�Yrt���`o�g|8s�9r�d|N�p6��"
��ިi���ч�>'���`�+�Ez���C��/�y(J����tȻ��cz�'���a����M��A��Wcm�+=R�}UJe�<��$�O�L��C��vR��[���9ي5��u�������������!��������H��J�2����C�M�[�ןX��i��9�٫�H���n��g�=�i*�x�`�pq��F{����K:�`��	��ߖ('����6,�IHl��r\��d�t��]*�����%�ϸ<jy*�z�Z��'��*E���3P�r�ϧ9�3PT[�oO�W�qnx�����P4����n��IL�/�T-��x���O�8뇘�n��<��ѯ9΄XB��k��!�d/�X�O=���1X�j���x�"���mw뺘 J����#�o�qV�/N��%��6�r_��Z�ŀ��9���BO�:cW�����G�`��9����.�3};�"������Ke�HYt��4��a{P�zUm��e�"�!q똄�W�Y����ז�`f���@�`3�~��ׄvS��dr�.����J���.��DY0���]�YE�J�F@�Uv\x{�=����A� ����}���>�w(t�ZH%����i3��MA���";���l�Z3ݵT�bbb�i�H�*�m>49#����!�pl>���P���}i�Ҫ��/3��]����O:ʰD�m�,����d�� 3��ӓ�<�w��IN�f����"��o$
���`q���C�ћ*�j����p�}���
(�͟�D�h�MD���,%h�!���11�T�յ�b�3.�..���\4AC�H���"׭�YT�&�������o��9�]/�"�����T���$'��x���5l��y�[�O-���A��9~�x�?> x&D[���+<3���y� u�*�߻�%�:���TLR�\��+����v���s���a4ՋU'	vY�B�)ni��6�"�!_�í� s]l)�~�s�B�6��d�Ɣ{��Ü�yxb�P��s4���cj'���:����>��eYm�^gkih ��wㄝ�N�������B�n��+P=�v��j�P�1̃]@O��Y���hL��`��tW��e�~��]r�t�jB���q�r������Y���ŦΧ4=��2;�!y�go�>�	�Uv��'I���3����\
��n�máОt�H��2�HC��A��Œs&|r|k����]��-�!��(���Թ�X��TC
��W�C��Ï�#J#��o��bq$�vc8���6?2�3��k@ �ⱆY&g{�]�U')�$�X����>��	N�jNrG]��6Gn3�I�"eK	�@���oG5��Y��r^(<���L�g/<�{d�f�뗅5��*X�#K��
�����歗�f����.�r�br�܃gZ¢y5Y����69��E��-�H�6iRA՜0X޾Kr������r���� ��Wa6��!5 ���*��9��yS�iҙ����QofF���)WB#Ѡ���o���PI�� �_�b�2O��|$Ho� ���?�@��`'�_�ʐ��g4R�gGd��C�"�VU�"�Zd��8�2�xg�K��L��Gv�\��P..����xUW_�����ջ� �i��7�����ʽ�{\�:��*�"�'���z�"R�(���|�#�C�"<�v�����b�g�u�t��q5m|��@�G���d����D��I���w�9IxLR��|�5�k,������S���u�x�-����|i��]h� ��2D�x�^�"���Y���8D�VbT����
���w#%�`HH��Z�wpqד;���JU.������(G#v�)RϷ��t)q�I?�ѵ�����l��-����#��4<k�0��.���{x����z3���66�`�8(��_��/~�%��|?�����;|���7H��|��M�zJ&r&���ьrR����]�W�|F��,|e��q��hC�1�������sb�U�v �y���-2s�Al�1�_��4N5�	�J�A��tN!�ca��E����)��c�{�o�?��in_`yRO�����h��c�=)1�Ӥ�JѠI�K��KV|��<�B�����A��E�8���?��w	U�9���ϊ?ߔ��vED>����8�&�)�@3WqԴ�$Y���ŏ�f��?�t�	��U���cV6�8�RYj�|�3<�bRz�*�t_^�8�C�p!�Q-h	b�[�5%��+����:���M"���R�"^���?��l�|���k�(�/��5�S�u�N'���HӶ�.�����F��I�Yۂ�Y�q:�(��B������7 �%���ߋ���o�-7����ѲN@xl�
���$���٢��p<�I?�1�(<"�;;I�c�%Фh��)٢Qk"������������Aö���C�E�j}�.!��&T2��A����xk�r�漱O�{X�X[Gl�|�������n�ʼ%����x��ah+O��GDmQ��4��� ���C>g?��
+G��o����K}^�]��Ĳ~�Z`��l11@�Њ��D�H�*Qր���#��n�����F� ��/�ab�B�SԉI�R�΃�M0���>��Z�Sj��Hc�3�h&����NjB��!%*dU�yn�=��e|��UUХ񜦂w�<�s�z�~|�m�Չ��BX2����|V��sM`�/ԛ̪���/bXttN�o����?�H�0"k��7�.w@��qk)��#�W
��]�>w;�u
}���J�ce��w�����,�*3��s}�re�;d)#/Z*	Y�m�"Ė%x�-�l: h�!��`[%Q�	jͭ<��L���3�)�������v2?��_�R`���v�� ڞjL��2*}���P����ι��u(�Ӽ�sҫYe~?��%�-��_�89��:��U]d��gѨ�Pׯ"(�����h�)�b�֋r�8Ƥ�rd�7�ޥm�6�� *1r7*���	��7�lЉ4{lDdG����J7T���=��;�$�@�4�[��Ǡ|l#%���]��IUM����v���%�����>��z��L*����5�(�c����(�kfi?v�����k��VJ�\-4(�R�9$�S�x���C��6f9D~4�~��k�~KFL��,�W�-/W'w����j6�"�z�!��e�&f��51�9h�9H�A�O��)��Q5"�[�`�ҳ���b|QQ��@���������'��H�1Y��L��0��o(Z����5��i��ᙵL0��|VK��xK�7�~?���>�gp�� 1�""�Gx���zf7`0��_�A��� ��[OLܗ��#T�D�Y�;� N%�t�w��7���Z�������FgJN��	j�l�4L
f��c+1�-���aT��kJb��پoY�>"C�kH/Eo
�K6Ū߹���T�6m��h5;�~�J۩O�F�X�[:��\D��zG��\���x2�����U�����e��cR�@W7:2��}��w�=u)���H��C�+$�Z5��˔'�	��r��v$������v;�n��/U�M���H�G�{х25����T�a�n��Uh
�a�r.C�o��~h�)��[��У��j��_|b���O[^�PV��$�����>�9������а�,�<%[�Ƽ<�#�u����_��0����u�����l�r��`2
,��5�9�V8�y�7��ݫ��N>���R�x�mne^x���[Οl�
Z���t�Ϛ����s�]�Y#��B�6�A���FQ�J&�ٚt�IL�\E���aC��7Ѽ�:�G6���@f�j,O�s%jы8�j������ ��1'��a`�1�)�tG���>����}X��Ϭ��fXYSՃ7K�a7&?l��-��C )�/g���Xv�G�H����M��.1[�5��lS�j��y>UV ƅ�.�i��):�-?�[~>�m^8�Ww4����l����	r3C�p��;w���~��~��\g�C�z+ ���o4�<����IA�i�S�\UU�o����=��bjr�65�Ŵ|IP�����@@!})�Q�}��*u
� ����
z�+�Lj��[jŚ����u9����E�U�o���<\�*�r
o���)������K��w�L�Mk��h~��{�a'|�B����@Pk;�		]&����α����a�@��7���58���J�|l��g�P+8lk�����X�k0z��=!����Ei��a� �4��#��t˙�\�N=�A.�����i�s�3��R��r���Bf��,�%�Y���t)�[�9֊;M�/r��7�Q�C��#�����r�b���Ñ�S��>1��O��`���5t�������U�X���g%{1�z,�^�K}��a��Ref�\l�CP���� 6�u'��P_3�U��<E`y^�A�պ��[��)�1�~��j�
�GB>a{�W�l�Ɏ�����|�I�!���~�s+�HY���̌s�����{�Tq����h����"�W� *��=�tv��	coC�Π�md��В�-K�YJ�y.I��*e�j�\8m��-�����"	�����u�I��O�;��-�b���;t�	Xa�B]e��Ɍ>�_��E%jƎA��Ve�M��0�����t��~��+�K��!�T]ϳ�_k�N&�.�	|M]5R���4J�P2p�D"�V0�ٰI� �����Ç�S�D����/��2Mj���p�G>n�6e�Ǹf&��]3c��*X��F��U�'S�{@�a�!����\/�Ti=�_��w} ��C���*���c�d��b�gn�7%��!��N!�})y54D�9( >ϗeMh�#4�� s�$Q��ú�-�@S7#�$�hr��v����z_�)�A���˻S��}����򅨫Ќ�*��\T6F��r�	�)>L_,.1�����g0�G�9E�{Ő��]� BR���-�����*�[j�Ya�W����Yu�0n������j ��#zv�`i�,ŝs����p�����J3/LхԦ�wr��H��<�y���?����y�)�2INҀ�F���' �����y�����;L�a�v3Wm������V��f!� �����;>�HG��ú�"�OJw������� !�i��	%��|h�O���_�,܆�A�8�-_��5�䎢�J�>] ?�"�/�E.ؠ��å�4�RA��ى^�j�N���T20׮��`���B�O^�� ��E�� �� ��Lì]���YR|`�E����l�Rk�d� �@�D=n�e�~띁�gtS�0]�:D+t������`⵩KȟL�����kv;�WM��g��˥;�f>m�V{�Q�\����, EF��V���ޔ[����ټ���j:q�� ��Oʎ��E���Q�@`��+;@�	n�gMguò��f"@���0,82	�(�sIv�dƭ�c�Ӻ��9��,^��vm������/\�LLf�/��
�렚ѐ���m
�0�m�����k��QZG�/݌&��p�N�ې	F�@U0��R����j���q�l�M3ʈ�D����
�P IE�I۲)�����`�(���E~�x�mu�ht���֜��7��_�[{��Xey�.0���c�RUi��:�=� ����>l�S�YL�o���];��ʨ.�������P�$�����e5QN��^c��1p%sn��9-'C�����^�5��<�S*\`�\2Ɖ�7���*�Թ�T��<S:?��{�<���4�$�nOD@ )�a�L�����v�j<�?kҰ�?L>�ޏ3O<bp�j�5��~%��e��?�`�"W����
��%d��i��t�E�I1�B�xr�3l���1�$�
q<���\���pk����_3+j���/���������ݨ�, ҃���uMR�!�QY����J�Mn�_k������
-��C�.ӻ�c���'�����*�{��m#{��H}�
Z��K?��O&�O���-�kZ���<Y7�͟��f}tu����4�i8�-$���@ZZY�����kCW��X�s��[@=��Ѧ�3 n�뼻�����?���E>4�F-e�C��%K��z\ �P8��xB���+D�m�W�R]�\��H��c��752g�'�D��].p ����j4�SX��`�{�"�H��%6���+Ib���@T����O������uQ�ŗ�⮀���9�Tĸ�ߏ�z���M�M��i��V'b�������I*;����)��rF!���((p0u-��V�̶F�7��V�o+N��.m�g"Jw�a& �x�Ri���ɞ P���02谋+����,�iNfY����_w��w��1������9���`�e�_�5&-#�ɥK:���iC���߿���S�>�g3������?	P�C�9�)�Nb��}���ZH��:�<�,F[ҕ���D�uֽ"qm +��x�7��K�,(4Dq���<leL���܎�H2�����eϧ��]9ɹ�rѻ)w<͸�u�!͍����Dqk�o�ُS82�$�y�jn��ךK7�TBu�l����ߩ��h�� M�5Au>)E�L���^���Y�*kɔy�����Q1���aa���ދ}F�R#l�~�	??�M��2���� 4�K�@T���U[!���
Bզ9�T�<�w�����O���d��ޣ);��o�0���*ꞷLB���10��W���3��3�;��nt���'�@Gqs2��׽R��rH{\Uf�uE=K��8�f��DJ���4H������rv���>J�f�[oC7ST{N�'��(_�-��_�7�+�=�r�*�6RC%�Q��E�
:�}����':�"�� +�s;�����
�����_Af�HJ
�W'��*�=�l��*"��җ��u�34#8B���e�V/�(,)OmY+������ӣ*���zw��C��-#�NEd�����&4�@�s�-g�y�[��{���oT��+E��8�Wp۟j�`U�g%�Mj`�Yu��+P�	Y�����������,�[Q��ċ0��]��g�����si~�������s���!�[[,W�*�����Q��*�m��{���.q�8j���?C$C"d6��,F_䙫�<�<ł2,���G�iVpF�d�1�t]�����v�b��:��la�o�̓=��~Gµ��t�˚��;=Q�d�&��څ�?C���F��l�DT�<n�ڞ3���)VnK�O�}���W�~%]w����=���]9|'/��y�?�������k(����`�&�S(��#���	�!�Ab��Z�xL���)�t�l�nא��n�_y�"a�P�:mt8%��'L�0H2�6��eSO��f�#���Ƥ���[;��Io8E%��m�����l�^���Qp���U1�ͅ|���~V(���9:���N�ߦ����?��QC����k�����,n������W�[��}��n�R���S�͝8�Q��&ږ���S1�fK$ㆿc���T%����R���������ܒS��y`v�f6+:���0h@s}n<�p��u}?�
^��WKw$���G3���K�z����6�.4!S��mMU�0Lc��9�����ˎ�Z�)���~U{��]�"LY�G�-���%q4u�|�TC�}��w���� �ݲԃxnٕ0�Q�cq
<���`�x��: ��H"�˔A�UJgG��MW��:��T��� ��H��������,`s[plA9��,���f(��$2T+
)tyS`�z���5`�k�HDUtl���|_�>@�!�֤*̮p�%��\j �z��F��'l�� �bV�P�";d�`J6�ILvciK�8&�Wl�0�kd/;|�u�����F�,%�Pb��>�\�Z����&_BT_���J�q����xAObڣ&r�b�($�s�LCL�)�H���Ǌ�{�(���oh���E$����^����5����Su�yyT��äoYb\��9�:�(L�AI?o�x,��+}���<g�O��x����薜�q��C�3G�w�wށiq���B�`_�Wf��|�O��6,��V�Sp؈+y�؎��qc��j/ݟ��&L�.d3�����%zU���[�DΠ~=5��,l7���S�q��Loy-R3�T�]�8�Ϧ���r� �B[Γ>H��P�fwbgA5��1�τ��j���LUEW';���Ca�[
���ءzO�kj���n����mm>��.TЗ>�~��k���u�_mº@[?7�:C~��G��t�m���Q�"���'����Oe}�ͻ�����?~U����-��/�y�ݕs'��$xm� �Xghmc�S��w�t�@i��4�B;vs𘖐y5O@jY��{%,�I}������lS�dd;�3�*�ڠ�����S�������yB��jF�g�!`�M!|q��&�oُ� J�R.K�|~}v�3y՞}ʝ�B@�=©V�d�hj�~+ W+<�F�����B�
�&?�*�u"�_��ч��{�8�[������[�m��J/��]kҎĭ�G}���
��u�E�O���A�HsG��;ӌ{�����$7��&= ��m�M��9E��p@:�����Y���`#�l%���c���]T6��ki����/X�EH���'�g7� ��&�D^�T��ir�#xs��{c(A�ɴi�4M�_�K
��+ k�6�~�Bj��gX�oÔ�:�:N4+; Qe"�!cS}{���%��K�Qs�w�O��x-���˴���aP��AD�wm5���&��Җ���՗���]��d"З0^~w/���k ba|�����q�h�}]���s�(3p���׍��f:>@irD�Y�$!�j%)k6,�-u��}2��%��a�9Z}�U�C� ���#n�sЛY#U�c	*��x��j��BL�gP2Aq��x\�nk���U����$��>����WT}G�̾D�vȏF)I�!��c[c]���$�2kq����jf���lL\o��/��ߎw��Ǭf�,����9-��:8P|�p�-�t�G .�7����^��Ou�����Z!�-�W�3p0IZW�Ǆ%������!�mz�Yz���0>M/��qH�=`���dL؛ST]3ޢ�j�lC�׼*<�s�ɒI8�d	՚B��,p���fC���G��	��,����O �sš���oHR�������t-<C ���� }�6:b6�[ߕ-���9����i6���y~�3Gwb��\�CβY�&�	��{3�b���u�s�I�n	Cx-���k�X���:݁j�� �f��(�ĨR�e�H��<ТN� ���N�@]4��%�<�&�h#˂ڭ~���b��@��fN���� }��q��D��C�#W�Ѕ=��ĿQ}?�GN5�D��˼�V�q'M�? ?\�t���AgQ��5:	T��9���s@ H�;�~>SYD*���X��c/���b�@����u��= �7���C��QS�G��h�����Mp�1;PƆN��4�G �${Z�В�P��7�*R����$�14�loFSL�X%}&�����{�Jz8�(/�H�(�F���v�HJr���Q] t_f$M�c����F����/K�_�x������]R?/�+U2ow&)�ġSi��~(�V���(�e�QK6|�U�bUGk�T�T����i�2�t��K��T��U�T��|�4��"-9��o��=�R'�K�d�~��2Ό��\}�'�T�V���ܣI���#U��+U�KIK��>�"@���E�$]ɓwazӏ� ���R�ˍ��8x#dwdr4��HYvŰ���/��0ч�O�{����S��&�׻��OE��{7aD^#}�}������ߖ�3ϗ=Ȥ���+�b@,��kт5y<'�Dq���֘��)޸�������Ϯ$&�X�(-�<|��b�w����Jx^����
���+T�"xY�?5Y�����O�*��$�	D��PƦ^����}����`�������������g�,	�R�bi}R�&�s���Ϳ�e��	}��Hk�G��XmZs�H�Hf��/zk'�t�w�ǃ�������r��Y}�5-w2ȱ��m���L��J��r҄�;h��@l��)c xZ�ޮ.�IS��ēz�c���݋�?�����<x��\��@&1!�H�8��p�R�+S��|����ZS�t�����'��ehfD�p��Uˈ-�Ad�ġ��V�>[ֱ3́�~�k��ug(�ȷ)(�C�p�e�M����z����`x��1�7C�لM48l�	�8ů�Av����fq�[��W��!�Y�q�]4��#��]��L(���q�"�|�7�ӎ2�b�F�$�����ߵ�|�pz���вE��W"�u���s,�~X��*:��uL�?oh�)��F�0IŚ�V(��V����8]��X���Ty),�kĎRh�t���=�S���%.N�>�vW��&y|k&[S�T���B����jz~�hx��(�Z����L�F)�����۸ynL��Ǐ�oL�6<0��v�ğ�J��-믤9�t��J�O;���Ho����(����.�pؗ�R�	�N�G�T�66&�Q��L����_I���$ɉ��U�i%N�Yz���ϫ4,nw�!0mw��l�=��}����J��+���DVi�	��ێc�'BV��M���������͛�M����iz�L����K�3���L��|稁���C�|ʮ�	��v�sw���pͫ���(�4�.Ǻ���#b�5�𔜛W�j��H���4&6vg����yڜ�<؄�ְ�p�%&	_Z_�D�}��dJnm9��k�τ�]��rQwO���i�ĉ��t�]]I��FU��kTo����,��ME��օzA�n/4f|�l�~�u���W�1G��0�_^�pū�"E�O�)egQJJ%B�q��^��l�9x�;�9/]���c<Q�m[�阥��s�CQU鉵���meBoM�@�N�����l?�>:��U_�┆���m�O<>��g��0{i�<6�D��
S��[������ aK�e��j
	�Aڜ��-���*)���{�)���C� `v�5t�� زg��(����A��$5O�@���㖥�|^����e�}�J��7�)@���/��Qȁbʅ38	�7��e��ћk�^G�l$�΁����^����sLa�ub9 =�2��Q)ˈ���?���҄���z��V�-�Xe2;���9Ԏ�@��"��Q)c��Y&t`������p�qt�1�����P��H����v798b����A��ܼ_1��1�WP�V�Q�AE4�z|h�ی��s�E�%���z��8��oT?,����n��������l��xU2���[0�Tfr ��P_d���3duG,N������#���T�dћ˼�5A Hi�T�@v/��s.ͮ4��߃:s��<&�_�A���?�;���ЁA�H�n1���J����t>+�D�pO~��0k,. ��n���D�R>�S�]��z;���������H[�}�
3(�����~��e���W��N�v�g9M uy��s�\{R.�n6� ˫4�G��-�3Bй�WQJl�*�߀K� �:�'��A��� ����(�*qdi��ƣ9'��=>��'��]m�6u�q�$�6��:�w�λ=:r�@/M����Lc�ܵ���7�v�j�eߔ�?���Ӷ�VL�����~�� ��.��9�Gf��-��3\�8\�k~�����M���� *��B惭e����Y٢;������ȱR5�k�����Tv�y[�'�?A�V;��{�*��OYq6x-I.g���K�	��n~�qY{�d���K\<��X�0�9\��DL�C�z�`z�êq	��7���m <[�
���\�#��;䃨�L�Ł�,�2�^�1rr��K��Г�ȧ��fӳ��%��PKЖ҇a#�7��<+�/5hu��q �t�O��|�&>��w�C�7d��Ri�4,�5� }�I�/��|L�#�ze��R�L�7j����5Me.�X�3���I�-gx5�n��]��>)�)pS�~�Z�����p��R�G�m	��م����GI�u	��S�Е���;�i��Re����R#W��"݈@ER=�t�i@��X���m���G�Ns��i��k��i���J�e��/6��Q������:��e���90J��N��{�lP�-iV�`�ც�o%l�''>j[�RCj~6*�oS�O��+��ER֒s�M�z̜{�B��V/��5PiQ�jͲ�,��� ^���^Թ���gu�@�/�?����R�5!&4�^�N��X��O wu�M�;���H��s�'ߠ�嶻.�h]�X1p4>F-wP����� �6�G�	BeC9K�p����3^3ӟ`�ے��
����M�mʅ��]�R��x�<�,(�p��f\h��ɰ"�z<�M�J�Z�`[��D�[�nV�1���c��s^0�#᾵$��tV���1�ҏ�d5��ᩓw����%��z���e��a�v��ɦ�kI_�G���T�/�_A�����|�f�\���g�����M�]�47a"��t�_@Q�������'K�$zO��$w��T���L0�̎���za�Qf����/\d�d�J�l0�y��FX[�Q�G�|��I'�?����U���!~��Qޖ��Z�`���|�� ձu �T�o�ϋ���Y%Ųj�"���3.��w�#�D�#��u�P�����?���(T:��v{�]�X�=RAQ��Q!&! pQ�a��da���\�BKxE��Uԑ�O�
�V����B,�KU��x<8N�t;Lz�M��[��*�mAvǊ�e���q��|��6د�|�Ը�ݝ7�2%����n�JN|�醙��ZCx7�{�]�z�ۙ��q��W��"��<+� g�'Ȧp�)�1���KsFc}}�k(��6���r���on6�ױ���Jxk�
r`��W������Q-�e���x�'���|.7%8g�=<#��im�9�������0u��K�����`���(,XS�t����F��k"�3�(�Q��es2m+�� a9p~s�O�����h=1JR��NE��b���'��r`Deզ�dp��W���6�[k�?T �K���񶑔_rh�����<u��G#lJ]�8$���'Q�Y=�X��@8�t�܏�Q��ƕZŧ*fI��8���7�������Gu�Ub��~�c�BDT"�{�9%���9^γ2��E.e�/���
)Ĩ��O���̤]wNGX�3��7��Tl�����u�bÂ?ޑ�b����8�4+
���aK�Mӛ����V������L����r��tG ��-�c�F���+Z�6÷�݁���[�b��K�3��h�%F���@����S�0�
����jqo}$����z�Fg!���.��_�@�ǹ��	����A;�Ei	}VB}(~	��.��6����P ��mD�y���]ݜ�]i�M��<����� Q/�.~Vcr>#B��D����K������
Y�1��$�k�\�F��E�QmV�C^G;foz��?����z�m+�7��Jd�+UN���G>'[a]�ª�M���5���uR� xc��,��/����ø�K�7�����F])�y�O�l��MaC)r!V�!�`=�A��V/�U�5L�e6�>��m�ӿ	zd'
��y3���#6�G?m�A$�
��`���y�+����.�c�
��U���⭸����;ZC%�Z$��-�FM�v��*Mf5��b	йY��Pز�N�����z)�U	r���:jFq�W3�
�!�#��K�+���[.$g.#�P''ih�n���U/
�yPjĽn'/���V,ޢu���2}�ڑH*��+�ҭ�\����q)~�����I��F��ʖGo���]�� t1�c���.H5~�R��~;(��;��?m���=�V'�;ɕ��Xjn6��=����+!=Ȼ̢O����.�$��I�0 ��:�Q`�?��b��l���j<|�mJ�������b3��M��:y��AR;����z,��e�5$�P
2��ߧ���K蝲t�!ڤ�k{3�L?�mb��:�=x��@i���4i����tf�L�ELU�E�ff�֓v��������~��z��S����Fk��{���.�.A\*��%-5;|��Y��jߧA\9~�,��q��B�Ϛs�J�ˁ��"�2Z�)��d&�:�{/�U���Y�qg4�Z�|���lJ��Կ$�@Z2W`�|�;�.��}k�'7��A�LH`-��:9�Yn7�+��|��s�._���,X�͓�Y�N/��+>GmĿo���J5�yR�`���적��9l�~(�xj��Q��?�u�Q�Σ"���k�2K	��ץ|�]���pQ�RG�n��9P{��"fOl8�/�UBxj���{"���D�}�v�EK�K����t�y ���C��M��^�7Z�/��"ɮ�.�>!�Z+V�Zf{Nd :Ky!y� ǿ�<X��;��5J���^�k�/J�6�Ƽ����m���a�[qyf� �z�^/@w����@���L����Ҷ�}�N+_)�%<�-��������%���u�I}�:�
�,'%��k�=���t���X���-W.(��F�h?Km�ʪ#$��N�a��~4C�t� li�Ǡ���y�>uؽ޳Ѭ6�o��5�`̟�E��8��_�yRoxA��SK#e!a ���4�� �9���>�ǉ�	�y| '`���
3��ހ|�.`��bv>^�h�/2�M�G}G�",��.����+�h9IWj%᱔���?a��W"i��Vf���"#�������G�Cd���:����cY'_n�y㣌`4��W?J܋����'l�a���~��)7dBX �T}[;Mo����*4���k����F�G��1s4d[��vgj�]g�d*�� ���o�Q�O�i�So3���~��C�
Ëw�h�b�[Hx�Q+��s2S��4A�"�K'֘����)�O,�7+��7���T�s��L�l���:�m-��i�0��J#4E7&o�~�A����G��NR�,跮�'�AA�a�Ǡbo5)�is�����Vz��@�YpF_���
�0��I���TxN�ʥv�eX�y�0�F4&kBV�,8�{�W^x�A{��|�IW�Ύ�k9	C�P"� �
�� �2��4M��~J`<Q��b��ڱ�̅��2��q)��Ju5��]�6�0|~��r�9b�,W��e�0�{�ƳM�&]^�
�k�����ѿ����*\�!<�u��m�����:z�\�}�[�fY�(�����)�u���\!�����)����Ouq�90�db��$����Ϻ�,ɩs���5�J���CD'�:����W�9�,�̉N"w-��P���K3�p���Y(��cOZ��,q�8�5�?����E���O����T�z������v�A��B>��~h nO�D����谚�5�|����fݎ3}8�B��E�Ą�u�no[�1� cgS��t���(��0�JE�6�|�
�M�����vG�:�@��$�/_�'
�#<D�/6.8�������]�j���8�O���i��
��k����G�|i�N	Շ��/�FU�_�q��|;
X��S�T}�	�O+��w
���
�1A����?�7��Y��aQ�堽���o'3� ��b�s�~8i�
�`أHqx��2��u�����ݡ�gd��a��*�����5���X�M���@�-�����C:��,�n˗G�R��ov��Q!��ສ��P#�H���v4m�j٥^�U�ұ�z�}6�N"S3{-�:a]��|�QOȁ�0s.�8)��g��/Q���v)%Wo5l�c@|f6M���'�;>[>�^N�ΐ�QaGH��M"4kS�Pt/,����a�+w��4���Pӭ?�G�ڛk�E�	T��l�C�����xE��qtJ��V���&�F�q@.��E�����KT|x�C?{��&���v����q�9���T)a��j=A�䫧E9
�E����_2[�tn�郡������Vۑ�����eR�far��6�ã�I*gJ��r�ɝ��U?X��i/�/�G��I�*��/^C�������6�����Lq:y�5����v�G�(9z>goOlm�tͬ�wDQ�3ސuC�eIՐ������2���b����Glf�D�s8��
�?�� ��q�I䎢BV�$��3�k��sJu�C��_J��'�w�ϙ=��c�Sx���64���A4�G��-�<`�kg�UP��
�Y���f�}�_��K!e�[�2~^�˝�6Y�7�H��Ō�;�M�/,*A���e�d�+E���P1G������N0�>��Zڈ�=��9yaXU���sd+���d��Fx���u�o\�uh���)�J�>�W��7
#��q�f���G^3��d슖Q��:!n� !F���4I����8o����l?�sx��p#O^ a-��|e��p� ib�9v%mM<FXq�~.O�;�U����<n�b�@~�+��I�J�����HxmӬ
�ʵ�lM$f��;Nj��O^�*���<	��$���%�r�)�D���G*d�7ȝ�Y�S�!���Nq7�����R���H�B�����c����VG�)ixo������3cA�)����[9O�cEn4^�j ��ٙ�G<e^�Ƌ	``��D)E[��6r��'W\��T;|��t�v�/�������d6�~at/Ͳ�N���v�o���Az��l�(ۡ@+�7�-N�&1+@餺D_�n���Yhɟ-p�HW��� e�,���B��ٵ���$�=����_�����o���{�4��A 9�`���wT�~�'�+���	�[ɻ$}�vs0� $��Ri<��ju��[�`a�$$�vV����F��J{�Z�=�{n���z�72�����' �9�8�S1��͸=�j��4�=�����&ѧ�?LKK5G�����''Ҹϼ�Wx�f:�Q!ۄ&�DդM��f<�,<�XD^�k�D���-��n��Õ����tf���{�Q9Sk���-������<g^�_6!�w�a^�޼��i�!�����.�@�B�.����{����f m��!�����c�ʔ�	��E�������n8!��,��F�����qH����Z�@�(�=N=S��)7ȥFe�&�U���VS��W�7��E�2&�>��6[3BxЁ��tQI�ԭ�Eơ�b���l!������}�Rl��:^����%�L�D�{��wOȕ�yǁ�NO���_2\�!g�O�0*�	׶m��v�G��8N_L��8�># �W*P�ƻy
UV{����h,���g
��i�sml.���(]��t�.�/-��9����i_��o�Y�C
Y��)�c��3y֕�u��z�*(il���w
�²�7�#��8'/-+>F�܇��7��`7+?�+�
�BD 	�Z��g�����7�N��?��o1��8��b�,ZѴ vL�+i�7�9�w��ߢ�f6�,-�	.�W ұ�#����{��2�"���ذ��Wg9?9d( ���!^d�|X.͎�Í����PGM>��4��R��_ޠ�m1�I
B�R��D2�L�h��у�L7�+�{���K
��'_��4�;ǧ)�xb���-���=8�m:��P�o#4��X�H
ʝ����Py|!�>̛/$��JW:㿙PM���=�ZL��f��h(?�:+DG�C�K��0v�|���x�G�﹝�Uz�N9��#kp?M[7[��&[���a
.��gK��&�vPV��B�"[\f���@��[5 #\��gg�;l�/�M�d��^�LL(5�r$b*�w���]���ț��hB��V�M�7`���?d��ޚ��>w�cQ,#B�g������m��D>e`�����$WS��@�Ů�N<�T�y$
Og~��/�	�2(�HY���v0G�R�p_��{2W?��:����@ 8ۣ�	ہ5m7�~��=%�zE��@hi�����+�&��+.����������U�R�p��x�|���@��6a{��տ��Aח=�0�FY�˽h|���Ą�G��H��ķ�/�E���L: �:&��`��	�<6��f#	-8�2r/���T�h� ���-��G�G��S6����(ᔠ3dm��*�Au5�.�Ԯ=����߸
����KH��z	*�͵E��w�/_fNG\�֖�wu4�y`��ʓ��$��@�K��0���r�e��uٹ2 Bi�m�vhG�����^&W)\:��UnNP�<�s�^���z��붿s�Cq���O�L��W�#�**�9v���h�p��-�>�+�@��ˌ(ſD�F��� Dt�Z�\k�kJ��8��A�b|]Ҋ�)�hv7�:Q����`�2�\?Y�Z��xyM e���r��K@��íS��hU���������3�H��s�|[K\H-[u?}�.i�VD��H����a�2���0?�=�a�ĖbT�Ƶ�i��'8����D���`��Yj��F���	aQÐ[�_��1�^�s涁p@�}�^G�e�6M����	Ǫ�?��:��x�&�툯�}d��F��<C"�v0q��$<�䋅�B����)�,�gLAu����f-�UЫ�j���qSw4�3`����	����l9��ԛ���2����ӻ�8�j��x��3ay�u*@F ��92P<���]�.�a�\��?��P�N��M#�]�k���|���iy���p����
�s���b�ՔN�k��e��pUg���#/E�d'��E�4�9��@�>�Z�������ʚ#Ua��Y��t�5��=��Nw9��f�tl�`�4��0��Z,ؖ�\���#���������x�s�w&
��\P���ɛ��������n��;ZV�#k:x0ш�J�?��� އ^Qk5/VK�呣��ҹ���z T~>��Q�)�˺���U�K�؜R��r�����Z3���w�^b7��`�(Y%��>7�Pͦ�x�?]�΅�}F#�f�܊�4_���O��	T��c�#3(���"{̚@����N��oi����azv���M�j�zu[)$�Kwݝ�������+2<h��<a��Y]���_��.X1��9���Z;>5��VA��蒸S�V����j�(�?��bXފ; �u|6�	���}�i@�Z���!ч�
���#Z��*�����Z��8����f�&"3_��ܳWC E�q;�F��Ѯ�cG�x� �җ�=�3��� '&Y R�G�����w����?���a��SZ�?	��%t;<?�~�1T��U����&VĀ�`t4#�AC���^�$?�<:�-Js�q��զ\
}��py����Np�\1`_d��)���S�Xr(��k[�K皦\g�3�I ��`/�����3��K��+	w#���7���J���������u����R�*P�X1끦�	�g����E����NeSr/���Y
�'8~X�$j�LZ�&Ҙ�Z)]ra�]�ܣXv��M���N�ye`/��3�W�d6��m7E`�nx�Ю��h��&f�tHpR�8}�r�+Ĩ~
�x�����#�o��%	���FH!���w��[\o�a"���M�u�/��H� �q��p�^g|�dg�=��s�h)M�:ZZ2���halK�㽗��K�:}3й��Dӄ�~67���V�W�?s��\,qtR3�2W����1�_ݸ#_��I;��!��Y����D8���	f�\Y�����Į��o��-�"�����	V�^�/'��0�[��/kDT��G�Z��/��گ��b`ǆLM�j����h\>0���l��V3<�.�DT,}���-A�v��n%��$|�KU���*�Bƀ�Vr�!���K_��&�W�SVwٍ���Ģ�V���UaۻX	�/l0hA�͘O��l��2H��l��WC�o�=�a]2�cі�F��M�Q�!�(�H=��4=�M&,Ћc����9��5gjl>ʃB��V�|��
�8�R��G/�:'Zr����-�$�����C?L�nl}�\������6��g�i7jV�����Oy�L��i]K��a�4��T���5�<_�Z>�7��@B�b�()���V^~���
	�����R��Ӛ@����42O�݁�������[�A�W���*Dv�)Wͦ��B���Y�-�C� ۘH�����ȮA�H�$�vB�fi��˧>���	rv$'�"������]��w7��9ƺrl�)��_�����A ?U�R��=���:q/��ֵ�2�V+��(��}���#�\�>�<�՜�t��h)
e6�ڐ��8䴏����1,'�%민�M�L9$��#�Jm��D�uX�����0Mn�8\4�������< _9�L>hA��`p�ޑ�T ��{��-na���B�?P��U^�O���pЊҡ��KL����^ �|E�-7Ww�()��ez�����?ʃ�"��K���=\�M�պW`��Y����4!G�>�c��dK/n}���"ރ�8f9��ȒM���n�e��J�ݶDf�����2�s��D��#F�H!h?���d삨�������{��)����
���m�Av4���p��98��
�A�pyK
Q�ʨ<F�����h��^J��n�]�p8e�|%�׮�ک�N�Z���\�P��^�!�y�hT���� F�/\d�0鵥v��KZYѫ�,���ɋ9{��Q0�w��1��7�8VF-�3~�e1Y�膝9�Pل��6rE�"t=Â���[���3�u+q����t���/���.�
	f�-,���xV�����;��a������zҿQY�-�ao��y0Ү0UUxQ����yf�ah�R� Sn���w�
v"e�̤�5�T�䶶�{��\\�?.��l��H�Ē�T���"�K�m +�=���Y���Z̩�ta�B�zB8 ��p���q���tM�,v������H�z��;3��4*ʜ�Q]+���/�)���χ�#qL�1+����mGX-�(���X��	�R!?�,W]�2�S|༡�*U�/�T/U��{�	Y����k�6�()��|��=�P�<j��.���������$���7�
���PZ0�ƃ���L�K8���p�8��i�_��H)2pnբEƒ��L1}���/u�#���($e�8@<���8#rk2���<�F���/�j^�KG'*V�Ȭ�ع[iʯ�±l.E��-��	d������:�de^�0���0��b�������`�$�����'��H`�T�x��Ő�s��h��,�"ה�oq~� /�N��Z��B�9�
EJIo���*%�F4��?`f���ƒ"L d��E��fGj�A��>���E�ʣ%O����1ü�l��Xku�dѾ�?�u	JX��V]^\��ƕG��R��O�"�`�SL�@?�D��r�ʁ���'1�{Zjdy������r7�X���k�������闭��w��<I��DL3w3�)E7��� ���ʞۓ���m�c��c߫v7DfI�Τgt7"H�����%>i�hW��&�o���QK�X�.��,&�C��0ڊ0$���{��*��~��gDӔn�0�]�E�~_��t�	�M�D�>�����{S�l�=�?�m�&D?L�ۮ�&!O�(� �!��d�4K���m�:`�]=�7^d?�P[�o���O��m��/�Y	������/�v�� �9)k�*�O�l�%��.�7����Vv,p���7KV<�G�F6y���D�у���X��N�gY���큆D7���׹Խg���7ď�TB�s���X���$�6k�Ur�vR���9�xF�J�(Ȅ���q,%;,�4>��`RF��CX�9[�����f�71<1�>��L���W]��W���CS, ��)zm��8��b"p���"̉�����U�[�l��&�i�U�p+]�G	G��̚��	>/ dÃp˞�5V��-��^�B��~2��ϳ�ޟ�ث|�`yQ:ޕOm�P'�����ť�J�ܪ!v����=Ay��	n�GE3=J��ꆟ{�χ��!q8��Z��F唼 ���,B?���uf�ʓ�~289�a�Ɉ,նAa�ĬP{גU��Z�Btl݄S���E�B��w:C"�쉏������'=�H��<�h����������A����ˌ�V�/U׋�<��f�,���q�0��<R�e����Fd5�F�O	�Q�_��@K�B++E���4V�_�F�N�G\��ja7��D������4u"�J=��Bu�$��`�D�З��p�;]Oap�P*�J��گ���8=:�}��@m����V����R?�H[�h7��X�� ��I��<$/_��G>RK��B��7��t��E5�#Ӥ���EW�.��#�Cٕ�9 c�m�7%�t�}�yB����x�)�;?�І�n���T嗿����fX�iw�\]J���-�'�2��$�N�gxH���!ߓ�`<++���%2�Ҵ3�6�ͦ�z/k�õ�6HŨl��Zrc���EQ=�K��������$uF=�V��|�8b�,��5(��n�޾#oD�U>K����Ņ��5�1��"�x�Ӧ�o�w	��o�����B���e�O|�T��ȓtu\M+��J�Т�ɪ*���6^� v�g�'�a��BߗG����Jvw@����WJn��\Nf_�|Ű
z��N~�TÝvhLc'v���?Cg��U�"����R��Y����U
#OxzQ��S."�/�p,z�.�N�z���;ʘ�����;�ʥc����Y?��l_���L_ő f^ �Il�j
-��H��k�i���v�������]�|>�I����p��3mӁ�
U�8�TY���C*-�#Y����)M�*=��+f;M��|� t�W)މ1�4{}��O���79Q��(a�b���9�S;�˝Q;-�ŞB*j��"x���'�*�~}�N�̨�|قN�҄qhn����1���@?��֒{�|��,<!���(������E���̔m��vvEA�81�������tA[\}Zg�!i6r����1��2��������a���&�4GF�v��sv��[����Vw"1f��-[�i��g����bg�/�0�'��Yߏ��B؄@1n�?kH�$Z�'��_ُH<��1K��a�`J�N�n<`:�w�0��S ��k�韜ųjۧ����/�-�΢�E�gf#I�p��"����1ې��^`�Yx�"<Jw�Gj3���P�n6���v-'���p�3U���דRrl����EA��|���Q��{S�a�����	���ҴV�]�Opo�)T{�	�_�m��C�2�ڼA^\#ǔO�LM�}�����I:��:�N{��p��R��hK�)��j�x{{%FGN?�cI�Ʈ��}+]��1Psd��߭a�-T6�	�L'�M͑������v=��:����Y�!mL-�Cdoe����`IA�d}�F�i���
�Ae�]3Kɬ�Π�_�S�����?#�8�ZI�A���`��s����'� '�ܬ~�;,g,�DO7�#&�o��s���>�Rv�d�Y(O&yK��}7���\�!+�}݁���ߟ!M��XϿd(�x��u_�e���fIf�%�{z���i�Q�:�E���L�G�8�ݔ62��PX@�����oM�h���]W��qp�gP%��^���
���݁1}.#�`�g����,W�x�W�8S5#�'��P@�N����b��2Hj@łJ�gK���f4�^�k��o��K���r���!Pi��E7�����`��_�K���`ka���cJ�n!�ΐ�
ްA��4/�ϖ��$��{����������Y��d&E6Ŕ�D-^���謳��J�W�~R�}E���x��yt}q�@��p�i�_rN0��I.?�A�r9�� �0m��O|@̜����"�6%���o�H�YK081X+PUnNR/�4�� FC���TP�/ö�"��}��t�
�b�%���XN���Wj��s���`�
�~(���V���U���x����a�M�N�o(���2�����7D�����L��E71w.��/�F^'�T��q�H<�\���Z�a��]@I�]}k���
��	ݑ��є�����CXs;j*��:;�(����i\��UxG�B�x9�!fwGnvv׶����<Q~��~���M�yC�Alc���9u���U5鰃a[���}����z���L�I�^�R��h���v(�����"�QK��1Ne܁l/y(�R�|ꔂ��uWZ"}s���e�ۦ	:1{
����S c��$�Sk���s�e��6O��p)���!#�xQ��=�0��t�Q���"�� B�^f��#<�c�?�l�]˺�_ٹzZ��D�W�:H���a�i��܄u�Mi\����3s��	"�
��\�	����b�/��3��(��'�r��_S�{�E2�e�%��͎�N�T�Z���X�'0�Qy]10�@�Zo��Q���5��#�4�/�+�����u���l��U]FHW1��-�\���	�9��r�e��w;�M�89i�E-*�09�K9H?���Wɒ��9�� �G3K�	�2���q��0p��e�\�`�v���H\�i~c�[�3�/)ۙ� Ze5}�*~4�E�i���9�΂�ciN!tD�m z�2�ټ��$����9q����_>mAtA��΍$�9��⍅���D�
�mT�?ts��q�L�e�L�o`��{��Ɲ�j��W��U�"��+A�(���u8��Q2v���U轓 ��I��#�]i��d��9㨡�U��� ���q^�����s�Y�I��|9��u=h95ã� �o��ZTZ���9 ��X�h+�qZ�+��鮭�+������*�c��v��M����y^�̆�"t�\>�y�ъ�B���G��W��>��ju3���|���׾����l�Iʯ��`���$�Q�v�X���ޯ��B`c{���T�l��/@�x�)2�8�S���ܐ	�sg��>�et�h�|���e���@2b�Ft�:��-��V�x�4�v\}X(������
�"��wp��G�5�F�2�A��=o2 �ދ{3���Ag
3 �|�&f���ؙC��lA���2=�7�瞽ϊC�-��PO	"AZ���������3��l;�$52[�7�*�/���9�I�����YN�"��yp�|<@p��^!�}a��ډe�L����<�?��hOc�6ȯ���@ '��~׀��41��.�4�D�h|9�#�g�D��=g*� *� ��!]�3�p��в���?�B�w���Ŵ��N��G�2ʈM�&9��\�D߿��s���C=��B�/D�t{",�B���_25���?!2�Ĝ�G���$3�����;��]s�^��Zt;����˯�^�v���vھQ�|�
�l�S/�Ya1ٝz�D�$Nzr];�FPUC�q� �~::�F���u�n�:�L�A�5�ي�����!vpP:벋�7B�}n�]����w*�)���M�Z,�d��?���鹃&��i��i��<�JG+��E�YM��B�'����3?��e�*^T���kY7�Se�?�X}�R�9��`�8����g[<�c�TZn��-�Ѽ��<Z���H���n��P��� [G	�[5a���%�|���t±E��6S^z��c����u@H��GlX���&Hگ��?vY4������"���k�����!��H8.�S��1�w��ٴ��o(��s�Ƞ�g&���J��LM�[�ܗ�=`�i��RX��򯨄��oз:����tZa?йQ�^'ٿ��|J�omż���4$\p�ahQ{���ð�a$���e�ZŁ���Θ�R�K�O�;�G����a7����Uj�~�K(��>E��y���u�6%�J���j��>
W�([#D/��ЬE�ɛW���R.���xJͰ�e͞�.��Y��1��4`9Z�Ľ�a:�����{5JO,MӜ�YA��ߩJ��}x&��Y���������Ќ��b�#���E��gf�"���b)���ZV�CP��E��ϫ4jh ش���A�w�}�Mh��3C�O-\����9^��^�n��"k��f�}V" �E���7�� O�p��0�A.�H��2Z��-�����̫�j��e'�	!�Ù�4OZkR1X��2f��Yjb�댔2!�?L��������n�{Y�֫��#ʦO�1�`Y3m΂,�'[�^ȸ\Ƒ�T�аu�Y�����8o���%b�#�#�3�-s�Pxq��R(���P-���EE
H����ԈC�p���
t;��P�?*�sg�O|�;-����Iv4l`+��r��z^�~��Ûm��O���O@O�E��H9}�CO߈ߎ�f�^���ͺa���+���/(�8�����s�~���u��`>���0����I�A���l�|7U�Z皐�g`aC�p��W���ڠ��`-Yڐ}�p���e�|B'�P��b�*��fF��3��g���5�R\�R �_������1�!	��pS"�%^*]ץ�11��d$������)U����ٷNL���̘!&Ѳ��Ab�kK��~��kC���+���$�� ���ǃ͇��/�Mf��X��I���S>�G��ф���V�N})r�R*���h��g�$Pb���0�W"��E��󨚶FE}c�-����������O���)[�p��2���� 3KB�+��4TT	��a�
�q�,�L�yB���*�!PN�ug�XA�(��/�(ܴU��	�/Z����
̂>/���Ah���T+�_�
���+�ra�J^ފ��
�����fR�ݱ�4��LR_ZMI��7�:�\1^�l=�Z�z6g�y�т�H`���c}N#�C��	2�	*�V^�"�g	T�����&� +����V���@N`d�������T�1����S���7ϳIp����`Pv��ؑ�đh�gF���B�Z\i��0bb�kw75�g)t*-foM���v��P�>�q��bM̧�3�*�O|DB�$�"��F@�����b\;�du���Q'\���b�4ލ5d<���|Z�'����$Y�M�H)iv����4�����nT�'h��C�
��A-�>���<���������^���]�80>�؂����m�����2kE�$���60�S����[g��dR�5*��_�BP�����E�l��VH$i��%<k�)(��߽�[?H�>Y��f[i)����F$��|���^���5t�5U����������ks1�`ɜ��n>k-�˝nb��9�S�EQ�_̉�TL�*�J����������S7
������+:��ʊZ���c�@.[����߅���S�rJ^�ɹF���Z����r��s��z�\3�#�h��2��J���8.%�M\�H�@��m����I��3�;�Ak�}*��3i�Zo����0	\~?_�n������C��Ƽ��Wu
pR� �zQh�;)~W�P��N2\���r������K!��N� 7�̌1��d*��\�����K�9�X譑 �8���YRAC��TNHC Eb��y5md.�d��4����-]�?g ��0�&�D8���ik{P��_1S��oN��K��+��~#���_��&��Hp��}' ~lj�զ��ƝP��h����HS�N\ ��~�� 6Gm�+^
aG��@A�7l6ĵu5կ(]�>��8�3\<��	��wF�9&L�<94>[`g`GAT�:k�Yߜ܏ku؍s�REf����D�5�{-�����!��q�xL"�z�Ŕ%dӨ_
�(F���.��BэȎ40��
�V������1��������|c��fM�Izƿ�.��a6����K%��<��o�I��;��d�-*q�]p�ȏ�P���7��O���J5���Ɩ7.�����s^^!lB��*mJ�g��e�z)��c^$��;`��>�皯�˚tz*^qvL�`��2�i��p�bEv�t�+�}`YlC2�n"����&/���[8$Z���m+��5�_����<-��`��>���rZ1z2�����S9�:^Q��7�h2'��|@Ե��fU����&c�HL,f�x�L2�^0��iF�.�����c8)����؃� 4�y���o��G'�%iU�@f�e�D=��>��_�����Ap�Y>)(
�&a@1;U$�'=����:���L��T������%(b�fM�Ȣ�[��d��e7�!�4�z�q��c�40?��gM��0	��Y�5�����&I4
Dq����=Sr���zîg�d�*UB���>oRo6�����s%��MD�~��Y�y�-�k�>��Q��&:��0��4�߯�)Z����q�j9�ɖȚ%���Ow.Z7��B��u��)��'�"<��~�WIՓ����2�#�a0�q�.|�?$�wÂ4K*ʓ&!�7B�.�f=��BEE��CY������s�R�Yc���z��w��[I/���sMH����(Vi���薘d[Z.��$�C�Y8�]����|4�n�*��|�r��s%���7���24̚���5�4y�
(j
F��@���w]���������|��A�����f�i�s��򜵄F��Z�����M	O��vHwA�Q�SHIŷ�d��m֤f��s�gEJG�r)���v�1&���+^�k."W�(��f�LK���%���⼋��NtS��ۑ���5��~n�r��y5�g�J�^BF�Z���r�FkZ?\�@�=:@���ö^�.�x[�3.���I3�|�DMw2�rk"���	�D��04�)�%�R���~
��MC7�+D��z���[l��u�gH��V\�:f#	}����b�_V�J��%�̀�N��)���m&*U��T+[.6�5yM���T|���"�˫=Q<�%��صj�?�3�?1:�Ej��Ǚ�Лg¥�֘c���Oe�����l��Kw9k����Ԗ�m��&C���/y�
�֓�%KeX�`����Û|��0C����6���8���"g��_��?Er��ӎ�6�l��<4�XP2z_����+���f<��P�~���Y��lc/����)��d#�|=z	M?S���}�ļr�-��rg g�S�(C`w����ψЀ̳f���*���$��6��bT�H�*�����G�7�D/���k�sqalQ�S@&��A��v��?��%�+���Ի}���T�u,����5/�78�v ]ڇ��	�� �X��Z�k�Rr&�ˢ��I��at���t���z�S��5^C�C�4�d�Lv��*��賴���Pv)����Z���=?V�vxON]^��Af���u�{o�֪Ȇ9�,Τ����t����dX����,|�Xď����3�r�)��X�*�M�O�ɮ�wټ���_�������Sr�N��Nܩ��!�5N���1Fy"�P�zoiM��>5���Z�(��2us
e����v� �ے+��|W���z͢�H�!�)����L�>�OJR�!�zb>���ءz�i�rZ�n�2�i Ž��F�2B���t�7����?�a�	I��DaY\�����̇�W:hHPp���!s���'��.�
:	���N=T�}�gk���v!�F�қ7pz�9H(�Kb�D���{�zHƬ$�|z�}7C�H�&Zj�$�$C�SE7T���i�yxt64�*�X'��^��Y8Ž�?TM�^FѢ%Xg��/[���r��5IxLJ^ʕ�%�?��P�_���a�a���%
f�4���>��b������<��"�~N�(~�VF�<����m���F�S�"޽!�uY�'�Aq��Ɨ,�XO���Zi�f�t��{GK��Die��7�=���"��<���{���JeF�����$�v�?�2�~R"�s$��کa�>�bM�c'������f��7P�ㄳ�ӫ��F�U� ���2��Ԝ��2����NM��W�n�8�5�V5��u]�~ú��1H��\Eq���TF@�b�w�
a6;M0���å���)JvPbR{��?Ç��*0����jw	+]m���IcU�2י>B��=�^k*�'�ޝb�
��������B�6�)zU���DՐlNh{�D`�'e���!�lwǤg�q����h5*b�<�y�Y+;4A�H��J�+5&�8�7���j4��L���B��HjǋR��KM�����ɻ�Q�k!�ּ2��c6���L���_w��*H�O�Yl)�}
R�����ͬZ�ek2>�{�9E\�?�u�8�'o�@�:���!Zu/���%$m�Լ_|�l?�=2+fͥ��xw�kFCKaS��Xo�S��T��:�ᛗ'I�AP[�O$����DD�2&���T�t~�$�������5=�����a��:��G������J�34�W�D�;��)�Bv���E����D[4����w�Tm΅��J����u_e�Yb��Q6�)5�<�<����嘄ŷ��������K`�09�Z�%*�'*ڌ1zw���7��+b)���IlDx��?��>X��LH��i�X�[y\eE�:7@%
��%����� �ϸ��:+����C�>1?®��A�{���I"}ʇ�i�[y>Cv��&F�#�	C$�z��%GuJ�q���N"/�1c�������{�ioCfF�<V�ï��M�9���,�s���KG5�'}�I1����U�,���&�oc�{B�q�����Ͱ�_䙔NW��m�N�407p>��OU3uÚcQ�%��bC��Ͻe�� މ.���wqJ�'�C�(��=��*}0(B��_��:�5�I��=�=`�n1��b�@|�����6��ӕ1F����Oُ�eC�\oa>b2�$���L�(&���>��Kc��ϣ�+T����yt�U{���C��0�?Fpgڎ�?F����|���� �� ����p�'&+��������{�x��M�me��}|7�,�]�As S�(%ֳ�0]�f��Js:��͂��.���z1�<��ߡ�%�!���#"6����vs�s���(�l6� ��R�G���%��e֝��r!�M}FB��> f��am��h2�v���~�s��;T�n�
�G�$ �F��I:nw�� ���.������E|W/�Rx!�?|��yc��0Bp���ڲ��o����''��F���w�AG�L{4|��R�_�>�@GVA.�;{���K�}��	�F�{�H�q�EsasUnخT��W�rX�	4ݼ�[v��u2zX�����FG�1u�؄|Feҗ� �[חj�Pt�]���=�~.����H:�k�v �J��5�%�L�1*�����֧y��&��qݻȒ�ߩ���2νU��<3�w@?9�e�W�,�GR��������>�]�r�,���5��W-b�Ugٮ�σ�8EQ����VLK&�v ����_J���Ħ��z��XMK��s���\p$O��+i�!=V/'�G3ĳ��	��wL�ɍx�T�B�X^�ޞ�}���8'c�=f�)�~(����f�G�{�p�'�6

c
��a#o2Ɩ��9H���^�Q:�N�.pbᩋ����Kb4�u4}©I�8XW��V�{���*R Ƕ:'F�{�0�e�����	5p�x��W��& ���G�T�+.G�4&W����OF
����i���]k#��c5�.(dP�S�w�*��E�4D.���#$���@�ͥ�KvI���$��P.C|�b�,L���r�
�xa�S�=z��9�Ԋ�u��c�F���[2�D/�&��l����cW�Mt���$��'dU���y���.&nꌍ� �"r��U�EpX������������F�~~\����گS%
��Gw({�%��1�[op�\��M	W8�\_kGCOH���ܸ�NR�]
�H���M�������w���ri�X\�ySW��Rm+2��K�ig���h/S��sw��"?�L���.|�o[��������z�gԸ�j{��37���?&-�� ��S�Z�?�`&�������F�d!��&���i�U���3��H����Q������-'t�#���
 (R!�L�P��X<����Z\� }ͷ����e¼W�Oh�1�?:
>vm�J(������Kj*UhҚC
ӟ�s�/�'����zQ6g��go'�M��X�8�Xz5�����稜F�2����=�%�Y�
Gx�G���ΐI2 �y�} x�\��'O�b���>��Sϵfv�#|�h[r��
�A2C*�N��r�S�e폂Pw4�U�r�+��.�%��-U��4�����"���- �0�)�`X�������{� Get������F��e��u�qz����Q�` MI�l+k�/�r��#��}}x�"H��L�,k_��7���Xq�0܃Q ��QMÃ���^�s����)c�1�����\D����6N>Q�0/!��G~�ᤨ�I�D���/��g�h
'���8�Р�#��ih�+�+憱sfѯB�t�2��x��ꏂH;��l�jQLV�Q2��4hv�5K�F��04�o�T0�Ѽ�W�;HG.�"&���s���K�-Տ�ףQl��w��XI]�۳N��x��":j	G�,+�y�q�#�msC���µV�3�
�x��	�hr�oqt`Z����iV��$N*�эZ���N��Ez8������h�y��������I��Y�0 �s�3�+o����e�"��0�'p����w��G�)(���l�zF�Dݪ���C�M�t5K��I�;���)K�;{�H��L��v���G�O�=pe1���.����(Zz�G{�~�o�Q)��X�'T���?ɘ��_V��.�~Z�B�O�S�b�ّ�b2TXr�� �b(?,3SG��,gv��~�EyPA�
�r�bI�c�t���k��L���("�@w�2 {5�$�"�̚_��Z��c|��`E�5	� S��<bV��9 �ב����B(`�����>hZ�|�t4~�ƹ� |��ѵ�ؚS��y�ԙHyE�Ġ�:�6v?S�-~����)+- ���+��z��.�t�î�ͱ ,h�܁���d�)nW�~ŵ��Ô)V~b�@���?%�&��d�g�����R�~�W���
G���r~��w�?#����[�����	�Ҧ]��ʶ�GvӦjU��*�~��׉�� ���.�FM[Cۆ����[�v��t���GW?�F5��C������q�-�"�oF��'��R��π�ƣ���
����
�D��n���%��C<J�2���armD��=A��	���
�优�*8��]�t�@���'�OQ� 7t�d/V�T�ݼ���P��Ĵ�� ͉��|��W,&�G�xCspX{_4d�M&Rc����?#"�r��y��T(̾(�0�1h ��R�R���O�G�YZ�}����k}8�h�@�dp¥�U� ��؆
/��d&7����ZW��[���f�^�:>��v�_�%FV�-����	���ds�;��3vƋ�8���C�����m���7GfV�KdJ��Q�h/��켴h�Óƃ2/45_C�1����4l:ڼ�.`ٌR�#����I{8s9s�1V�4kK�Ѱ��HD��D1xçwL�_�lXL�~5x�	�t;uIvs[��#oma�����wX3 �x��gGX\��@�Ȼ�M&��Xּ�m��LDZ׻����,�
J�@��Fch��OEM:��_t8՘������Umo�*��pR����j�g�ٷm�j�d���SD�8ۈ~|"����KaS����Cw�uE�;�.X�e��t ���I�X_����踎zLrtO�� s= r?.ObA��D�m��R�m��f$o��Jh"~�?Ó��s�y������Z���8�|�UQ��^	�Xv�!�Uj�T�	+H�@F�?�T��-w둱�ǲƝ�#j�k:�CKw�~d�EV`F�[RG��p��2�G0� Km2f��qM$�s��.�⡦���
��M�Ҹ5��PT�4_�PK^��L���!&�!�&
����+N!��_��d�'��Tc��s;T�f��hH�I��Q����^��WߑD3�/`C�B�u&�,x!�܅��%�(�~C����m������qAWAu��ٸ1�"h�|M�P�Yq����5�7�(�"!Iv92'e"\���X#g��Ү��%в�3M��BO�E�s�(�l�D�$۰��w>1�tH�1��Ѣ	��TH0=���vc����=a��}���\���Ooz���l ��V��+hu�W�m�g]6�1���2�YlХ����C��/��1��� �����S��Nᷭb���<�KD���K3f����0 1X�ʤ.��Һyh��g�s�k���>f�>Ϫ�]�>�&鱭l���/���~��)��	x`��0��%���sG�f�Q���˳v�c4|b"cތ�:Bю���~f�K?ЏuU����YY�g��G��d����FN�[r%�yp4ܜ�/6�s�~�������,h	p�8�sJR�\�'�J��g�e!9���39�l��L�Їe��j���A(3`�gA=�s�SQ��v���ϗ}N�&Q�z\�p=���CB��$���gP�`L��Z�[C���s���W�sjd?���4�M[6ѯ/����&�ȗ��rv�Ą�����>'@R�Y�
�
?Ս�f�is��E����;!�uz�Y�C貨�5��\$a�<�3a2ϋe�K�uQ}/C��%M�ɫ�k�Ĉ�%t:u,\�Z1�T�'����=�Н�u�=T��b@�=�ӣ�YK�2E�<U�T����ۙ���Z���Q���6@��b�k��a}]�8#������b�+�f���b���VhaT�#��WR��Ow%��t!P��%\m��Q�MW/ʥq,�N�?��~����� �Ԟq��6V�M�1�RƦ�G}���=�3��������|�Y��:����,^�����̥����_׬ߐ�d���c'��!M�s��a��{�2���E��uFX"�Ex����������(��h }B=,�`�8h��lI�2�A"='�j�ϖ�a�O�a��i�!]���9>K�h��} VxP+�l����%;+2s$uS�O
k��S�i��=^y�j	�|�U��6���c�#�	~g��D=�Kݕ<܅�;�@�U}�i#�8�+]E�q�B8(���M*���^��^$/**.����*�����.�L���9Ii(�XS%<�N�W�~���eو,���d?F�7�"s�<?2����]���:�ƿ����9�f��dj�\#
�J*�%����N�NѓHe5�B�k�� �zk��Ɏְj��R}�*ۑA����6k��u��t�s���NN]L�7��_3��_�C$a���օ���@ՓN������K�<��S:�6�P�g�ˉ�/��z]�
�_�$����ݢp�(��N�y*�Z��|5u��G�i3�+����U%^��E�ľ/\�Z��3g�/HW�a��u���V�Q�}�*��!ZL�]�U$�n�NIHO�ܺ�TH
�b��U�DCݷu��ư����q�$��������0�m� �+Mޑþz�������s�#K?!Ä�3��h�r��COgO<����14�$y?u*E��A�s�n`��mS7G��>S�F�Z�#�����V�M_�Wʌ���}D&��|���3����Iœ��C���f@`�%���G��k��9v��3�&ʂg $y�\w4��{���f�Dȉ*9Xy�"߆���cu�-�chP��M�I=q�5+�cK�Lm��@�SYG��P��ɏ9p/n�(v@��k���81,��M�z�ə�cR�Qa���+�K���T���z��!(�Ӈ�t�b嘧�dߊ��6y�1�洷�bt��!E�z�J��lR����V�0F�t��z�>��5r]^t�Z�Q�2�4���jH�����쉨�w��|�����?G'|R�tt�.�]�:��$���H�a�$����� �k]W���)FH��T��)�x�ΑN�*@����X��6J���$��������5/�Z�C���@إf�v�I��# -�c��˅ZA#|Xa�N�������Y��"I�BE�^��,E����n�w
Qa�<�'���M����khf��7��٤��lA߄�ZK��j���w��h1��?��[MK.�
��}��y����4y�zK��z���9�+��L����\2����uKU�^��xq7�(NEm��t��ƪc�ZQ�z�s��9ي������1I)ym��3�|�ʺf�i��S��;�-��zð�1	w���D�2�?X�.�T�r �%'lr�4B�{��k�~2*�&@��a{��k�P�m��I���]�_��|>�C#z��>��/@
��.�W�;C"��I�?}P,�R*9�13;��3X��&���E�*���̖�Y�.�^H�/|�A�,^�-s$�f~8�l}
\�'ΰ"P��3m���SY�*.��'��
K�<�t^�9'F��!��!Y^�+U�Ԙ,����	���z/��k�/b�����M'���M���D��/i�t��b��>¢��R|����4r�x�YN��|1���;��9Ge��~�L�mŵ��m��S}����,�+$%c�����"_L�<a�{ri�S��dL�����;C�Ɔû�L�ŹLk�{���e�$��f��ۛ�@��M�P}���T�|n66�Rҡ�0Ζ��1+��U�A&�۽���:���̿:�E���!��g"�T�P�K�}��t��� ��+���pi�������P�T�).��u������t�zM��֞a��s��	S��@8�Յ|�Ҝ�����z�sLzyBV�Z���YSgO�k���g�f�0�&=�R����<1���B�@Huj��|YG���a��������b �q������&��x��5��L���p^������ʣ
���k�`'��n��,q2k[���\O4�)���j*�V�k4p�E��t����9!.�#"��TN{��P�u.ء�"NU.�� �l$�.�[�������
�h=_��&vQ,��"{~Zï$[�N{�{�J�6�6�	��z��"E0�^��'�!�����J����	��܁�H]�C	�Aë���roP�~�4�1��)v��եY�b��(�>I�d ��l�����U$һ&Anţ~A�w��_��=*ݽ�HBS��Lyݒ�N�W�%o!T��������t!a�w�:-b�~T3eTx��@KY�}f3ɘ�E����~s�)�_��K������]2̮#��h2�[��'PY£C����G�={��3�$)2����S�!�q| �V���DFȦ��}�6U���8l?v=���r�J�:���s����|2Li�ݟǥ���JI}�*a��$ʯKI�T!��$Hc=~<o��Hr�|���_n��� /9����.�e \}]�S���uB��%%���Ŋ�Os//�+�7�`�8}�m�u�KTL)ǋ?mJ��+��kzD z�=	K:��0��K���qCZm�sq3]p3-����-�Rh�E���͝�7(a���\V��Zhm�Q�.�e�$��\'1�`�2�g�"tvF�藛�!F�H�,;𶭩%�-��kͥ����.a[|�Z]�3!���u Q�'~_+0�����X���cN�I^����s�U�U��U^�U{0k�E�U&���Z��T3&}d!Ul�Ѳy��5Z�(&�� 6:�5,\~b���1�+f��¬����\����� 7ە��{�4����ѡ��&]��hp��z�E���J�v<��G��q����Rj�O�	r��fn#�#�n1k���}�p��ɛ���ɔ���m	��Ճ��hBQ|/~����ym_'�Kz
���_�<��y�-O@�{8s1�����*��R��'L�Q����4 ����k��[G.�tM�'s��F˜�$3W�MMx���Y�N�X���C�t�L����lU�⧝���"�~=Gd�ZA=б�r�~[��m�`�|���k�-�.��qW,�����(VшׅV<���O��BF^��X�q�w���Om���ꋰ�ף/"� �d7���<���t���2b��;���/���.KЕSݏ��W�U_��J}|��Hț�+V�U/���z��9�9��?�؃��m��~K���q�E�k$7*�A[1�kk}i�"-�%��%��/H�9A4�R�E�2�*ce�|e��ʎ��>���S�_1��\Lw����R�r���x��Ul�pN/��n,�P�	�!>���0����C�������;��T��L�!\�/�����ɟ)��@��<��f*��q��[� �ɭ|��En��=r�Q.�NP�����ذ5��dY1�!���J}®A���&�ʙ�h�Wn�	���Ӝ��n�I��O��G3$�&rG�7�I*��9�H;���N�\1(s����r)[�n����fDR*+�"2{��������<5<�(����2H���X�����x�)���sZI�2��xZ���_n�SK�¥����ڨ�c�>���cȝˢ�(l~㭗r<̆�9[!�[��`�#��Ogʩf�~����[�x�,����;�����O��)�h����Cş,^����#��yY'�҅ą�����䬉��o�{p�&�5~5�~���o�R�o0�
� �N�jh����W��Z�'��eB�Y>G��%E�����7�8�}�l�SN,�AGv'��)��m;!m�RL�J@�w�H/��QU�8���rU�Ϳnd��Y.w�g�JU�� ��?���A}I�%<�pr_	5�o�WQ
d�:�_^/��<|���4V��H��m�o��x�lh�*�/�<�u��2��Z"m�v���B*�<���G�y��f���r�i�C�D�3F�荼}Sn��(:T���W�5t�DW��r���@�`e�s���-A��D��uO�Z�g�:� ��j������DF��qaD �:��i硥i��l�����6X�)���,=�G���C܎����{YY��#���{��ԔC�W}���m3j���Xe.�������'�J!��Bu����B@��UVx�Ğ����0ڼ�e��!�R/�Vk����g��K�{�+��|`�Ǿ=Ƭ���9*�������#�^M�qr�~�쀡U��N����4�E͡QW���(ܧfb� ���f�a}�b��[��C���zJ4ۆ�ὼƞ�*j~� Q%�UqG�g���<�"�-3'��w6rQ�\�zY��:H��U�Ԏ������ƣ�*`d�&�5� ��Z���=��h�>��44K7kׅ��8I�L�+}�������㘺��PqVΎ���8�?�xi)u�8`�C��-ɑ�U8�$x���y;A����*�7	��a�N�U����γ�f?�Z��Zn����٧s����0�WF>ϭP�=�Ua�gL�$���p�`�B�]|S�J�E�m!��H����t�j� �7ÿ�13zG �y}k
A:cY^���sKo�&yQg����|�RÊU	���L��d�Ȑ�T+�[	�Q"B\=i��^��a��PY�ą�������ޝ�`���{����:9-+����+`.7Mf�2<��h"�_S{X8��H�7\��JD�E#��a#��#��f�g�J� ��͡�v����KtɎ�[��`"�3@�P��O�27]
v� ־*�r�E\xH�Ғ--�w��'� b�	�@� '�8;��m����x8���a��B��i���}�5��:	�7g_��Y7��Ɓn_2[��mS="B�.V?�,���IM�65�Ӽ�E�a���P��e�Q�~d�me��j���5HiUu?�r��!�+���'4e$U/U[�1�D��;#M��K�-��a�-�qVfjf�7M܁�<�b<ju��$gJ��}�:�j���SP�:ox�ٿ��Y:a�j�X�|��������V�N"^a�����`��ۃN�Yc���E�۟��K�88�͔K6��]���_�!p��X(d�9�ȣ�H�˲�rvzA�C cS�j���G�4��^�ےO��x��������HP��.	���lU&w�5؀G)r�_��@3e���d�R�<�0J��Rzr���)#>�eQ����<i>�w����%�6��F ���y�S>���|�9I��χփޤI���6����o���ݒ�#JTBz��sT�&��+=,&��"�B�����A�C�Xz�q��F��x���t�����=5����0�ڗ Sw�צ�YW^v�XҨ)�v�����:�"i���G�����P	���z����\B/=��f��"�)���˟䖡;�\U��1,r4�F"���\�qp5�`�O��d]hiY�/�YCK��_S���X�nĥ1�]����e@��$����"�O� t.���3\S@�Q�?P�/9�F��B��~>�u��� �H�����!�w�e|Z�O���T>�T�����k(��Sr��	g�5���̴h�<D��Zk5�{^�u��F?�F��~7<���[�t�Z��Q���j+�s�6�
�|� �)�m@��gz�5Mn�_�$�+m���d�{�/ԏ��.���Sc��}���c����x�㿼A�*��s�͓kbKy���?�l���`��B�i�}���6��Y&:?�6���\q+81f��EJ�����8y���+#�#w��j����3�������R�8��<��+��9�к:��Tf�P0ͼ攻|����(�B,E=�f̌^��`���	�3����{`�:G�N3��R����T��m�1m��!�Ϟ���-�?�4d�ӑ=O��q�y�+��]?�� us�ܚ��z��J���$�k���M����A�˥dc��C��!��g�t8��ͯR�ɹ����1�u��a�tq��9�췘�s`�4AZ�ײ������.od ��i��5l}�h�r��w0Z�9;�w�ty��{�S��8��l��g��7��A��syZ9����B�*� �g�d�UP�֥�`��]N�Oy�����t�\[L���þA�w�R1�iA��z��{?���Z��44E,*�&M,� ���&x6������A,b#��tg<�F��"̆��Z��9�р���F!#Ƶ9�/U���YQ�U��ifDG���, �����eb�y��ZYĝ(9��
o!�5pI�yQ#���k��� �L(n1�G6?P�t�K�!�{���.�(!RyІ|i���nOq�8�*�#+N)���7UmEp߼�d��$X�W^�	�5%�@��A*�~-!	Y�&<��=����J����K�򊉝��in�}᱀��*dDq���Z��/#�Bѐ���R
��Q�|*�g�|�h�C��;>V��(�ա���%�L�����D3�)���DЀdIz6��ְ��:�|>�m�W��#�!2s��t��	��,`l�	�)(�J���B��U
U��u)�û��∓<�|�ȗ����Wy&(l�۷U�c� �۰l��������}�ޓ"���y�{�7ɡ���+��Ei�j>.�:���8����9�xN~��y�5zB,VIv��
w�_��z%�Y�_n����?�h�^�t�KW��
�F�Y����`v����AZ���wC�4/�7MK��@u� ��ui^��	`�����;ֹS�76��j5h�V׶R|����x5���a�wVRVV ��－�Ok�<���̂r�ݳW�[�¨��ZT�=�����B �vL3)�w��ޑ�W�GO�!�=0���]�B��_�/?��0�Sg�d��I0�Bj~ks�P�e*Ά��0%�"�Gvzg~���n^��/i޸��o�):I���H�:]o���k�2���A%P0���W�Ȯ����/�`<��ѐ)�|��-@�,����9�β�6p�)	hWo�=Ӄ�A�mڗ!io���C��1�DNf��Zz��Dkl���]f,����!����+���ej���tOa�U%Q2�<�'~옋��%��Ŵ�=�y����D�nk�I�B�%~`�W8�9�Ӎ!֯����C�	z��=V��i�}�;�uOo*�Đ���COz|Z.Ʈa��ς��A5v���D_�_x����Ak0�8��7�n��v�̶��Y���Pr�y3ߤL�Ps�J��9Wd�K�C�<3<�sT����*Q��7 Z$*��6��L?7���jǆ�`�5�����Q�}Cj��ѼWg�O��pC��g�tG
o���>h��sD��2-K+�h���K%^`J�����M�4��n��p����v\2Umҗnb�����Wp|��;GF�������^�ݎ�\��ɴ{�ȹ�7��>Mն�J,K��FB��#�(�+C�x���j�����j��n-��o�=EZ�*�f���(�0x�Z���\C�5���٧%Q"��/an���8��<j�0<���H{����$����9��(X6��>��l���+i�(�Ɍ9'&�� :.s����2�c�X(���\�މ']�Y��Z�qׁ�����֎[c���8˫h�8�� ԼM����Yy^\o5�� 
�!'�E���?/4��A��0�����F�aɰ��Ҥ����l��+�!&7���˟ Ic�
BK X��-��Wu��b1��[�JI�������/�S�+IpgcJ��� ��b�e.���W�Y���ae 1L֩,B%��H��_�y�v|�e�|�EsZͪ��.��=�3u{7����aW�gb?��J�u���)�u�;�Q�r���y��k�,nq�T��v�����-�!��.��UP�wx ��tS? +չ��-��n
*�OB2AI(��;�K�V�8;>iMbo���^ ����n5G'd�:Y���'�l�tW^$��r�E���ӵ�%�|��^�M�H�^^y=a.m�>�ft�X�1�h<, N��*�1��Ro6J��=�{�5g������[�0U�t�<	�/ǽ ����Jr[p��B��>��#�P�ȷ\�ܴڊ�-^eR�9�؉6SZ@�ݝct8hє�s9�0�≧֥Ȃ����[Sf��;�j�{��%����U3��C7=[�;܏)�:�G�nl��+�TT�����[7ؒ_���
(J�{�v���݌�b�<y���l�9g_���_#��zEF��DT%�vf��|��	��u$������-s����\s�CQ M��%�PEm�]i�p�$~���
�
f1�^�W/�\��p\���a���A �:r@�M���؍�|�u+H���n��l�/�m�&c�6,;��t�ݘ�� �b�o>���P��d��Lu�W��!YZY/J^KQu�E���H��Jr8=�Ɇ́���t�\v��`��|T=���'&�q�>X�ݝ�4�X5UO��Tܕ�vw�M�g �� 2͈/Zb���F�Y��T,>r�v3�+�>`���?�"D�V5������������ᔟ������B4c�A�v�ud��PO�0�vD�$�~-/;w
�WdtG�,=g�7t�5t�Whs��e��F�I-16�9D��ND�'��>��ѥ�����M�2O��{��a*��nEPt4���z^]��b>�l�1ym���5.��f9�h�;*b��:~�M�)�d?Ry��G�ȟ�o�G�4�E���Ll���/�!Sޖ)����*w�s��C�;�7�Q�2��t�I:���XuX-Wv�D�b���vq8N�@��� rha+�_[��N��N6Q�̧|
�xnq�N���o��<��F�BF�����B^�+s�)�՟�d��J���͖H�O���O��Ҁ76�%�9�B5'���>���wZ�y��.=�tr�ޫSW)�Ǩ����֞(p��z��z��ŝ��hs�@��
��nQ�7��d�M��ǢR�H~sԊ|J�I�vTf�Xf�H�g�h]�/�6P�$�"������]���T�}�糼��2��4z!d��Z���߬��v�#�5�p�-��8��k���R�1��~J�a`k��0/28�xւ6�0B�����r!�'_-�,�>�_���N��@v;n��NJ.P	0�.�����!�uZ�y�a���b���Z�����u�B�)��e��L�����D�ģg����n�"�h*�d�ToS�]�TG�AZ�W\��9��g�xT����eO�ɮEp��W�ZS���&yE!��i"�.�_m��X�� �L-�co��O�QKB����Ԩ�����_�JA�������J}�T�r�L3�V;m�[:�
j^��g�{a~����m;'Bo�g��cѺ�YĈ�˟p��B�D���Hu�?�A"'��B����쐥>�T���Y�p���~��ή��aS����ﺋ��){xn��2��Z�(���C2`Dױ����V~y�t�.�?��)��`�"���V+ �T�����[M�.2�l�'��~���Z�����QyO/�Z���Y�I���ϡ�l�/�n� �+����?�
!�<�&1d:�����z��*0U&�7`��!�a�wom$
QM$�,�w8�f�?��[��\��3%Q�E�h�d"�GP%�'ÝῊ/F����G�FF,"Ӈ��g<%�M��jVQ*~��c�_P������B�G�3<��Hp4^cl[C��$�4#��f�p�&[Z�aŗӎ/��4jL�e��d�Sfv��坼4��?u��l����$if�[��2L��/����}l��N=~�쯞�*ٖT*'�������1Sm�'�ʦ�`-�Ta>��4�����]N�0Hm�q���+���$'W2�YYc�a�n�nB��RV��¶�9w���	>2�J�c2�	Z�G���
ύ��E�2��^��nĦc��T3��i�_��Q^2�Co�w9𝦐rP�e�6iE�]�\S��&�qj/(���A����0(D�_����L?v�ٹ�$��e	��lӆr�3EZ���+,�Zu�Lγ~|ʾ������ �q���':|���	�G^.�r�h�$�T,�uSrP"�)SW�˭�Z�5+k�\�aЮ�{u!ǻX~F����j�O���M&�H��q�U�Z�7�͙�c���uZ�հ���=_���$��QG�z$R��ؕs���y�r�Mŗ��%�s�Ax8�g��6_U>�s��¶D��(���N�z0?��6�gmG�M�̃=��d. ��f��5���b�>�|�=�b͆��ˋ��,�}�Z��K�D�辫�zY�� k���5�a$�Y�/|�/n $�[L���,P���u8FV��Ub6w��.�G$��b��y!��85�V���\iM��N"C}f��-���V>"�D(B{zP�
%�V���?ۈ0������#��u��(� ����D����q�*�?!�s�%?��W	�Y����������ٺ�]���ʳ�ex�g�.���F�4n;}0�*�7�*Sv���h�·h���Җ4vE���`��S��X����A�p����KV��
�R�/P\
��D> ��fA�{��"㰰�	�Q�X?� d>ѩ�ǌ��0tfM�ē9�a	�o��6i厸:�l��Q
�X��I�6��:���0������g���/�؍4t�$vf 6b�`,����Fֲp�<�wW�DH]D?�x�]#�)�_+����e��/T��:��WSl]Zk�A7I��d�C��т�����Q�f9�x�іe�I���y���!���p��,���\��Jl	���}�n>Q?n�����X�GKGe�T��DrPgo��,�+jf}�AE��c\Lc��ۡr/�N;η�pҿ/������s����-�� Z� ����Gc6|�I>��nY9�WYʲ�2�N���Bu��tCϑ��b v���\��{�0p������+&WЈ�(J[�t-�<Ǒ���[~D�z�T�,{�g�1P3��E������iI�^<p� 2�"�e�g��N��[�ϛw��,�8M:S�q#�����D�@�/�om�l�i��i�k0���a�V;_H���mg��9/5Y�#��g���܌�ʰh%��&�X�i.��T����������C�]%���Y���(Ғu ~%���M�KG5���Va��к��K�@��0)�>T['G=�RC��Q����'4���`9�����s�6�&N$�9�6�D��?T�����o����ujq�J��ழ;.l�G��/����Ng�W��I[
fB�J�X	��k5�Ȧ��C��V��m�;�}8b�2ϩI���w{�
a6�C�t݅�ah�~5@���;�r���ԉ" ����o���O���F�����3VȾ�/����0�������5�v��G�=�@�=�]��2�H����"/��zL��1��u�F��x���S��9��@�TnEC<�Y���^��X�,2׋%��E�S�ku� F���C�=ދ��D����f�_����^uF�p�ζ���#��+��;]&�	�r$�� ��^_�� �;��D�O;2 ے��]g�a�Ͷ۾C���E�S �����Ңl�_�v�>��~�?��-����*��_���Tm<o��������%9�^^C�n�J�[�==!��"�g���嵚!@��p�/Ú2ؔ�1ڵ�r!�^�I$��w�N�	ج6���V���_�a�LfR>�䲑>:�S4�Mxc�Cy���;�U񫬐��#�Da?�+&#�q��Ȱ>��A1�����T�VI��&-��v��|��uh͆"�L�*�YS����bƳJڐ��u����̶$8:\�}��o��W�� ���?yH���\z����&@:{.lPC��C��P⊡�a�l2��� U5@f��ϡJD�J��#i�- ��q�_iL�,��c!'u5�� ʙ�κ-��k7�h1��z� ��`�ΐ�~Q�z�3{�#����S�.z7����ߨ��{��S*'I�=I�-�Y �ցGaed���3��"���������u����u؃��n��J�I�E���˘�(���q���mm��b�<h�#���T'��.�#m

�?��.���4��@�
�Y]r���.m�����3�+���]9�6 �Fu��==
�1>7f�(~$ੀ�4g3�%R�^}�x���Ui��v�a�ޯ����N��z��'3���u�,Vx�֘3�6C@3[A�g�y��%w�Wz�&i6����j+
�B��]OG�NC�"J·�"2� x�5�[u�P���أ�e,F�J����!ä��5��sj�)u�o�I*B;C@-�%�Uy�B���>P�-xw��� �r��m/�/i`ٰ�(���yTN�>�m�&i*,����U�ԓo���D#�^e\D�
�,!�Q[����w�:E��4��k�U8�"j�����!��	� ښ�� qq�k� �/9,�>�L���>��R�h��}}��q�3�E�p�� ���&�}�l���m�m���@�������mW����`ed��86O��-:j];\z�v������b�D�)��զN����k�K��P}�&�[��a�o��|��Z��n���Q�Y�������rvG�l*ȍ��W
4�	L���6F�bpyμ�r�.Z�x�9Yu�Լ�.�,��񝿑_�lE	��:rB�l/�x��0��Rgk���7~F8�~�:���;}�?���5������'���W�Ʃ�X��2Q�:Yt���uQ�/�s�'gedB����o�]<���h'O�Z�bc:xy�WO����%���(Q�TH-'�n��b���4x�,���m
9L��]�i�Q��a#ƞ&iȄ..�L��!!*��{pA�r�2������Qra_��������6���ͳ���g�94(WR ٍl��D��E�ט�,�	��z�bV���I���*�ڥ],v�CS��7-@��\aΐ�|w�y���D��G����-����_n����J.
Y������Ie\0I0w&��9Y=M&���*,BR�P��,�HN���]�A�[�|��N ��S֢'�ˉ����t�����ɯ��A�	�4PQ ��s���z��`�M�vsJp��q2)fp�K�Z�f����q��S3��Y!��>�*�PX��LvW���B��%>g�]h��a�-j\j�ɻ����� E�)0`���n�:ѡr'I)��]��I� Lwy!<�6���sa6�f����l9�	� sh��7�d@���2o���h�+1º����1�k���:60��Y��j!���.e�B��&����@�]C�8��ba�h_��Pba�{E��m����'*�y��5�(��}�74��W�|����l�f�u��7l��Ԏ�x�̊������`ഔ��g� �K;V�]D���E�d�ח���w�:a��Ӈ@q�(�=P�Nd�k��6	n�+4AXM�/�����L7���N�g#cH�1���5k�YkZ �z�֠��S	�:�'�$8(�)�"L�J�c��U�ř9�KǙG_!؎Ǉ#������}Y��ƨ�B�E~8'z`�خN8�m�����X!y��#�i�;������'i\]�Ϟ��$O���`�fz�g|i�6����
���V��\��d�A*J����hjaV艻y��
���KUn��&m�r��Z1;?��㵾٭����{;4��|B�G��'5�rkX*�ǿ�vu��Q��x!����|Q���	�#Pa"� �f������b���.`tA*���qLvgz?�2X��JE���ϊ�*)��Hx�����ƚ]H_%�2M�>�������6�VZ4�%��u`���]����u�p�?���N�����7�3�=ބR�=��,���u��4!m�񣱘�­��̭�u�6���{G��PerA�q�|%�#�g�2
]�h���t��"vԎ��y¹�2a{�\�U$՚�L�A,;1��Ϙ}�ܹy��� ��fIq���mqX�d���n��|_������cy��Nu?��{�q��r�\�x�^�\¿���j���p
��,�[�~1Q��k���x?km[����W��3@�������\@L�J�d#6b��;tQX[i�Ukk<����~��y���&dL��+,^^�Z��"�_�C�o�o��V�b��d =���xm�]�<��pz���h�� �wCT�j!�n��Z(�%�֓�U��W��7+��*�w�X�Lǝ\\wY�=�G��v�gSly���Yz��g�I^==�BL�I�3|z"cMx��ɍ)�|l�N�D�D�(7_�#^_� g�s|�e�x��2��M��q���j�t��
�6g�}��+���̥�^�J?E�X��z
��|ey�b#�L�
�C������:���5F9ؕH��,�ܯv����>u������&��	1mj;�*�Ԣ����t৐x�:I� ��'J�XL�r8uz`���׌rZJ��Γ������5��p�v>xtY�\v��9|(UV�]A��s��#{��a��T_�Y1����Y��a��0`��m�+e>ҁm����pǽ�d6]�� ��_aѷ57aV��[h\������!�X�!pxa�nC�\��_���T7��`�q?}8�!���;m����93հ�O(a���l�������r3��l+��w�>ۄ~򢩚L(�H���P#r C�k��;y7E���ٚVD�lNt	�_D���0ֳ��1���.���{�<V���χ�
���D;,�
IªǱP8�z����4G�GN�|�#�9{�F+��"�3��P��X��Zf�q!fSM�=�*8�y��h��Eʜ2��-���tV����:
���$��Y�,G�Q?���7�E6�Wh��^f�d���)%U����8Vf��Fxv�'��g�!#�4h�3�A�<M?+3���#ݼɺ�K�z�۶]4-���)��FK�ʁ�*{&�*�ݒS�h��|oU�Ce�v�7�� ��Za,O������2��`�Pw�����<��a3��6�g5;�R��	%��{�����M~C\���ڽ��.�"�z���Nh���NOsyЉ�
;T�dܱT�T����I��r[�i��g��m��sa��fH5�FD��v���?]�ƽ���t���q@�*CɫT�;�ѿ�9�=ƭF�śF��~���5L�����.[h 2�@�f������U<�^x�Υ��ڒ�X�O�Ơ4l+f�@f-r��/a���k���FZ��iUf�F���0�}��Z)4�^�rsۙ��L�TU�n������M=��F8i�������pVe�3���HHv��Q�W��Ǎp��F5���l��p��W�0o��(ݲN��:�NhU��[���[�>�o�hc�'�"%���Aqţ��7�t<�
q�m<l�1�(���byL$�4�!����Lv:��3'���\E`�8�9�w�h�#�a:��{ECP�D=�`�r'�r_���-$Q�'�n�n�.l7��Ƽ8ӟ��a��ǘW]���6�:3�j�����xr��	C.�w��{jY�i���3�<6�	���2�T���2,'ޞ!f�
Z�6��M�#������m"�xY�:O�S�Z Q��M<]�sK�n�,K���7�f@5+X�<شת=�2�W9�����eVϧ��E��Ԋ&d�G>@Z�2SO�T��[ʔ��F����tc�lg�����N=Uq��t����~��O0J(@i'V�M�����}֋<3�v
P�Нa��\��a�z)�������^A���O�_�@U'R�/�I�P��e雮y*y�b�ӿ��%r��AݢT�L�3:V������d�;��A��Qz�Ȱ!:�^*8��F�پ�Ζx����,�<vb���Y�,nĎ��HzfDt�5|Q9[�4�R"F�|�>k�yT�R�� ,���R�a�ۋgU1��5t�9סdy���+��/���W	[���$��L�Ⱥ�"�A�,-��+�`� db-�B!���b�����E�V
��X0��y�et��������,U����׻�$�|��<�`�@�i��6��E>L�57h��� iଳmf�'gE_��'W��妚^�ng�D2���1�Dgo(q�Q��]��L�UX��R�L�	}�>ۇA�-�b��Ab�c	�꜄������3?q�G�ꈨ)��ռz��vf��~�,=��#��= �:�**��o��:Z��Ac|�Z;|�h�w�cӈ���0-_�R���j��-.өw��ǔ�p��7	�I;2�^����ی ��E� I	0��Q��~�0:��pΣ�ShyD������Tސ��������%��� H��`�B��Q��I`P�c�v-��}��%uH�,�#Äa~�f�Q?��q�B��ɓ��V���O1#�3������m� ���ܪ�M��v��<�Fޝ0�&d�!�Cb%Y��d\�~�Ra�1�mҿ;��D�krx�Eכ�7�8���Q_z��o�k�,]���5�o�q�k�O�.pZ;����� �_�d7,i�+�^�\�' �WS	����-�WA\?d����j0���0$�USmf�c����Y)�v������!�f*A���ixu�Z��&���%=��4N��\U� >��3�u�k�'9������>w�ø�7VX7��m*��<#����]JK��t�|��E�in3��$@���"*���S+�<.b�O�~@N>/��oc��Cj!��Z��jz�6�?5ìO��)t���q�	`K]O��.��[���寰��u��$���c�k��_P&u�b� %�gQÓd�K%���������M���P�Ř+d����F�[4�BFrW*�Q��8~��<4�L��%F�������2��λ �<�F��!*����{��>^lݟ3���4���i��=�I����cR��L�9	3]Y�l�J�(���h�G�C�ɶ���n��R��Y�d�E������G�Uϟ�v�g'�$	Q&����*���O��E��}�p���0�`�a�L��
;���M�$�����h����w�����(!�g�g�� ���i�K ��U�Ȥ���7�/���Ӊol���h��2e�W~S+Km`�������ɦª{Jv��@8�N��v�U'��G��fq;�|�65o(�c�?��W=4�
s{�ٓ��B�?���>�r���Ō�d��S1�K��&S�^-x�$�7�Ej�7�&~����EXo7%�;����j���(h^���ꎟ��b�?�ѭ���xݜ�#>�w4+����O�0���3Ȥ����^�E����4�Z�$;�����p̬�Pg̴���)��;�� �43�_��Cl�cH�*�u%/N�
T��������UF�"X�dԷOQ�3X�8uZ1�>39������o���x����y�������#���\�����yi���^j�{��*m\E�	W�Z^ψ�W����w��Xܪ��p~e#m�Ve�3��:|���wIkv��?O��ԣiR�ΥF9՟��Q��YM�,J�?j��B.���,����,��J�� �4'�^�%߀*����)u̟�O =i <��~��73P��_�ϙ�˅ѻ����n�t��A���,�K�cD!}��ލ.�Ӭ�Ȗ�8^si6n��Yf�J���潔�"Ѕ�����_S/,Ċv``��e��i7�m��D�G�vXn��F�i�e��xH/c&��Z%���P�&�a�	�?�o/����䥿�'i0|bկTx�qtO�4[du�����5{�2aF��q�[҃���W�"f��U���L��$e�EI��P�V��1fJ˵g!3c�}�莊��9�U��$���=��H�h$!|�Y��^~���`�;f^h��$'Y�o����"#�>�Y�Ucۇy�Hp�
��QMgJ}�v]Pb2Ő� 0H�^�)Y�����Vs�{�g�\��wL�ĺ�SH4B�h ���XS�^�9"�:f�8�j�	����&0���g,*�;�3��>�qI��&�!����z�1��,
~xYq6,r�A�.6�,��H��+x�R5n�΀���f<׬YY���S�%��
��r�h�`��Et(��]�P!K�HU<�~�A�F/\/����r*����0Vƨ�Z��J[���#N{������ga��9F���U멿�[�R�h%�'ilq�k��N$Ϭ��p��G��� �9ؘ�.��}��;�^�.���m�U��bAtL�)���F>ؖ_M:�nl�p
>"{��3L���2�+��3O~��HU�����1�
v���::D�����F:���1z(	˫������$�����B�.���r��s�p�k�MD/?��ꆽa'[}�m�یK���\6� Ygi�����s�hiفl�5�j�	�Z��Ӻ��'9�2~��zr4wkו̢ѵ�6=����KWPs�[��2�J�<�!�X��7���n���,���l�և��i'ܮ���5��U��qJ�}?�GS��DEZ�R�𺏀	�߸y��"�Y$��V�CT]
��n?��l2��{W�\��q��.�0?g��[�C�W��V��*�;�
W��e��*�D:H������Y��_n��D�~r�����[�>����	��DzW�#����v	`g�<�,�V�? ��و���aF��
��O��g�?�A�F��a���W��ac{_��O_0A�h|���
�q�` l��*�-7�<��)Te�-��Yy���us��m��?��gj|ɔX��i�Y�q�t.f]ǯS�G3��KC2fJ[�`�E�`�x�m��wH��FF�i~����K�&�c��#<��С�u6�L�L�u�]]�\e��3�_��CT�%�PЉQ>X)�YIV�,��%k��%D����33P�-"d���h{~rF���_�/��*��/ww���m�~�{��I#W2�U��?��@����9�f$h'r���PE�(�&Z!")������H�+��q�b�e
6���S��å>���+	n�V�t�0'�7�ϟ�l��.�����w��ulݤ#�ؙl����w��{�]�F^�|��&��UQ��,�r����D���,y��Pk觟��I�0�%s�4�>���=�#S�s(���(���{��^Z�+�>�ҝgʍqd���e�
��=�0���Wv��3�&��/ս��ajl��en4` 0B�,��@��������ݗ����L~�0^�Xbu��?Rۛz��MD���^�t�ճ��g<,.|�{�L�7v8}�}ijm�f켹0�U��@�P�G�0�6|\
(PP��Z �$'^�¬��q��c�ᡆi4�N�,�A�/O�^˵PF���g��&�#!Ho�̀��@��#4��Tո��Ez��	&��=�`#+ � t�h�ݭ(�eT����''[�j��@�p�MQ���.7T0���i�Ơ�ɂYBUxaω���C�yw5���� V��򤪅����J;!Ɨ�j`*�����H���͗�o�n��H�H"��#B
��[J�����~�؍�w���h���t��̅�Dms�;#���j��|�S�;��>�E� ��+,��vNEL����"���+҅�n�7�Dg|�K���z7`4_B���X�T�*��=v�3,G�=�r[��1Ͱ�i���}� �RI�)K��������i��(�b~�H1d$��g-�2��ɝG�$�/<��U�z����C�6�VS��v����+��� ������b#���s��J|�k���l:=͡olf(�`7�-�]��3��Zdw�!P��̧���$�˗mb��So��7g�. Hf؇ϞF��9�0: �L2�,� A�"���&�5�B�~�T��E�<��nu���1[�\�������a��嬷Q���Zã��Ư�Z��i&�[��A�����"����O���������o�l,��"�
����l����j�+��ډ�ý��%�d�U4 n)������z�IJ�i`�)n[�%��_��s�T�f`��-�����6$@�!�sZ�1;�N�xf�N�s�)�D8��Z��x��F� ���d��t�9�~�+2N[ y�X�~F��[%����.�Yx�f)yP�\e��l�2��iM�M:��P�=~d�e� ���C����w�$JRu��� �;���e�AǍz�ѧjbf�ӱs�oT�>_$�}�cfF1F;۫�]�Tg]��?�\X��Hxx�&�nn�gJ5�%?�x`����P�H嵿?D݆{�/�H2d������ݛ;8S�D�����w	W;��m{�U��/I�������?^��;��o�çќ%n��K2��r�.E�ɥ �ؼ�k|���mJ ё�2F!"��o�I�p@��GO>�v������SL�I�_��yr�����6f��t�L��\=������)d�v�_�hU9T� kn4��j-,:I�4�d�(9�����e����M�)��Ux/͐[O;La�y�7-J�ÿX����I(ah�*���Ϭ[s�(���Q�������T�S{q�%t�G���.ؠ������+�t��=�z���IO�Q�z��X�u�-�\����^���E���o���������ס�4��ш�菜I��R��E�x�ASE_j<6Ä��ֹi��h�:/(��ʅ+���ÅI��s����a���PI�S���{��$I�
9���jۅ�����x�6�W�WJ��9ɖҸk��b~��Li��Jf�y�_a���E߀�RuӃ�:�'�g��Z�$�oZS��fee���( �+/Ӎ�7@{g�ˁg�g�׈V~s��ܟ����o@r�M� ?z��E�zk����1XY��(�<���<'=ƹ)+1��r�8!Z(wF��I�Qj�OD��H-����䪒[��(�F�x���"v�K������B,��J�H"�v���aBOtS�t*{]�Q�	���
q�?R53�4�<X�b%�����VM�c
��@�f����y�)DNF��M-��'��tޚk
 �B(qa���6<ֶ��}S�R�;<�L2�Rڑ�x���TL;ر�z����� !���_'�T�!��ɿ�yB�cvn?������ 2�rK@���5���oܐ�(���K9K�r��|���a��͕�����`�=I���,UؔR�b�)�_`4�hGgQ�-�L��Sɪu�ͯ����hk�F���L�F�KF�W&��I8�$J|ߧu	l�ϕ� =�3�^�L���0��[�F��Y�1lR�Ro���aBD���vK��?P�d���,�|��_\'�w�]�V���ܓ(���H�Z��}�o����������l�L�GΗ~l�+[
���c����M�|�֊,��Xg��\�nJ�^�d]��8>ΌlY��tS��T_�-�*޿��� ����5�vO������Lm8�� O
f�+��Z$#�_'�㸻<�I�YQ*�de4R�3Y$e�x�j��p�|��Q!%r;�|cV�c�2_�{��
��ߪ��oh��t�U<D0j����o���O?��7���6o'�N���%GġO�XJ��SZ�F�v�`�jw�����kH�[=�r1�PcNr�#�Ha���i� ��(H;����Ϸ�f���)Ў�5d��.��@���8kɂ+��LS����{����7$���&W�b���
��j����� Q8��qz8����r%(�>���ѷf{������W]8,�m�io���b4|�=pE'���yX�}�����(�3EO{���9�<�@���7hWc�}j��m���n��^�9w�o�����ދ+�$�ܡX!Ek��%������c��CO�b/���yN�X��4yI��ɧS���0Z�FeG�-<xP�7VM��`h�fd�����N��D�N�1	.�@Q�������Q�pQ,f�=X�L0�-1��e6�$�]��a�;>9��&\I�������W4��?L�|��c�,EB�!eCf��AL4�H�z7��$6�~h@w�2��N��6Ix��/C�,���H#��u�4��i"�cct�;�ϥ,�eX�QֱP����Ĥ�4�6V����@:�Z�9TuI<%�=^�U��ó�S�T�5?��ȧ))_�!���u�.���ܒ�����?y�)���<4�l����Q��ߟ�����Ẽ��s��X�k�B���j#9�j�qB�{�қ5�������8�{�=Y�a�2!��(�H���~�jOh��5]�̫*w����B��5!�دFъ���������F�|�i��G�Ģ�D=�� ��o��p{{جu�{֋�xg��>�)�܃{�
8)������&)��C��H[�l���{�*���@ ���&�JR��(���n�&�����3�j� X5��&e.[�h��΅�P�ј>~~�QH��G��ob�d������a�Ϝ��6��O �������QI���d��.�-����KE�:���s��m���(�Zޠ��1P?��(zu5 Y2��$2�̈	%8b��B�K����#���W3E	�e�4^�\��0M�;Ea��K�ܛԦ�W�8	�����ciB�.��q���0~4�t!��e8����E�Q�qL�%���+T�򌽩��A~�"��=�O���&~��[�>�ՃU7��z\\�W���xP��X��QMI.�i�jvx�c;���v���N�Ѿ誒��$��n����||K��1���
�X���8��ī�Kj�*j���r��Ogh�F9lR@��s��GR�^uh�؜3e
�ͥ�f�0�N�qE�b3���X��\�� ��_v�_yH7���8_��3n��+t��7�sg���hB��P]�H���%�s`zc���ݟ)8MJ�����M��׫�u���e�֞�p�K��Ge����\�O� ��"�5qhLqK���a��L0  п��&w?͖���ӂ��}&��B��W_w���XZ��
�Ɔ89���^F��S�I!\���(
ɾ��4���$6�� t�����4��g�a#�Z���@��?��I��@riX,ܡ�'Bz�M��Z"�R09����9�ԉX���k�<��jʾ9V�/���c��T�dN�c=b�_^�= aWg[`��3YJ(�;1�䄣��a����s�"٘+wi�Ոv�ml�aZ���O�P����ؔd����
^�X�G��w:x�}?0��HT�.����޼J L�ո����h�;8p>�R!v����5�-(��6n���.�D�}_�%�s
=p�g�ٔ�JTa>UqLm?�8 (+�L�4Ǘ�o�zĊj�R��Z?ե�&R���]�b��;M�%*xj�X&~M��C��N]��2cI�r)��!8����P}��}��I����_�����cTV�_� ��V�ʿӻ~S�ev����,Z;CDM8l��
�R�՘n�������*��ے�
JA��g����|u꼮��'�!�� Y�Oa�l�>nX��)����A�C�7z���A��>�uzcTӋ��}�L��QB�&���|���4�A� �v��ū�F�1�wl�1>Z�gF����2�6A���3�R(F���n|D��9�r��6a�H��L~�Dh�ǩ�xZ���K&D7��ͳ`˼#7V��H.�3Ok�
~��$�,�r�[~�m��1O�p��_jWRH������弅W?Ϗ(k<�;��L��Ǆ=�.=~VK��^�3������ڏ9�YRSjj,=��\���x>̉������/h�S��B�.?`�8�6)�O�|Nzѝb��L��� z_6dP���;����K�gb1&�׷���%���Ŕ8�����-YC#�ɨ�U�ʲA� jR��g\���6��#N�z�8k�|Fk�a0��=ڪ"b��vǩ`˒F���ŉ��u$�9&V_�~	��g	C�����1��?��0�Od��R ��?�XƦʛ�:;#�}��u�;աܷ�H$�U��F��Lg0�H���*��ѮG5�A���~6W�p�m��z,� {~,��5�M`����qi�\7� �뱸3��"��
����wCg���=4�5C��6^����r�f�/���6��ߒ�ܮ��G7��P9̝�;�U�;���u#�f�]qc���=�	w���Xb�۶�!`&�-��!�9>�Ò��"��M��7'�>H�Y��DUŜ�������J�� �&2����S�4 f��Cms���D��ą�_��[ԅ��]BY��_P������1#�%s-��DÂ��xE25��ⱽd�p� +b���&3��}�z>�ٳ��9�D��X'/���3�%WHk���K����w<�{#�s{U7�Y�R�4��f:�jpV�4�ΟM����aV�/^a���\�����p�R��5!�YQ�8qϼwVnм�ԃ�j�]����0�y`����)n�|4ZH����q[�^;a�|r�����L�z#��v��*��{XI����T�L����5��j54ԯ���yNX��L�����g���gћ[#��E��yEb{'#�뽲f�{�5�ߑ$C�;��l�$��_�0t�-@=���z���.�R�>w��G���� -?��iX��������$���A�.~{΃�U���ݗ�ucѱ(dH��P=���A��'��=֬q�҂�d1�UIA�j�=�f�p���EJ�{�\xA!�qt��Q�yx<:kzgşk{ryc#�S�U�lCy�{�?b�ڕ9L�u���q�eX��鏗X��7=�+I�;�c��+Յ�<���	��;\�����"��y��o���[��)�k����Ԣ~q��U��/����|�jǶ�v����33�v�$:Cp"K�&Fzl~��z��xG���������5�D��}K��#؄��e�j�̰�*�������k��4Ȋ�>Z����]'���i�6!���T�$μm�ӵ�K�qi%����1i��e�B�p��m���ܺ��!jZ�=Y
ُ�����Γ/�{�[���E�����TJf��
@�����j�m�|>��>�m�j��A�0Ұ_%�x�jFZ�),��u���Ь�3�>$<�<��qM�� E��nd3��|���C��&�î����9����a�EOs^�iH8�Yƹf���}�� m�b��3q<�\�7{���R�0�.$��k(�t�{�IXF�$-p6SS�\0*qՀ)�%&�&5 ٿ�}��ύU�K�H�R"��mL<k�����v�O���ۧݩ��$�i^(y�B�諝���]y6� Bw�J�z�d�- W�^W�D=Kʃ(������k���4�����D��&|Tôz�|p6- H�{^]v�6o"�?(��+��2�T1�kр��*Қ��;f~�Ȧ�T{�H��4�4^�����\E��+#l��HQ���ݫ���X��ꤼ>fHo~ �Ds�J=���۸�y�-�c�鵅���7�7s�2?�ќo��m�Հ�T����6�nQ0�k��֠��s��&�Z���̒�%[Pks*��O�f�c��Y3h�%8NW���.�&������-�p���������wr�p�P8ʣ�K��_:v��z��\ޟ���e�%��zܢk�g��=��n��5�HE
��.1�Rڽ�`��'���|r�^��?���ffJ�>�	2���3�j���2zΉ(zm�0G��]"<�U���r�'�BvhWL������Wgcg�[�R/Vꝋ���+�AK��B$��bUw #2�}r��2�.�?��@Fu�q!��?����T���~W�n
�U�Kͭ~��z�~�BAH�.�����+�
t*�����X���ڰk����j�8A�!I�i+�ǡ��=��)I�ujN����A)h���t���u�x�����!Q�o4YY�;J��P�7�H�t.h����Ti�pE�A��\�n���GN�K �m�8��v��Oa��x��~�]�T��+���$Ϛx�;מ�-#.k.~�͒�ۊGü�ٌ��z0t"%a�$.&���!�1C-��#���=M�ck�M��Bv�we��6{�ǧ�yΈ?���M�h��ȁ� f����Sk�x�k�&^^
j��uG	���՝����]�:�{LP�g��sS��3"�]�V_�B>s�Oo��+g�{q�2n�}BrwՑh�e}@9�Y��<��NmLa��Js)��x����!�C�E�-��<�%��@F�� ݸ�
|K7M�U*#?b_�B�lm�X��?�fH�Rr�7��A'R8�����j:v d̈́ Ug;�[�
6~Z���%��֋6�f�~-yw��o�{��-g�����RI�D��~Ɍ��0��v:��UpW�is�	�4�����,��ur��T��1>=���4��%ӳ��}�UL�WPK�e�~�C0���b��˚
M�6��0
N``�y���*,�5��HqK�;��W7G!����V�@�N<�����%W�Ry��=��-aY���	�ˆ �onBy���������%d��ܿ��вQ�����շ���_��kgx$�I�Q��5B<�Z�ث�\߲��_�ͭ��z�08+��a䍼(������U"] aHb�2�� '��n�e��%=2%,�T ��I!-�!2B���^��PvP���X3Q�� �M5�F,�r|+(��ݘ6���bWsQ�!���U��U���A�0dj��|4���q%��@�����^(�Aȿ}��zL�ۅ������B��a_z�l��+:u>"��)&tӲtT/>��-����P�]�%8�*t�Q?���θcjHo7�[d�GF �z��S�@�O�(h��w��jhZ��mem���ٌ�����`���$LdX*+�\��6㱒Pe�kP�x2���-��UF��Z�����_��n�g�R.�P�ф�'�����W^:!�A|<��Ow�^Z��/� P�v���ݰ��I����
m��p���j����&��o mI�/���D�<�eKe��+gw�s�|&�.�;⏨x~W���lW6]g��{n�k����1�;F�]Rp%���r�5�.��J�A~!�]H1$�'G
����` ��b]^)j�y�	�|�1Z@�r}�K;�j�-�V�E|]������#&��5�z��{}����PP<���p(��A�'���)���jx|(�{���T�.��KZS%��D�&� ���w+�3J����X�����39�$n�}���^���E���U�HYY��#��^�u@��V��AgN�^�r���w� �;)�pX�-@��[]�TP���,�:���3ޞ�1a �D�f�ۘ�D�o/|3�O)Qo]�2PC���
��x��f�gAs���
q��9�#��� ��<uJ"��5Z\`���~3����O[��~K�[�U�ƈ��N-�Do������|�p�I����g�q�`���kZ'�Z��):��[å�;.�I��}��!�}v�u�C������ټ�풜���.\c�.�p���aUE���j����4����4~j��x�%(�����5�X�b�m{+�<�砰������C���B����J���E������J���N˲-����^y+)nOԍy2Q�H�� ��E�x��Ǉ�Mg7Rg�3'c];��]H��'��UY�7���a룆-sR�^����c�m��;�,(�yd����5J�(���B�����[��#h|gK��xu-
z/	��fQ�1����9�k�/��9���N�4�}��2�x�c�n"��e��R{~���{�ǘ�_+kW�r+�9Y!@����z��Fg)�K���m	i���.��O��_yr�ӭf�]�������نm"0Mð�M��}Ւ�̒4���|�P�m�M��Y|`��W�PC&���S�uA��MNj|���C��L~f%zݛ�1U>�������Z�:��R�5�86"�c�Iփ�}����`#x�a��*��2�ֶ���/�o�ۉ�3��9��ҹ	�&Ё�k��-Ͻ��ic˧���7�L�Ǚ�hp�aјm(�B����i�pZ�S���m�f!����!l����5*���8��b#�430�bK�,�,۫�5��d2�S���2)�!�#N+%̊��O�w;�����~Y��Z��QL��eWXP8�A�|��@�-`�:K�}L?ИǼ��;�::hS� ��>t��zV�^I��t����韢���s�E(h6�r)(Qt��p��*	��
~_o�~C��bSl�Nħ��3�]�������Bo��u��7�������2�,Ļ�\�|�llU�X��μ5��s�`��׶Ac��w5�Z�0U�k�T��ŷL�3\������A��\_��]c���2��E,�e�Qa�ģ�K.RV��X2���O��z��D��C��;T7����-�b�W�M�R8�]@�|��Ϛ�e�(Q�U�Ѻ��WFيˍ�ݤ�����L�iF���~jI�绰�94��-��#cL��,�a��py�&����ԬU�)y��,Z!�����\$T�0
1�L�X��H���M�:u��P�	����] 3G�0^�ư�@'��E����-v6�:�VA�i���p=��Gv~�=�9���"���8ؗ�����7wT�B��jϴ�׿r�3H@��~3j�l�	3�-oF7&����������"t�RC����`eԏ�`���g�m^|nw~�����_ ��6���5aG�����_�f���f��n��,��SGc�ٯ�h*OJ�N��O{ʰ\Bd7e��v�G�ēhv�j9!���ߕ�V�6����.�4���Nչ+XKq��+���z��^j+�".j��U���]�?��@��B����&]"��Bg�$�$]�Y�9!�%�wcG[��첟���N��"ÿؖ^�HjBclPFFbg�$_�l�w����%�l�Ü9s�i�R�s��"Y���]���)�s�5D�K�"����D�vxU�d�x�D6̤K� �=cP�Z�]�n�g��>�~�Ͱ��f��>,���@K���y��j,��)��ps9|�险C���=�X�;0;v��w�bU9��s\��7�vi����M�2_���Y�0�7HP�}Z�&J*`��� ^�����1�T�/��DƐ��o���2�g�E�"�wb�\���(�F�ߍ�H��un��~�NY%܎Ǉ�~I�ط�x�|�P��:��	���jw�U	1Fd�!p��3Cq�l"5N�-�����;�2E]Np��]��)$���M��`)���Tҩ��f\k��|����W�+[��[�>�̙�"�^��1�Hu�~��7�w�Q�zB"�\޻2;.������Ě�N��� ��:g,��E��uⷤ���"�%�}�`�1Ԏ.�w����U��p���S̣���I<�ٔV�z���l�|�/���j�@2v��C�A��#����\�Iz:o�O����Є�W�L#cՋ���-�!�`��5�{��!�l[ػ���
�sHäQ�H���Cj?'"����z��k����s��CT������t��@,2���q݊_�j��B�� ׅ���m� O,9����qyϹ������=�x-B�t_�`�b�%]@�ND��ߩ�qsșU���̀�/��30�ԣr*�R�3� ˧QX%z���>ȱ����yZ=�-��tC)���G�Gv�)���%�i_���0	|+�=�|��p�K�[����M^iGiJ@���{*�Fcl{��tJ����z@p,QwGܔ{���ӟߐ0x�s�/�r���;d�̒�6/���ڡ��lP�"��<̶"�8Q�]y@�� ����}X��2n��y��R�/�5�%'8ٯ�>�,x��˺}��%�P���		p\����g��)W{�ћ�5�N��֊
�����e�"����ü*p>�^Q���U+ϋ&AF�^z���+p��.s�+L&���Iֲ��_�~�����X�:o�"nrXwq��
(UE����b�f�m)ޭ�q�5b�4{�Ԉd�pZ{g��`��m��GZ7mǉql��D�p�,�f$(��w��+sP���E�.�����J�0�2��T�k��t�N�`�$��>l��N����Bf�K�*��7���l�;<��3=�%4�+���$���5���-�V7tޜV�)��b�Kk��t�,Pf�c�y�k�PH��~O�V��5�y�\�T�̘�h�BT*�}�c4��	,:����wX䦳>tw9v�ZFk=P���Bh�J��.!���	���w�ʈ`.�����5a�ᄸ$qh�!�PY���<��'�8��!�ߌS ����o�Y��d\�J���[�\�8 G^N)��;��jc�(u�����u���6�k_� 4��4��C0^�ڄoL�h%��$$�����ۭ-Pn׫<W�1̺pC9h�Q�
��1G�Ac	uŌ�h?C���h*�i��``���1�ؘ��b��|��2V��l�b���&��}Z�D��E����;�X{��@Ƶ7
��8s�C���I-o�0��e$�W�O#�a�YmF�>���C�������/F���lNJ]���S��"s�����Ip���!AU�$Ġ���w�[y'�]	���O��=nzZGcK�6���X\"��Ç�HT���.�/�%suݼWV eN���x}��oBW�)ukԞ����6���f��>�ύa~-1������ �%3�?��#		B��o�%}�B�|��\ i��3��W�*G�}x��6��#�r:���%������[���2�Ac�bd*�%o���m��,[O��G��w3|&x�
H��#O�ʤ�7bm���.�`?*z	X�`��+,�y�Ij�۞�����5-��|�@�)���k-(O��f�&�������U��̿��إ<a0J�"y�
�e�xTB�d�՛��&D-A�� /f�N�+8�"�`��S��ޱ)�mӘ�-��5R[i���v�kCH�p�c��J8��h��'��%gF﮺��oMڐxhd0y����W�)������A�I ��K�0Ī�cl��<�G�*eiEOa�MBN?�ٞbR$WEhj����I�*E]�U_��,Û��e��̽��@y�w�*q�����Ƀ̦�1l]l��y�$> �v��	q1e4�b	��:}�
e�_��7u�a����#��b'm _ r��[��m�]�)M�>�m�����GP�>�w���䅤`�����ɟTJ��1��[����p�:��*Tͧ�WK��z�_�rT�Lf�+�kD�V�>i�1����r&Ev��zM�t�$~�R���*�,�`��y\�/��9Ӧ�Aۼ�G��#���s��	#�7C�}7n�� ɾ�2ș<Av,�����;)��!5�纂2&�@��/� (R]ysp�����nu�sA�4�����_�.B�nIL�!Kh����"�r�C�ˬ��w�J����ܔ�I�ƹ6e��!�@����-��n�j\��<�q@�8��4~;Cb��6+�d�����pP(���%�G���������7K%�7'�c�%��xG� خ��7|-x��0v����B��%P�~9p���n�1.9(�\h"#F���r5K���.N�Y��;��4LM%D$s6���ǼI��t�|h>Zt�@����TgH����:F��+���(���뉋8ژ�<U��К29��_�N$7��la����r�Fb+�C��*�ct�/Uu��iV��%z,��Fr���΃�x��Gp�(��B.�S�I���V:��Q١�0�^�|Ľ���5O#a�i�V�lg�$�t�vd�0ڳ�ҧ��B0ܱN�9P�$̠�j���Ԫ�ɱ>�A�(+��^]�q�v�453\i �s���ycF)	����<�Aו�^�	S�KV�K�Ok�W�ˁL��{�S�]�h�)�Uj��I��p�q_��a�v�ܿr�:-w�;��@&T@����>����]h�`���77 �"\��n���I!=-vT��-�pۋ�۪2PN�����6�v���������^W����5f5S�T�B܇[�و�V�L���>Ҩ
sŞ��O��ED��&Xnъ	�� 6H�>�k��AᇊӀ�eu���L���f�؎5��_�zn#����������N��	���V�n�|��)>Z~��o��Y}`.ԼZ��)ل������8���hѡ�\~�4�gЮFF#V��|�Xy�����g�H��l����֔�Y�$_�v�V3���@u@u/��cP����H��cR�`jm#��%\���$�}�*�c?���k���H6�'�����TX�>bNE����;$E��_o���`�P�)Y��W�W��I� �=+q�)�I�6���FSѿ]f�7�x�[��܅(J��a�͚!�Ʃ2n���-�b˙{��hO�I�U�>�x����}������_ϡ]�7�Gu�������R��(��!l6�c'ѻ��h~���l��U���^9!����3زq	�p��]�'���օ�6U����o2��y��U�������ys�۱Cɸ���7�|�8�M,H����el+77���'��&�=��%���j�G4�#i$�l�$@����ߕ�v���WPx7w��*�b.�]k�kIqJ*ɱ�w��AS�k�\��1C��D�[�����t��>�?f�<&��f���Gp>�b5�[3�I��˴j`��f/O݌���"o���jXk[�הp��<A��Ź�5�U�=pP�>�;9�a�mC2�1� 0q���EL��8��V��#ӂ̻�	jۆ����ϜM�	�����}��3����s�f���"OY?�JR��}�-�k[��Sx�{�,H\BT���� �`y�P���p�,�0V��83����yK%�� ׸�(*�$g�(s�nӆF���}�K�F�C˨H�֘����T{{��3�����V3~f@�뢛@�VdH���K(U3/�ҲR�F�7��m���M�}sxh˾Y�O�	9v
'�B��rjǻ�����oG�A�o,�:ow_M"&���v՘�'l�:o�/ݹ�i�Lr��HA$�Q鼪�������_��N?y_֦�"<yr�X"-��ʌ�4OjAX�G�]�g����z�Ŵ�7,?���z��1b.��[�a��eP�V;�#>-��~i�ϑ��v�@��x_U z9H���@�.8�?�I!�|��T蹒MG0���s�+Z�������O�dr?����k1��t@Ju�7%�9?ܝV;��b[B��8_.s��a$�_-���z"�����Z$g����	++Ba�݃��e5��4�`���F�y�-X�d|Ԝ�#���>&rɔ�'_�U,E��g���(T7hBܼi�P7��Ǡ��0���)9o�����M{�$Xdm�AK���x�}c�Q8>z9���ֱ;'b��a'�*��^ DM.���،��W�]q���=p%�T���k,���EV1�@�<Ԡ�	�N�R���
L��y"�o�3���@t^��H�OF��j>�������uK��o�i��v�M�k��gSР�Kt�EZ@��R���.�6�e5>f���ꦛ�K�Epji���bGm(=�H��L|xRK�h)` ��[%Bo���&�����K�+�U�*p��~���]�GG�6�s�u,JMU�K���pF���p��.Lv���/�J�>�%�|�.�� ��~�=�;���D��@����gT��ZL��"ـh�vRAk�Y�A����q%-�n�����:U�֒�x�8�bW:d��++_t�5���^,�4x���O:�#'�+��e��I��.�O�(��Io�#�:^A��[��G-�vƸ�zS:�����3�N��H���H��m��8V {w�� �qW!oz-�DXD��gD_��9M�`��9h���6���Q)D�����c��(=��D%��3�:��tԡ�x�[���߷c܏2���7��� 4� �A��B�
}o�3`�H��h��~6���v�V{��.� �o���W�Y��A�g���WPH�J����Ww���ʆ!�iT9o�?�yU6W�����b����-S�imq$s�FV? �"L�G�.�}oUS��6p��C�鸳t�x�R?q��`t�����m1P���x&�^7��F�u #=(FV�w��F��{WB{��qx\m9���,>�\a0���8<bg��6�-U�'�r������
׀x���J*O�j��ShB����b KJ-I��4#�@,�7p3Q�@�����
⯑�Z�%C��곜�����Ԕ��-�����/HV�>�h�@�)VJ4��]�?�/k��?[����t��GO� q�bSU��H��*���k
�a�ݳ]-k��uDA��	)s��ʄ�/���&gG]jҡ�(>3��1����������L���^�#��˳귭j���W����n_ז�F��[}��g�U�)Y�o��)��e��M\������� ΁�
�#�(9Υ�e%p���c�^��Ĩ��߻�OHe���T:����x�|��MI�&''Zeބsr���=u��f�噯4���9��2�U&D`�~�"@���i�-�G�� ����Ƶ��z)X�U��0�8��/(����1ɺ*-��I;?��1�ب��F��uA~J�0�=�3�C�#�ɠ������(��2S��fb2YR���jY����7�Gdd����M�Q}���*/��҄��Ӽ��zg��[Nng�/s�~2� g�袓nctο> ��"A}j�U�Okg�
�x9��Ċ�5��S"#V��xVԝ	Q� �2�і�|a�j��B�V*�Y-�+S�4��{ �!TJ�����^�2OJЭ��D]�q�V9ZI�ڱ	L��M�N�{���j�
�&����t?bA>0��zMϬ�*I>m�a־#����+�g�:N��2=#���#v���a�
й�M
�E>��L�����jA�r*�(�U��h����Ob����G͜�?h��j"z{0�y6��`'��ֈȠ�Uh�e��h���_۫�%�d�t�/�x��Ŷi��{�oz��sw�=�O�ק=�*����%�{5��k쫖�gخ2�Ke��1��t�pp�o<Zr����T�+�������x�+�J3+���쮣�KqX���cU�-c=%]�v���j���r��d�˻	0����q��K�N�ۡ�|w4v�=�B~Ba����y�8������X>8�~����̝@P]+��p�%�(����<[��j�����^O�<تG�!��K��x�̩���/S3��]�&j����j��c�� �D�э�.2Ne�l����א�ٷ(�PkB�Oh,�&�,�ܘv�D|�(�=>���_��h{��:~ ��.�b��k�|�Y3�u�4�'Jqf�X�3��Ծ�[[�'�E�9��Q����P\H�YȌ��~��T0�#�2�54�K`��1� � hd���.�r ʙ�`^p�D_��ʳ�.�z��Vå��ݏ��o����/+b�H��p?��6}���7K�:t�;W9\�ϒdR���a���)Ȭ��,�*�,n��g�<���U�V�gw��Sp����/�-h�5�T���~-8)���^��>�Q�ĶEhN�;ӛhxF@V��}���=0�U�=��
�6s]t��?���[�OB�Ȝ�ȟcd�稚�Bw�ӆ��,�3�����_PK��z3zx��|���f�t,Q�B*d!�E��3�.�M�9�����B/���bEc����(_ܗ1l�#�j�"G[�Rz�V):t�36P'/��H�t���~3�ꈃ�	����i�c�_�������/�yM�u�
S��~U`2e��ʆ+���7���1w��V��ʱLF�}�S��)��)C��̢������� 9qU����by�@�7�t�4�D�Ou|��f	v�-׭�e�+����V���襄=��l���KJ$��*#������gqCb���"�/!�S��U�
��;���m�3 ,��K��V!T�_�o�5��T�ˤI(Ewi�-_�Fk������v��[=96y�}J�zN��(���T��M��{�(�[s�/s�Jp�3^{�F 0֬�vN>H�qB�]z1�@H�#�)Y�ܿ�E�|Gw4��r�b$8�g�#�F'�r�Z/Kd2;�HF�ጤ��k�.h�N����_����{k?�d_Sg0.� 0Zg�q��ԥ������14�m��5�$~�ˊ��8�1��b��hY�C�R, ��G���/�"^:����"n]Z��1���y��BD���A�����|1���;,�'�X�-5=zLUi�z��p�������e�0K��5R���46u�<���K��@~{�?+�
v���ӯ�fF@^v�SgWH��-y��V	!���$�q�8�I'KM�Be��T��b�|�RS������2�P���S����E�i8 ��$�BEzթ��AY��x������r\��}��靖�)� w��A�X�6`��S�%�$�4i�f�����b�w�������7t�~���E�Ǘz���� \��NW��U��6�qR}�H���+���U��EP��F��H�/9�����\*1sR��[��%ȝy��_�7$�p$K��Al�YO4L�&;
}�(�U ��+l��Ňl	��\���I�
G�EޫM8�=P@�K��|\�R�\>�z�dT��G	�]ҩ��+�Ҵ�X�J�ߑl�X;��܎��
)`�/�DLx���!�_/5k/�Ġ�H	Z�8���W��	S{������ C�<O�ծ���{�k
S����!2�EVnH�����1��M<�/8}�����Zfa��J@0ͺ%qSD o���=T�#{.��l�M�JVT���������wr�b;\�8��ʛ�/#��"�M ��k�X��p@���!�C5����ֆ"X�L�I�`��]�=����>��1\x1>��rh��!�]�9*BO��^m��t�aߚ��uP[��2��6��l'wJVd(u���y�Z���7���}�}Uo�����1KC���2�Q��8@ ! C�h�Ȝ�ԯ�I�t� gw��lfL�������6���x�иr��-�O{�Rߚ���)�k���\b ��S����U�ϐ4�E���l�$�v�Ĉ�݄6���ǔ�ߍ[H���F������r��6����kDCvږ�`��Q�Y�7��;�4���[�X�^8<�n�
�b�C�g�7$���:W��5�93��D�Eql9Î��Bm�m���ʶq�Tn��.黾˩A�����IԮ}�j�#(�r�C?|�����u#�B�{�PmHL�$�tGx�c�� i,�>/Gd���:�`a�#=xG��QBD z˺5�g�)�&�;^ v��ּ�a�ԾJ���"
���K���G(�r���vR���>녝PMQ���zL׽ɴ>�g��uLh�S���G�V�}f��V�ͅ0�I6u!����yi�BV���N�rԥ�ن����_��&�"�4m�p;�j@�M���gߺB�Ģ?���k���#
��7�M�i��l��a���K�r]9� ����Iˏ�A
�#e�s�b0�s�����4IN$eeT��Aj(l�mn����<���`����ߛ��6�Y8��B�F��_�M>8 !��eh@Z_�j^��JE{kp*8���h��*9coWo˘�ݵi������&�ݮ|r�-�Nd�K�]��
CΈ�����V��L��צ�ó�4~�i� n�Df$������	<q�j��y.t�H܊�i\ki�<�Oypg̹����Yc�\��p���ݷkG�ؓQ���gcq/����!����?���������m��n[�3�@��9�˵�,K�s���
�]��S�	���K"={fj�hg�(z/]面&t�\LQ���5���=u�5C7X3w0V��%c�B�Fx��Y�by����L�t1/;[���IR��~�U��X4��`2��p�H�^0r?O��O�����c4�`�Pz��^�
I���O�8n�I".���Q�v�>XS��J��{��3�����K�e�CX=-�)�=&�Zf+��V3���2 ��X�
v�K��쉽��:��A��cnY'D�o!����\LYRt�G��5�oH�-:���]�kPǖ �{���%~�z�B��[%Cl]=j?ֲ�_d܌�����L�+����$��t��yw��o ��$��(ėcN����a@�]֏2�����'6��K������K:��oH�pV
ޚ��eD�JD.8h��Y�^����e:�p���J�z��Rf!���w��\�r�/9p���C�DH;C��n�UnA�~�cL@�gz��!-	���<�iC�w�i�.�z�E�Ng ���Z�Qi�ߣ@��"ICU�8��ɒ�ķ��MIF"�V"�>�i�xp���O��|#HBЛ8vy�W�4'�bn�
�����/��)�<���o'h�M��D� �o��2� O�h9�0%yԠ�i=|�'ᰇS[�ѷ�Z2���Mi��'_a�D�9Gәk�a���R� ]el6��5��z�Ғ9��d�sR�h�Q�V
��ST���� �+5����5떳9%�g�D�xݒ� E��@���hH��:�X
���j<�p���@�Er�p���j�	|��4�s���VH����f]R�{�V��<���VM��F�^yĥ$^a��Q����J
%w I!�e|�������5k~f�_�k��>���PV=׮��x�B�0��TS�צv��p��M��X�'��r�Zi}��(�6�?N8��)���a�dMD�r-�X�UE�^l�=F'�l�7�}�����u�1$Tã���=/�u8��Cg�6ؐ����r@�ڬ���ي�Ύ6�S�PY|�L����gs�]֎�a?vJt��'rI���K�����y��pb�s0����R��<26�o�A���tt�B��h$n���X�5��;tݭ����?
�i�w9�ՎT�q����2�z�#��l�c�V�	�u]G6h�W�ʆ<��1�IV�ɟ�G	R�E��\ �5ug�=�W�,�SY�,X�Xܱ!u�`�[��
�<1�p��A�cIlN��>W�VC�F� �������m_���a*<2���qψAőԚ͠�����=V�О�T���!.5��
)��E�n����CLl����'�$!�|�ɗ�8y�^�,�Ӵ�e �a���x�;�f�C���*d��A�d�Tm��u?�I��}FuDs�	��]	�;:�j�6���GM�ah"��1�2\^�{%}ܘ���7v��Kc5�K�-r���JB�~�������&�7z��Uۨ�c�C���q[QA M���y��,��|��b|8�Kg{UU�j��MM^�D�
���|}+�h�@<穸g�K�6�9�)��[��A��թ7�]#�Va���ɲY6:`C�aFK��BQ�:_mOG���_����1p���{�^��rI�?(�Ux�̨��U_1ο�'� ��+�E)�f����3�b��@��fL���Ò��� &�ʃ{���	�}m����1J�c�I&�M	�&��P��w�8�S�Se��1%Cm��T�c���U-v�ڊ�=�Bq�u�q�e��]�ک�K��k��������;�����z�wăg&X[7�J�n�gWL��u"���i�6�%#�	�j��If������ A2Bg�:��$x%8���e[j�H�9a���@p|�l|��=�["��p�V��>GV�JQ�� �7�oJ/���~\(���!�bj��B ��z�,��](�BBV�a(n�٪f3t�lU������qQ�3q�S�L�Ԋ�%b��N�Ι�	{�����Fq\][�ՖZD���520^��=������W:��8���� <��7�#f��-j�B�	qA*M	�������}/�p�l�>���P�eS��������S����"*vCe��a�M�>I���Lso���Ũ���/����6��k{�|h�������\7]o;-���K� R'4f5P���Si�ͳ�<(�8 iv�"��:�,G-�~���~I���N�s敦ks�8�@`P�f�"�?4�e�]��{~Si���'�<セ���xBô�@I����Tpck�g_Y7�Q�I����g���� ֌�?��S��"���a��7�@$?sG��DI�^���/�F!'Պ�6�OdK逅K�,��Bm�SW����P����
����Fӝ�\�����(iM�xۜDW��~�^��z^�a9��0�vr�\�Qʬa���S�e�h�ϿJnNf�β�<S��vG��ƽ���7�j�@H�|��ZB� t���im���ı��'u���]��W�F�j-����dk�o?Ip�,��*is�Ӵ�ݻ�"wX�p���XB�?M��Co_@�9	��l�ls���ޮ9�i�-�׵�8i��4�B�6Q�a�|��vW�Sv���:�� ���,�7sAV�0ǳ/&ع<~�ac���ELF��Mkݺ�J�(۽���Dt�L�H>_��4���t����Vlc�4�!<�k e�
x0��D�Q̑��A�5"<�U�O-Ʌ�4R�Y��|��4F�\����궗�J|� }�>��/.s�VFD֓�+�O��3q����C5����!�}nj3��J�uB�াn�!lZ�i���%����n�Q�F ����	�JiT<a������]ѓ��N1Mx��8����*O
�p�*�d9/ʨ��L��`����!�sb�a��ޤZ^�|����fκ4��$�OF�z��"��Ⱦr���L��&�~V�n����NN�8�u����`k2�P�vy4emr�y�ּ�%@��a��"Q�9���g�D��/Fd���� ��Mt��E<��H�3BLE� U�3Y��1�=4/]�M�i��a݁'������p_#颮n�M�'<mz[Mc�Z�݄Gb��)N��YYSZ����VTS�孱�*�M��=��
GV�LXq"�:;L{�c��Zu�S�� ��g�, �ƛ]�b,ƥ@���&��d�d�9�QLd�"Uw��@w]L�����0e8w��q��z�X*>
,�l�:�JY��	�x���R�JO�������29<��	�ї�B�/�˧��K
;B�ЦD�_{�s*x�~�
=~�ȕ�}���#�FK�Ȳ�Z����Q� �b4�9wF��D�R�\���9�d�p����rʝ�����2�{%�4jf�8X�H'Q0�����I�QK�<�k��dHĒ8���cW���]͆ۮ��|�Ʉ$;�Q�@���H�|���\�c����ɫ���_�K����t�4��k~�I�y�Ɓ�fQ9����!=���B���J�Z���v����m�5��-x"m�j��-Wg&5����]���\��Ȳ\ywC��ݥ8op���d���W��%�;�j@�\''"i"�'!��s��ߘ�d�D�d0����渌�0$˒�.�/�%�Z_�6Jz*�9�n�3g��}�}�k��g���WW�/��Ts��>5��~0�<}w�l`��?�ai��mD�^��o��@s��V3pP�"VC2�8��g`�Ш��\�;ٕa�Ө�w+uh��ٙ<@�+*홲t���V�2�L�ԃi�0�?`vh��:~�>l7�OY�i����̎�Η����Sb6�$�5Qp�ڒ0��[�Dʎ�.���E��m'ٍ,f�E���e#ؠ*M_��AN*�[1�P'�D����s�1
�h�I_2����*i�gJ�8t�0�g�Bb��<��Pb}��_���SOT�c���K��j;����N(�Hcä�NW������Z�H��=��ZV2��Z��j����;����a��qrշ8�b�B��R��#�6&�-)e�}��ŕ˶^M��[/���=n�R����	�g3Btޒ&)��F�P�,���Z;;��bG��tG	��������`�I�y��nX��	������@Gi�b\h�Ē쫧j��0=DC4ӻ�qi�b���m#�}~5r���ؕ�����x� 8�u ��
S5=.x����|>�l"h��Ć�1�Z�i��ʔ��� @-��S��_����(H�Ҳ�^�t������.�pmR7�&�X_''�E�:�*����S�^��e�&a4D���iʓ�����F��5��87[l��8��n!��ڔ��T�)�󵈼�ȣUau]�ɝn�Q�*���~𥪈�Ax�^�om�lV`�������P�
��Ǿ:��1�;t�h�63"_'��(�0;�k���TfWd7�
)H?C_�A!^\0门�A�ܣ^,=�dn��w��ql�th�Hg?z5�Lg	�i�����D��e�E�4�5Q���N�{�D��Hkv@�ڔ��9�/���ڠ����� :�lN@�4Kv�yډkJ��ە�
y��}�W"m��:������F4k��p�&Z�6�6�O��1$��̂0R�P�� 5�>�3����v����g[�U�`��M�m8�c��e�!.�3D,�5���kc�����+��d���ZɖS��#�>���Ի�h1�h��[��6��w$��R��VN�X�{��{�יj��h�	�'i���a�	58_O���Nc�t-��	<h��O�7iW� �E~.�[�0�䖟�g �֬p��)��/���=���&`�XʳzQl8�:*�j��jK���+򌙡��i/z��i��`Sv[n��aX!T"���ە��VE�$��]��w8:������p��ψ���'�H�骇XK���!����4�;gWNҳ�oZw������0��7x�ą�hg���0yO�*M� ����qg���:���>�g^JG��� ��������0!7}��u
�M���� M�L���҅b���� ��s���Dgp�W����/�5�6����e���c���ѧ�܍wJ�c���Z��F��>Y�D@(����1�DU4�Q
�f.q|���Z�I��`tآ��	{*���]
#�6*y*%0e1[�h%�����ϠB[��&�C�,{-եx�5u�A�$��&�����q룴w�Q�����8�$2&�&�-�n�ϑ*=��Yŕ�F7���� �-)v��T#Ł�?���a��G�(��&"4�)�F�c�(����$�d2: ��h���.׶ݝ�boO�f�B��[��׳i2("���#Bw�Pqf��!��	� ����T��Xv���{�X������0�+��¼�a(�	��'�4"�tV���Ocˢ"�w�p(E|Jg[~<��''�pYΒ��Bo�J�A���Z&F��C�$�Ge<i��߇Uf�2y�\Lp���BZ=��=��(��Z��E�_�c_B�+!e(��Y��
6���Y��xk<|JC0zI���q��l{��_k#!�Ժ#��n��c��2h��/�������t ic!���֍s|�BH���>�B�����H��0��y��Cu���2�+�G�J=�Ky����R���]�e빹��;�� ��ț%=ɛ��>d4��J�Y���e@��|�ժ��0
��.Zq�VLԑ�2.�g[~O@���szc��n8L�+�L�'~���
%p���E��Ь�)�����K.Y��xVhZ(�fG̆tN*�FS�g�$$U�����L+�r�� }�XD�����RX�������`��M1��tEȲ8w�9b����@�}���R�K	/�Em�z�3��t�K+͹GH^(��骝����T-�@�����Z�Hs�&��B����I�+���P'�d�)�g��d��j�'���-�W	!�G[����gd���2�����
�db������xV�n+���k���{��C���ʳ<�#����?Q ����@�]�G�sؙj��z�����1�J�HJsZ\)ԑ�%��l�G�];��=)"P�g��>��6��x�G��f����<
��x��%J��fE��IO��_sx��"�tP%͞k��:u�eX�޻�_�M�i�Mܱ���VTl����˾���ӧ�}�!Q��C�h�=�d�&�L����ΰ��a,֙��[g�%m������"��F��2k�c�t-�\X��4j��,j�hPd(1Ŵ��E��v�!��$<̉-���(�T�m���7q6�2����Z �e�gB���V��v�ղER �~��5R��fA��L�^�[n�_�ݒ�����_�ZvM�3j�$��\M��0�����:�4tg$,�������`�޹���?N.�VD�2&WM��
y=��ٱ�(6OB��N\�2��m�H�F#ŏ����O��y�K���Ts`�I�n%
��֙��Qy��>��;�� ���C�ǜz�|[X	��w�\�P&,gq�ld��G�ܵ}#--�`�F��N�Ufs#��W��G����N�** >N��)vpq�ʐ��[!c�1�g�0z��\N�����re�#���1���U9�UA���E?A�`E<Rۋ���Rƣ�Ӂ��5�����������b��f"��O�N1�&����m��!Ԁ��qٟ�� y�7������B�Tİ���+�.�j���Mq�$ ��(G���,�֥��Y����f��pH�ظ9��<A��fѣ7X�W�gpJ5���m���!,���`r�׆E�/��V���-S���q���A_�r� ��"�ț�=K
���	|��U�f���K�|���M�G���I&�џ��]����/�
N�tS���?��b��Y�( Eop�1���U�<�	
Ɓ�{�2Xt�򁝭$ʘݓ����C�߃��$U��	}�kV% ��͇V_Bĺ�b�x�]�..�_ss
�r�1�������%�"]�?�p ��̧(�?�+��>��׎������x�[#�/�x":�mI+m��0yuh{
9��e`�I��M�L���F
y|����Hwk���]m�T��-`�����q��&^q��G�����a�_BJ�ǎ�A3��A���S�n �-��V3��0H-P	<U�O:�=�Gh�.M�Э��78�����L/{���S!}avp�}�g���t�Y�.�D��}A�/��GA�p�6&=��h��eQ��*�K{�0{3���ֺ́;���� Sr�n�^����x�&�lǘo�ل�\�O�/I�+?v
�خG��@��L�]����^P �%�����&p�\}5R� .I�B��H=^!����<��"����#���j-���������+�~��=Y���\�@�D�/iy����D���ቁ]��w1��U��H~IBC��� �C��Ju�T�׊V�A0�igG��y�]���,��Ah�tM;�R�6����5�*�����3`��<�R���.0ؤ�e/~U3U��o2݀A��8��3�6�7����9"Lc� �˾�8	!S�W)T`5XQ�κ���J�H�M��s�!p�c��'.�9�}(�;,fFt*$���M��m[%IT03fw_&�*��~ca�W|lC�xP�E���7:�ӓ�Wr�y���U��0�KV������y���N�#Kt&5y���HXd�S��h�"S=�k�R�"���L����L��B9Q���HF�D�^�Ȅe0풰8�_{w����+���T�*b�<z�����qE�C�"q|� q�cwjр���b�m�+��������=0Ъe�P�-�W�*�Y�dx�I��*0;�O�h��p�ͬ
�� �{�f'%uJr�28D�A����PIfj.�[#o�|e+Ir�l`bA�w!�F�~U����Xˆ�@3:�s��%�;e֫{���vZ'R���g��7��������B b�����VL�B��M���w����A�����,�~9NA�kȂ��*�|a �z�u�?��R?�?���n��7�(,���	�'c�������y!�>�5�p
�L0� HRg}�ػ�H���d�an�_��6�������l�g��(�5�-����6B0(m\��B�u*���$�7Q@3�Ȗ����m�1�� ��"���CB�Z��ɈS�+ ^g�60g-D�@�T�����Ɛ8�ʒl�`�BM
��{%���"�Nї`:�;���@��EQZ�ت�֭*��E�nZ��.U�Գ��x�r�
!��yGٝa,�.>��:���K� �%]d/ *_���A�i�S�]��|�c�N�W���e�5Ni1ѯQQy�>��F�=�I�w�W��N����c��yR�s,��]����"��يi��$K%�x��J�|jc�&{X4�}>���I��[3���ۂ��_���Е9̓A��S������.�;Y���}|ձe/O�LӸ$[�o�h&� w~��.�[6��b���5	o����U��I�Fm,�CZ�u�U�hn$��9��z�=?��2�ʕ���k���������Hm�4D��V\��a�+D''����᱖[��`G��خ�x� b>]�.l%v{�WA�A��e����D��h3V��~�rt������{ޚ���W��M���GB:��B���CI�1��M��`�g�.1J�� �M;	<t�i��n�Z�F&��!���+�_�7��.� ���H�/� �Y����b�~iu������z���۽���C�XPw�0`R�+d 	F��\&N`��"yk༌F����G7*㺱�����KWQE<WRo��Zv���w�#w�h�W�]�7z�d����&V��@z�{k�"yp����x.�����Nv��jr)??J�5':+�t�Jt�����b1�"/��9S`?Y��������8�MiI�۟j-fz����Ѥ)��@��	�O���i8�*��V)�g	����6�����9�n�B�:�8�JH�\��Lq�#�$A��֢v7A�涓r����2
1?����T���2	4r�FA���6{�z̏���g���jE�ܮ�|0>�k��~�,8`mFd�H%'����@�6?�6М�y-�r��9�����/u��;��.��@��]'a���&z�x�{֙��l����Bר'�F����7GmA5�2��*�
�z�}��9 {j����S���s��Tu��
 ����KT����	�Q�e(�蹟V-hԠެN��ov�7wVd􃺪d���O��?G35�"��o�1�B��������`g�%�ր�J�q��#�l�p�s+ŏ�����aϯ�	��݂Z7(n�D�$�&Uy��8��ix>�8�,j����ێ�{~V�RC§N׿��l�_쪻f��E(�`���ʯ뾑R��;B2�������;�/F���t�g�ݒ'�O��Ӷ�ĩ䨴��8=���M~N>6�l`�0%���������]�dY��\ֈzv͟63��Z��$ʣc��f
���}�]C� ��|^�(11-K:.VrU�d��u�!�h�i����6�(F�@���u�r0<�x֞/[ �'%Ű���8l�,L5 A!-`	�$�����N��7G������F)`'a�3�'A��)Χ�oЪ���r�Q�=�h��[z	TC�+A�;s�j��>������>�n
�Rr?+iŗ�&9Y��-�����ǀ�D]t "fI͊_/�)�tc*�� B��󮘖Q`�����Er�/���L���P�P�: ĕ�p�3@�6��<�!k{SfM��ow���/�7�0aZ��&���o+�8^s�Mr�Ϫ�_��Ch�2�ʑ����%?���,k0�6 ��{� ���Z9jWeX��������ֳ���O�C�Vc�Wc]@�����ѻ��?9�A�gs�(�f�XjI�s9�y�6�1��튝-��.Ky�����u��.Ag�xb4�Q����f)f�_����_����b��
:��fhH�/gd�p�@L�Ԍ���M�k��P�� �WAa��2���sy����ia��$��X˺���Hy}�>Fy�o����x�n���oĠBcK9Ί��KN�2�q����1�E�UԼ�6���X�e�m�wW�'[2ip-�nt� Ổ;�V�(���G�T �**��=�]���_���wc�wCG����d���{T��8�	v�p��Uݭ'�X�É��+(jX�t�ٝ�7\��#Ruc��%.^����I9k�+5��!�5�IC�[�:R	3��+�K.����ĳ��@h^�� ҽ7�U�<�(ꮢ!�͚?ceņmG�HYmV����#�>t�XvqC������/K_�a�yS*��~k��)'q&*hG@1�c�~�c)�_1����uv�6
��>׵�	'
h��퍭ᐝh��dn��R�Z)	�����C�{f )��/��o��+�0	߳���6z_��1�T`��I8 ��ȜqQ�����O'κ��?C��,��6x���Y�&� ]��l��K�?m���^g\e$L2�ݡ�0%N�+�Pc���y�U��C��'�窅h�0OB��4yS��CR�p�kjk[1�H�o�ʕ���\a`��]rXη�`����!�灀N�C����k�����ؙ��� =P4��7�gf/�vG��S�J��Z8�Y^�p�lI�'�b��+�:�94�hK�N�@�7��Kk3����a����rEBQ*=]��5�����W��W[0��%�1h{Ot9��>���wb����[�h��@'D��A)g�~A��
8��ȋ�XKs�r�n �E��_ʭ�X�m߿�(f�tU�~�Ywj�_9��tb���CV6��%Q~~�<�o��Z1fY�o4���V��\��pN��f�͹�#����Lܕ�\?��A5+2D%~�ݣ���?'�|�1p`N[���e��pI�U���eHP�KC�,؁ܨEv`;��m�ڀjEe
��a}؇?�oIHe�$��~�9"���2O@1jԷЁ��?1��Ć)��+z�[���H�A2�9������rJD��4�%F��9�4���Գ�UzBt&3����B#R���CU�%xRl�in��_�Ru��)�͑|&��Lj�p6�b��7�j܍\����
N���t�z\�\�$r�<���,x���S�B��e;����p�t�����af3�kݦ\e�h�וP�s�Z�Yp��S���h�޽�A�u�0� ���M0d��*X4�і*�EЃLpL�33v�� i�1Yq��Q���(�=�S��Ҁ�[��@�������]��]��T��PqL�t�Փ�xr$�c����G�*�����;|��Q�>ظ�tq��^�1� c�b�.���"��jS�H�XE���6�y �)�v���=��������T�L�B�'�Ve���@3���whS="ފY ������	翶(4�\H�|���?��U������%�L��$���N��<B�)�ϩ���8����5�Q��a�C^^�|2�(Gg�D�I��v�3c�-��$��@Ms���àb��M�X��!�~��F
lo<�igB�%�&������y��,	���^eM�Pe~=vi�}�ed�%�1_�X��k)�R�a\�`�YO$?u�af�oZQ��NW����Z��5���N��!w�aH��4�SP]�*�khA��0E�|#�ٹ�kv����ᩔЖ	R ������MG��8��S�7�p8:�e�$F�l��F�l��F���ڌ�����^h�C�_$�`��`"ۋ䅪'��fv)z &��b�2�N.,K��&�:Q[�pp�<�v��=&����R;	&�4�*o��E�i,���Q��HٙwC7�Y㙩� $a�Skgo��t�Ij��R�.;�F�3�V��4��~���C����h��F;��祬�b���P�<ͣ|��_\�c@A��@�Mx�0ٕcɻe&<�^����W���1$��ֱ����s*�y
�kr�C(Q ��CZ��@дu���%E���+�z=[.p�t�L�C�+�r��I�k�P�J�tgfv�	3�yR��x������0���Uiەl�H���9۞�w^=u�Hf�Y~�m�̲�$��O-������x���`���^��g���gŃ�o(C�u6�a��[�C��r�;¹�������D�l�������<�X�%4�Nex.��V�4��y�����<{� ЍBc�A� *7�QfB���0O�Ͱ]�1��:�2�
�z��g��iÝі����+ j������Ϋ�!�$�4{ʹBW���c�b/�c���c���#CQ cm�����L#�l�S=JPϲC��.�>�/z� *'ǆ�g�8ԹS�$E�H}��.9���XY�zQ5���x�X���k1�sr[e�=g�L^)��k�`���!	h�_ʐ
C`a{��Z�?*�b~t1\�x�I��]��4��T��H�u�,oR��M���)lLJڵ]��JP҅g�J�P �6�X���� ��&�|�hx�Y��lmo��fp�:e��%�o�=B��:i �T�>j�q���ϝ�}jo��Z�#��>r������?E��U�v��.� ��N@;��m����X�o*��'�Ӭy(g�z����FB�c5�N�s~��JU-MJ���O��Y�a�ޭȌ�d�"�V�|�����1Rp��kb�G����<d"'�cvK@5L<���[w���x�1���D����K	��K(l��<W��P�R",�뎪R%9�\����7W�*�]8/�F��3���F���6gH�Ru���I@���!���<�A�:���ix^� ҈��w`��s�5h�Ad�Y�ѳR�/�<&��N`[`_^��{���ٺ��實C�Iue{�/A[�J�K��M��P<L��I7u LDNz]$�
Ow�=�� �p3v^�;�ЂzM�� ��]��N��(�����Efja����{�1J-t�ѻ�k��M��T~�6��1�p�r@�|�h��Ce#��{^�1��9��'b6?Uۤ�#<6�D�Z�O�iv3���`ڂ�����-��6��!��XW�qJ�li�)�&pα+\Ǎ��v��t|'9�/� �j��oԳ�k�(�f�sc�˼;Gn�w5t+{{�я%?�N����i�T��x]N�D|�?<%�G؍ ��8�'�*d�k�J�SXK��Mm$��yn�����@���?glk�g��EX��H��߀��G�:�F8�7_r��S�l�4��yH�j�� �p��!ר��W�MQL�N����&��-w�;wZ�/I��\�M̂	:m��FQ�3��nmn�؁�wk�q���7�m�~H)�v�?����إ������4�o�ٿ�c��V�V���܅f���!v�m�,)�4&�������Y*�CEz�'rjxt���Zޙ��H�pC9PR��T��\�ؑ��&��@#���TO�<d�������lpUR���|d���{#�Eh��Q�-h���Ƞ`����M1�R%��k�9�#����6��=i��4�z�Yk� c1â_�=y��|�?�O�����Om��1����vZ�5D�� y���^�% I_�%��k���B]��;]E,L١���]o��\	D�1HE��P\�����w��3����-�� ^F��!�[�m�ό��|V����aF;Zo!� ��i����F`��Ik<z��w4�!QD��s�>�ة�(�B�Fb�S�^�r�WH��a�lhDC�tL	ؾ\����Qv���P^3�A9+���(�țZ-yiN���q(*�{(�iC[�wP�nd��i�"A��@����Uw��H�:Q)]��]���~G��녦�af�B�8�q�����QpQ(�
���L�ԯ7q�L�L\~��1dA� �W ��|<�y���5� ��j��݁�[@�)gi/�J����/3������S��aBG��7���R�@>�d��Z������� M����S_Z��������44r;[�l]B,1��vJpCB-��[G]2�7:�Ju�:O����;t.c�7�~ň~z��R�e��3<�����/�=xRyxHB�"��((�X���w�s��;��!H�q�'�����s����$�9��c� ��H����
Y|ˊ���l��SI�s�����4�~#ǧ�'`��U����VYc�_�U9Y��%ӎ��>e�g����NL�RN�����@�;v��)'<�G%��F�
܍?9�Y^5t8:�l뺏��m��P8�<�	�߷������/S9��R9�L-(�9���S#L�C! �
�.�Vm*��S/�rB����!�1�o[��We?_xg? ��P6�a�_ti{Ȃ?�jL�a��������oQ����������G�&r%S�o}����0�ô.����_�~۝����N�m���s�����*��7������-�	h��,<D�!d߳��i:
j�h��N[��)�Kw�YV�����$0賸��.E�c����X�r�VY��B�.�*ֶ��j��:.��wj�]�)S�7��}��5J]e�$� E�s)���Fj;|F�� |����$��%W8�o��u�]O�>�U6ǊU;	�%3&�cL���',�S��V�Z�Y�CBLÍ��k��1,,eJ�y��J�@��1Z#]�~��٘���^�CH�pBj*��k|��3�V�'EE��R��f��|c���*�X0|�Шӷ��)�O��[�b��#�>�x||aQ���l����m/?�jXy�R
��ϊ�~�aH9�aЂ��ƀ� ��
M�^w��a��}�-HlZL+Z-,]e>��w�nhQ�a��C5b�:����r�Q'��c���º%��9ߵ4(�C�����6v 9~���Lt���j��Եu�fb@�	y�*<������\hW2�X�P�.9�%������.F���sq��A�@%T�Ħ�ҹ}���?u$�2�
'��$2>���(�������"8�C�i���*	�g�������f�S��� ��I��N��c��͚�b{8�� �����`�Qp�J��>R�r*�������kUZ:�
Q���}��iK��$`D�(�֝�q[��tS����(O�HǅO8��6�>z�r�}ŵn�(F\��n[�`���8*�W_A(ؓZ���յq��V�w�׾�׍��}����V���N1w9����9�'>�G�E����ߖn,�){���9��u$�J+��c�b�IqH��:;�l�s�(ku���g�MNN)iuW��'띗{8
�kU���*W��L�>�zϰ�%�,�z9�(��q�����Z���k,��|e7!+����eU���K��}�guh�I5r���a�!xs�X3:�"_��ph� y��'����̑��I��b��U���BO��=FPX���0�C�ْ�iG��>��xp]��G����L�`���ѴQ��O�h?�	��̴-��\�f��.\k�`*��h�Q�R≋����m6���"1��ڽ�LU����&�d����7�~�wl�uCd�b�W��D2�Y%��T��J�=]�%�*{L��!q�j�DT�K �Йp���Y�
�YD�Go��Y�u�3E�o4Rw2R��g�wlӖ\�����uk�lp�j�k�p� ~�wR.�Y�h��Jԓ `����S��'^����O��{�d���?�֊��ׅ�A�ɖk���Y��۽^ۤ��	�_�v/��'��^�ߒ}at���S����`�f�n�瓬�n���	A�)X9�HA��`Nu����빗���_�V6�5�'�"&�R�iK8�M��LV��!}��A!��`�JKr�޵n�I�
kPެ�QA�D�υ ��l����w���of� %��~$��t|�cy���d����%��	����Ȣ�c�e���� *��!Y�B/F�=S-��=�������ƪSo�8��G��!�-_�=���"/����7�_�u3�'��5`�5�P�]7��8�$���1���AE��I��(���!>���f�r;�J_����a�i�57�yl�J%(]����-�����$[�XN�3mZ��mc}�r�ۚ$¸W�l�GI@��W5U����{	��C#�np�i;}>xm�nl�.����*Dx�u��'����Lj-X���@S#���$�H#�����p/ b�da�iO0��Eh����-��N�Tz��t�~li�� ��L�("?��b���sJ���5ͳ�-c��Xxo�n�tm��$�U�����Fyy�"�t>�X���{�|PR�̰�2J�<7h�������/�!J�
�j{�5�F0�oEmUj�����v��gE"��-ZD~��$z�q�m��h��+���˭S2�jm�%d��"��lX�W*��c
E���<����SH�������菗G���Z��$`�EflFe3���4&��;硨�V����f8T#|�"MG� �>������	T�7P�v���~�p�k-W��o�� !g�@���C��>���1%��·��<����_a��ϊ�\�
����jgU�p��¿5;�/�� fOժ�QŻL�8e�K]�;�|$f��~�ժ,M�]���t�gls���9o�R����0���Z�b�&�9S�z������]��ɖ�P�յ���:{�MQͯ��E��k�m$�kx@!�s�<����F'�.����j���2�@r�%�{?[��ChK&Ja=Q_?�a��b�VwyF٫�M}�\I�:�5��n�����id���{$`�'b��#�Ʒ9f��HR�"7�m���?� ǽ����$ |^e����R�l��M��o��v��US�����	n0�79e{Ql[��y�X�>��E�����ǿ��&S���G3i��W?��$pŀd���~nY6,�/I�0[�퇅���M�����&����EF��Ji:���ڋ�e謾J��o�a�b#���[��`�'s-	ެ7k�!G&H�6w.������uE�,h6�<ȶ
�JV�ӡ ��*i|] \~*���OO�����j���}��6ǧ�$�t~� ����������DY-�c9jd�m�Z"�d0�`��[����e�50��6�1Q]LedD�Z~��,�ƓV����=���8��H�ZT9g%��p��؇m���y����L������Y^�-!�)���[?:4O.��Fo#�W����b A�c�U[y�"p]:���P�H-���j��� �������ĸRY$S
�c�KA���A��௲O����ݷr)Ӧ�c�$}@�([M�L�m���H�̌iA��A����?�u�9���n�{�,�%+P�Y����) -8�=���}:\X
�� 7��/��2i�EPC��3,���M�cJЉ`{`�#�*��Y���j�8�#�Qj�!]|n;�K�c�E��3M��-���~�A�.��|�"�B�=!n��(-�K)�:�D�U	����y�>��_q�Ĩ�(��CA���%���_s��EO�'��#%�!�4;#7 ���BSɶ���	M=���E����٥r���ο)[5A�8H�b���H��:�7�p?�\4R�R�syc8�S�ϪYv,���[R�cB�amLS�z�k�����sVA܇8��{��sM��
S�L�P�Z��K7_���/��5�8N�P�	��W�8^Ff����x��0f�e�ܲZ}ſ ��.w�*u�[Z�N��W�}��7Q:��u\�FC�T����b9'MDgi�T��A$g�0� ��P�/7�x
���(B� 7dw�T=(	e���<h����H&w����&��sƷ��rc��MW&����橘��̗+�6�`��	��g� !��q�����T��~QFqԯ�j�b��L^����ڸ������'�xV�L8��49%�FTs�y�k-.j�1W�I�4����YHx}��)e��&B����:G�I�v�>� DE����� @k�w	�'%�T���D/�tl3l���D*A���ְ>7F�C"@�J)!��˱ V)����^��0[+�z�.�R��l����S7%�U�"�G������3�ضт�n��"���X��$�R�b:���JdG��s�4G����^`֪̌3��O��s���>�7#\����.���!�+(�e5H�b�zH"�+��QuҜp.�'wC�54#�e8���WWD�WsAi���P�^pѯX��]�A��!��#�f�o8f�7��6�uY���2�n�������s��	g1(����xH;�s��4���"SG��6�,�i�O����䎖DpY*2�u���5�0�����FZ1��3ߵ:�y�����?����/$�O��{�[������ã��+=X�HP-�#X�8O�nS_;�Յdd�Z��L�B��-/��Z�M�W# A��O���&��gJ�}�`'����"��LDj>NP�-ɑT����ON�FL��^ާZg���I\Z�`�l�gx.���߿m��n�_h��3]�<[A+�wO�ȕO���*��:�7LkR�
c�_m!�ƈ�SC��5�N�X`7�M�������>��31��w��3<#�����l�m߇k�1%o����˯Y|j��y���(3%3a��?�7��gݙ�!0��"��^"�Djv/T�*x&ݔa����'%��էM�j�����oN������M�a��s@AA01m��@�PN09�4W"[�f������"��.����|���ρ� (�'L������v@/T�2���g%���y$����ց�Z�����s�I��|?;Y���,�\�~4hZ��@�x��W2?���HC'b���%Y#�^����R�]�xwռR/U�dm����sW�7��}N�����ǎ'�����,�4�M��������qc���,uC7�Cu")��o*��MIf�����0����,^(�ᘴg��=	��H|�
� *�Kꚩ��0n��W�Fػ��} +:�}\a.�j�d�ǽ^�k �$aΙ�胩��L��s���3���@G�e�O�aWFm��7��5�F$�Mjs�+m=Ȇ����J�RQi�j�-)h%��ę�0\H^3ST�rPk\�E��&N������G������b��8n	g��k���\ �Æ�����Δ)����PN$Ԣ�M��i��"���'�#�C&���]3DF�^��S�*fY����"A�5����U_��^ַg���ϭE?.7&H����zv~�A�w/���p�Dܵ¡�ٗ���u>ǫX%E�OM?�a�[��������W<�����ǐ�fe����⎶x+���a��Tz"��aF�_�j�*m;�9 �@BZ H��;q��9%�?3Ț0���N�͓�Dm�+�}��Ø),�SVܢ6��%�h<�x��N��p�vP8�6[7�VΚz��7�&��%^�ʏf}�x�h�76B��r�$��i��7�k�1��nC wQm�"LR��J�meT���0nI�4���o����g> L��ֺ�O���mR·ͱ����E���^���G�r=Hh~ٟi��{O���?r�CV��]�(�i�$�!����c�@X��:!y6����N����hg΍!�a&ٕ���c��ބr�xj�9��@,��'��̿��$f�!�J1zBr>�5��b뼣��'�={- .�Ij��N�	>a��5�6$�ki)6GZ�����Q��/��$ƽȕ���w����!��|-`��Y�{����)��ǭ�R������H�>�ฌg��g޺���<6z/?`U�U(qi�g �鯼l��]���M��RJVT�.���g��NsM�i�-�/����	�a����/�j�z:6Y�0>�4�y�����#���h�Q+]��?I�]�T�"�J�v@Mr,��/�v�p�ܯ^1�rƹr�r	}�� ��'"��y0�cN?�R�Uڰ��%���0�"���C0�C�2
CLȦ�i/�r��-��ɱU���mƾ��e�����[-�����X�i���������L`պ.D��.��z�]$/[`�|����H�c���L����U}�U���w�$gl��s}N���Ӣ���w^[7I8��w)��1�����T���5s74]B܃+�&� xf��L��\�)��62�$�����!���}ա��>Y�$���}jy�tAď����RN#ɩ=��ɂ~�ѵ���<x��0(��Y�;=��L@��{|Dc�w�P�(���ix^�����ڒ�p/���s��N!��,6��S$E,��o�:F���l��|
�iE;G��q�a���p���ɀ��+g�i��N��G1-@Ar@\s&��yQ^sq{I�w�>Yd�!�M0�!W��h��fю��Q��xS`?pk�XE���v�h���t���xZ�Ѵ�E��e�Ɨ%���aR�Mӱ�AYD��쀝�"���k�+v9 t�r���9��3^ř t0��!uKG�l'��K)�d��w��慪v-��^�� ߀�yo�9��}�m����f�(%�%�=h"��mwh�&#�}�<;����g�H����k�8��JO�'�0��e)'�7�gp�At(w�7���	��x��sC��.�F$����D��h�,r����B|�Χ�p�9�0ѳ���]ӺHr�uفn��N� ��ۆ[!$�Ƴ�O/�`VF���4�;}�: �9`�qF���ৎ�V��&8�������;�B��"��"C7A�ߐ���\��m�E1�@^{�z��&���<��#:Z9:>�}ς�~T��;Q�l���F�i��`��]�����ر�0ğ��&%|�,Mu�����/����_o�7@z����f�	�]Vc�К�"�� 2�-5'g��/$3����bN�����_t!�d�s���G�����v^hjN%�U�N�8��εT�W�Rs�	�$(6����Mܢ�N��g�����Sh�a6���̜ׯL&��
�"fOS6��*��-��z_������q���s	�f2�.K�P2�cN>�.}���99gB���j�����;C5�JT4��D��K���>$��j�~���Z��~J���:q�sO�|�'�ݩ��Ί��R�ς�W�+����,��Â^T�P"��R1n� �UI��4N�On��D`�a*͈�,�2��&s��Ri�DA�ݲ�7�=�#���M~����.��[��
�FX���e=B�*gS�~��Ԛm+�O�r��$�x�r����e��SoO�𵉶x^��HD�T� ܩixZRIm��ݡ
,�7f�愱��᫊���\Z1�9�.�b��*��
g����֍�C�%3�]�$v<�j2�x��ڒc�۲���i�6�����`� u��#��Җ�2o��oҤ������zQ�"��!�W�d�|���օ���� �b����$#�El#��+U�� �n��%��}T��!#��R�s+���]�r�¢�p~���ƕ� �cf�96���D��wV�eA��<:�FWa�}�O��ߝ��_���p���%U��]pϧ��&j_�q����
�u���z _���.��w����=�4���NMI�VF��z�Q�-` ��j/"�Ӈ~�C�`NO?X/��)�)������Tb'N�X.&��2;�=���.S�0bb��4���Ǉb���)�������7�K�g�Es t�5\ܛK+�KD�s���:��bWڟ��t뇒5<>��t7駷���"�����U�,R��hӘB�F.On�Ǫ	�fSjě���s�����w517��3�����r�ye0#X�g�p0$�J �b���I���Eo�0?�^���7�+O~�ѝFI,�p�0iu�>r+L^!|;ߛ� .�<c7P��Y�f.�!G�� p�?�����Cs�[� Tז=on0�֏�u�< Ҷ�Di�6������J(�0iW��##��Dz����d���6֕E��1]��� �:l�t�?�.4�h���~܂���Tό!!��ł�w3�>�%���1�p1	fMo��ʳn��t���A����[�"��'��1e���GgM�+�~�/��O�q�>"����%t3��|��l�b0C�Qm(�5�@���!xK<"��n3�kv�B«�۟F�^Hǂ��P0��q�SE�� �>fџc��3�1�j+�5�/� �!���`���{���@����q��Z�O��-.� �vs��n �� ��s�"��K!�*1�*��*����(���R��lJFN.��9���'y�q��5��z��D��L�|�����I]�`Z(%�vW\_��\�&lP1����1;f��L-��Ok���S��!��4��88�Wz�sA�9�u������`�'�ywګ9W���?8�c1�V��?ڹ���W���ߔ�K�آ�?��I4�����=m�B�*�R���+��|�W�xH=���Un���N�9��	�B�z���ZN�M�b�����&��>ʷ�E�/;��(�����e�	��7@j\�p��D���UDY��K/�dΩ�܅���Ł�����rh��/�i'\��ʥ��D��A�o1�@^rJ��k����ʹ5��`X]���F\<�� ֠�[��_�}v�7U�13Ҧ%��[8�/:�]Y���e���e��HH�a�K;���#reG�lh�1�	1V����~�s[�gg�D\�7�A�e`Q��8�Z,l�aR�� 6V�l(rF'{?q�n�A����Y�|��A66� �z;�	V�W����m��.��X����A����S��(�=!�o��2�'�K��b!���qߺ�s����M���e��#h�,a��.�p���;eM7�>͌GV%ܺ^5u&P���\����L�"~��p���@�f-	3ۑ�򙣣�՚��XB�U���{g��O�F[|�!�����d�Y�r�aw�E��6����?��2�V�R���OvH�ҚO�P��
��[��D�+:[D@���g"�ě��R�BN�֨��,*�~�̇��}�<hr=3�{i��a5�l�%~Cz3F]���_*�{���q�`L����4�y+_Rk��#���J!҄\N$>#5�v�_TْW��Po6�Ɇ���	LC!eQw[ܡU}ef��v��
�ͬ�|Hq��wޝ�T� ʫ�I5�K�}���dmڢ�O������,��o>-��Q�N��J?JKʕ�J��y���{�0b�l�g�,�b�B�"�F샪�X�����ۯp���IљX�_p����-˄��dtL눬�J���&˕H�]i�z��ܕPm��2��a���G�g�!�E+��!�&.eb��u��/r{��sv��ş�G��!5峃1�e{k�c๜�#;Lq��b��lI��[�����O��(g��-u�0P�+�#�<7q��U�y��^s=�;����N졎�7�n��wF|���SI�43N��?�Y�����[�v6k�B���*�c�4><����V��Ү��xNP�ul� ���E�ƪ����?[u���{�v�gm�0 �)��F�2�f�_1�����	�@ ] �(@	�&�z��кA,![Ke�O��n���P)��5���-	:��3�Ib��e+��P�j"�<������hn �R�
���$U-�k�a���O��vK��g g��+�K~��W������Q�J�Hq�kC\�9%��[`UeO)��(6�����\F��^(�B�Q����O����qٲL:�7�A7�
�j7�BXE�tTh%��;�tql9�zDIbp�Z-� �?��Fj��/=$Ւg'�>����Zq�EΫ�܀�.ubM�G��U=��)�����GU���E��_��W��4��4C���*ʫ������ƺ��-����0[���*rx����d_2���������.��b���C������o�@;Z�6�-�hJ�@���$Pp���-S���K�Ճå�b�N;�R]N�m�h��ߞ���V+��V25�ZU�{�k�i����*�@�`���U���F�rA�������6�Ь+7�AON|��lg���:��B?��/0S��֙H��C�+dj0��ex?����2�PD�s?�c�U��|n���R��j��I	Q�,א2��Pd'���0(���@��Q"�WÁ_&��v�W3`n?$FJ�xx0,�փ��q+�s;��+I�ƿP�MeV�������	��JR�`�hMۄSNxy/9��*r���$���ǶDw�]����w����-�W��dB�	�(d! "����8�M�rH"�m��Ԑ�Qy�m�����r�q/
�L"j�%OVHJ���D���v�C7��4g$'
�4LT��6��"��dE����&��ю}�6�d�S!7�2�@	�c8���ޣ猔r�2�`���C�-��uG��y�#��R���j����Y̭e������B��x�~���F�[���IO=n�Q(j����(��jcy��:���f`dy ��(����(�>�[ذO:�X����i�e��W>
��I4r
˂�VY^4�Ǟ�T4��[�g�̡ ���4��F�-���"����$�ks+e�B� �w�?�G�(&�e����ѽ�������Cx�����ɘ�bVԷf����4私�5t����bm+��{�����[l-�_WXĳ�P�h���t�Y�7�ִ]�S+g���"��B�:d���X��8���τ��� �!��'u�o'!;N*��v��*����K����8��"��=�%a����ߥ^��D��B2-��'P���1L��a��]*QD��w}4�d/�蟐[N������w�m,��2*�4�WZ�]2��۬��=�R0R���S��Թ�n��D �c��y>�>������/��3^w�fLJϙׇY������s����u��+�!���a��p��~���a��j�	��4�娲*��7����g}&�0>�DXh�K���c8i��O"�W���Ƃ��y���b�?�	�S��
��H�\@��Af�P/��G��T5'E������2
�8��1˹��]�-�����n�q`�F=�eկjE��l�-��f>�V�BE�%������-�=��Jg�̂��o��#�9���@n��g���]d��=�k%y]d�3����W�ݚ^�Yb�<�֧��E�����z�Y�OĻ.M��|����D2Ң�]T��Ŵ�ZO����=P ��tn���/�̺v-�}� X��)&(a�aȣ���A��6]�ѓk88�Pɀ���#�+?ft��]�5۠0�ܼvO�nZ�O��-�ջ��)Nv���^��'�V2b5�F�u���v���I
A����f�Lx��G�ԁ\�*��lߗ��=z�����إvȼ���My�M��s��F1�}̨��e+���{���R>��X��iW	� ٝx�:�ն��-���������Л�j�i���Y�X�b��.��K�3?�-&�t?8s\�:�Y��qǛ'�� ��t�o,�	B�+�Z-jK�^�*�Wu��[�E����n�Ln6{0��|\�/&JsI)�l����e��xT��kq�=jUt}�|�#�[��,}�L���\��LԆc΢��JR/�=o��X����M ����J�GR+D�ٞ���>�"SXq�����������t\e޿�ݞM�1z�L�:<zq1y_����iFB��<��q�^�۶�#+�X�L`�1����!���3�<��ζ�&�A��ye�� f� ���B�K�3�n�����ϔ�ɢ�A'N�,��1y ����(O�7tIZd$St6�<� �=D ���P���g�CiT `�&'ɮ��q��wt?w�+��t�!*0TF 6��fnRH4�G��.������E����Pҡ��)!�a)Sny�H��˖�a��-Df�F棩�)�384@Rߑ������E �������N���{wi��"�)�9�J1��w�X�^�7�������m��ק�/rA4���|���/�-�ϸ#��2�ǘ��{��}4R*Eh���|b@�#��<Xgw�[�s� ���R������ސ8�d,5УԊfU�c�K���\M8�$�,c��u�)�~�׳��n5��=�硩#lopA��pQz�8���zf�����>�������?>VX�wMam�+u0{S�(���΄������l6 P^,O:&"�,��gF�)��͆+)��g�}Je�rgy�ۏo��C��,����������z�5�+����6A@N.f@L��K��n��S;��0�Lg���e�(�"��U��#�	�����I��77s:_�N	�������,<j�J\�CG��5�P��=��#�t?F�Z{vxA�!�r���8Qr�Upuv���P@�$%��>!�Z`�����y�6k����յ5P��`b��X����S俜����ҙ�cd�] k��Z���)����5�����=9��;��#��6�H�(/��2'ń$�$F�v�ZY�iх50�t,0ܭY�iq�IY`�p�U��/C����@#t���g���ݦ�H��ƿ`	xk�!'��dpE+я�y��ǒ�QG �v�S���N:�f�' �8�]�{�n��V�����+���$i�c�����H�-�k�� j#`��J|$��!}a���yr�"�G�#����&��9����q�V�{
��?��D8�mV���c4[�P��6M�Ѯ�(�+�4|�Tjh{l_nb���<�;���7��@VZ�σ�~�U�8��6���a؝/(�����2�'�l(��S���#pDt��U�2_��Ƅt��P��)8䣨W�h��5a�I�&c�D7��忪��`����A�0��N��YbU�{���svI��B�b�r��H?�%�d%>�嶶<�����m����oJ�/j�>w�s�����秴�Ř�B���9��W�6�s�/�q_;Կ[��q&O[��F���|�m硩 ���\��K��I�w"�=�5Jy�3F���p�]��8j�`a�q�l����'f�Լ"��/�(C��m��Pˢ��$:O��a���.'}�F+T/1�g<N`�u���_�CK�S�±�t:��LE��F��?�>�Ui���)��"�w��:ΰ�<��選�����R0nߌ����u1S�Kd�"�mz]�ů�b�Z�i���r��l�1��� �G�W�Ss
)kBn�̀�D�{f��l��EK�Fo#���B�`	�1!�"��/L�������.�K���S/G5O�ߡ2H��P��!|���� *	��w���x�O�N��q����N��P��[�J���IXg��S�9?L=d�^�J[!�������dH�P=�g���fe���}{��\��4S�ō�1�^Lc 5{G����
�受��� +��m��}�0��igM��*��;�V��W�Yu琶R�q�h�:�N���C;�����ʜ��v��g��+3���ho�L��Eu�c�
��b��������x.#ܴ����T�x�E�uQ�]�x~��Z�\�"^�?{6fLi�%�|�՗���'	��M�L��oۺn�����~�����#���F���L�p���i�o�9���	��y�	���d�n�$xt�E#��l4
mW�� ��Z�~k �Y&�Q����	9��4�9���ʎ����M�쉥G[�B@F����!�r���]c�� ��̍sDj�_�j��Û)���%[ ���ј�KBM2"Z��5H�\�+��χ}��>uu�F�@1/�ߢ�����j��!�GP;#iu��"A�Qb}Έ��J7��~(ս�HӀ��b9� %㥚��x~�ٶ��Q���ƙëM��t⺚_�~�u�V-h&��\���9w���OZ�A~��UjK��p���%���]HhXL�TV.E�29`��弄���X�.#5�Zhٷ���=������^'��,=K��M|����p�ڵH�b۠tt�fã��5��|/+n��~�+>�E�I�$ْrsVd'��+��H�kL�B���1AH���`�%*_�}]�#@!�`�ۦ��.P�E�7�����tE�B��,��8�ߝ�� ΑOɳ���O��� �s���F"�@J�Hs��XY��^����$��i=Jd�Sj��?Dmy���r:�Q��߽/�zҞ(�t�k]5�<�}oD�H�h�C�p��H�V�T�4�H���_� zM���;g�B �TjH���ر�>�=��]c���X��_"Mq*�Y�*�S��֑:#��*��*BSp�aź�����z��U�&I������`g��3lu�� ��G��!��}���М��T	���-��XT����^���9w�٨PmQ�����@��B�W�){�#�Ϡ��mXiBJ�ji>�}���$˕���FG%e�ϖJ�ԁ��9�1�_�	�J�)��^J���C@�:�;i��х[~y�jm�C��퓏d]l�����,r���L�S�ґwҩ����!Ơ�w_L��'���z����_އfj|R1:p�v�>��YfA�~x=2�t�����y��{w������@�D�>n���t���f/�,�<�
��"�uX��p2���I���q>��̙c���$lX���7�:�����vԬ4-냱���A�A��F�T&�\�8��2�|��g*�$)�P�Ɇ>g5�`:Z��0Xt%k���a�"#=�p�`�1��(q&��UAx
�&����6�e6�؞�����P�K��?�9!�PZ��M���Ra�)��[�/]��Zc|1Q��Mh";�(y+��+'.�)�HUӂ�i��@�鯸��]���9e�ֆ<��dR(��L�6���>�e�F�e��~��y��)Ea�jxo�ք�0F��Qڰ�2������L�\_`�f 6�Z�JW��Ap[>�O)(��W_���R���L���@x�!%���,.�14P5��ɿ Y�4�tI戗�f�j�7ӆ����l8�ߦ`*���1��� t["��={�k��h 08s#��մ�H��VB��K��o�>]�@���|�!�Lp��D�mGL��c�/k��[��<�QZ�d�N��(t�\P�EL[�JM^����:?����
�
-`GRs���1�jz~�"�6��!$j���Eq.�P
�E���P#������g������<�}�oY�A�7��b)��Y&V5ƭlb�5�T�1K_>�_=d�CW�:���k�U��=��}�%F�
�W���I*5�����`���-AGm�l��q0$�䱳}�r_\�}u�XT5S��{���[
�Ϯ ���B��z���n��rF�[F��΅C^����j�l�7ڝ������{�����?"^�Cg����A)6����H�k?H����2�:��Y'�H"K��UZ�<� ��s��[T^��HN���V�0Ȍ �w0"p���=��\6�{��R�r��D��A��L}&�(]2��*G|��OA��G0,e�=M��e��d�D�~^|%���d���<����㚐Hw(��/��yiv���9?�FB݌a�Y���Ԉ��p��@�-8�ԧG���T)�i�3����y ���	[��I.���0#ۼܒ��ܖ���7��7<�F�@�����$�v]-�hF�u"G;
�8!~��)@�>u�ѻ�_VK�	�	v"��1��WE<�j2���FȇHN����c��4�1%PH�'�N%7��xв�ZB���+v��,�s�ml�l�	�x����յ���Ua�5%�5$-��-������
B$����DdH�u{�<��yp�;w/�dC��p�n���f��N��|��R��F�Wmv�U�[��;��u���%�q�]�sU ZBN8�� N��
^�\,�`��ű��R��W��uJ���(p{����t�#@�9�	V�7e0��gA��pO��g�w����N�Q�m�W� N��`�Iu�Ñ* >�pÉ�	ƣ
���|e L�`��1����髸�%ͺԀyILa�����V��[�5���PX U!Y2����,I�1a�; ��}χ X�g�O�ጏ
%��f��G�8��嬹��p�9��� -��c�bf��w��1wQ��{F_����s,�t_65M�ޔv��4�Ak!@�ռ���+�.�x���g��P���S���!��e��}���4]�.O5��P���!/[�<S�Q���$d)�\A��0z� �5H�f��6h ��¿Ԉ�ɓ�x�X�1TJ�&�16%<T=�?�cG"#ͫ��VD�zhAkl#H"�����}tI��ң&����磗�>v�6إ����hl�"6�Y�Hzm����L��'#�0��>��FM��/$4�;!t�;,Os
�f��n�XS�����x;�Y+{��o?��Y3z�v��e���F�!���K����C�z��������t>ZD#�q�!4��?�iw��9����^�f��[��txD98	ZLL'��
'	���ɥ�FWJU��m�^�C<(�F����1�Ѝ�tf�u��t����� �;{/��
NЂ��Y�
��R�C���`��� p��@��65'858�w��v/֨�V�g[�+��mO ���x�~�ԛ; ��=a9�`��(l!L�;_���@ �|ɐT�Q;WC�7�	���©^�V@���e�N����p��h�b�cT$�:�)�3/ηU�z���d�BE�&_ �uU$���C�7�4���|�2^�8ŧ��'�Uɤj�!�4u��R_�2�X��چxW�'s	Ͱ(`V?�O3đ~�Q��sn����#)�B!�5�x��7F�}w�M������J��ٯ�o�ϻ����`G�=�]�˟��; ��-U-)G�o��kך0p��w	tc�ٔ4=�]�G��Ib@��8U�:F7f*���s�o���Fz��CQO:O�"����n��S����ӏb��wdn�{{*4���M�Ó���F���W�1�ЏI��~�m�P��p\dj����.��z	���;](;����2d>���� �ϣĒ�����e�[�˙:d�g4��J��&☊�÷���nh����'���� n
J���F�S�"��� O���D����Y�%����w��s�9��
ptԗ��kbO\��Gp��"Κ����3]���rS�m����� ��x�<�:{d�n"�Q��Xw����|��84"�$��'GeB:v��\�����Ρ|FN������%'�2�7#|]+Ք���d+��#s�V�4uI��>a��%*O��"M,n��H���r��6}�C��Ɔ6�h �� \�}q=��&Վ#�yW$T�m��}s+<=���0Q��Pd/
��
5ZH��������8AևtXB�åIY���Lϳ�E�~]�XK��K�����F[�<xD�:�����ySDS�/�)����C*�9�ܦs��X�j�	9}�B�g=���
�TѬ������ֆ��N�^	�z9ͫ�*�_�}�#��9v��w�\�,;��4��5��a5��p��j8i�q7{���Z9NP�ǥ�&"�a�3�EӼ�����9�z��ϓ����J���8�_����>e��?�L�}�d�}B����x>&�Rֽ��RJ=���A�T�7yZ$���Z<���
��q�ʫ�L �7�;�1��}CCl��A�h�4D[�[�F���C�m�~q��Of:��ȓҿ�~��V��������/7�Ts��g���e����"�4$шO��������-�ɫ���ț#d�	[/�����)-%�+�N�k��CjE&�v�/�F��m[���M�ÍhTZ
����lzjV��m7P�m���N�J���-w�E���.�X�
:�EUg���t��w S1�œ��ҧh��m�U���m˥DA��I�I���Ub�`i�JS�l�7e�vTt'ŉ�����zG�C��F�(D�G��[E�3%_��<�U@����9�}C�	Mԕ:e�k$�sǂ<n�|̤帄��~B��x3�H���N�",��(1���j��f�9����(\s�6=��S`�2�>�B���������
�1��`����^U]WEJn��/��*���l;�i�KO��i����`"����Z��)����{���>�:2��J��xp�#����c��&1&eּ��jKd �6�2m�����:�����}Q=A<�O6�9����&�r`��;���>xHY��L�ԍ�#C^��^i�^]�r\�ݶZH�F�c'�<6=���/�z�)~���#Jp����`�r�(@�A��-�&T��L�r��76J��w��_𫸅�ƚ������%tJCZ��9���6Z��N �5=�#�&�Vdc��4���K(A2��Τ�5�c��e��Isݸ`���p��� L�f��f#)r�\G:]d�Ɣ�Aml��G]Μ5�!�{�PŰj�R*�~
ג�x�<�y�۵�c�D�+ʌ�~����������6�7=y�"@�)���)���o]N��KR��Ɇ�Ϗd�W̳s
b�Y��EJ�SF��F/ ��p?f��U��S�揖�E+��Z��νeAܟ{)��-�lkh�wy�E;NO�j��t��	�A؝qG�6�S9~�/�!��T���"������1��xD��AH�rѴ�n�w�p�6�Kf�ؼ��o�]2Òq�"�'�N� ʚ�
ё���w��T��fցo�
7��T���S�M�H��3�l8J�B`-�!�$�Z�;
[��f����2-,��sR��ӭm�J�[����3��8��N�=��9+�޽ݣ��Z�0�*��o��[�7� 6=fm}kY�+�fJ��}�Yu�)GVJ����v��o�-I��T���y5�JXR�Ap�Q�(v��~��η����9���
���M�X0p�4���h�e	�49�c"�쬆4y�����-��(�e�&_�"���Ӷ���?3)�E�2W��e
��{9���1`~?;�v?���� �J�=��=�
4�:$3��91:dj��>,z�˜��&m)�;��J�sO�C�_��B�V��ZuH^2�^0��AA���L�rm%1�T)���r��Tʾ�t����_g�;��"� �Uo��~����*��ę�Vv���̝pK"[w�y�/_3���8�MJ|��$�`�x�D����Ӌ�Sl�<���[��@+Lh�-�s�n�U�"T�&��]��KT!%vT��}�@?�9XI��W��� =���`�IDG����<xKM��W�,�O>L�? kV>!Jz�R�#<1�B���l������Ӳ実b���N<�-�BB��H��J'.�I�a�ͽ��;��u��Ny|-�W\��, H� ���o=Ɍ7���ؾH��0�r5Cm(=�@bFS��d
T`�M�
�d�ʦ" 5 ��ۗm[���J͈~��m/�n2���f2-���U`)�����S�M��	�P;����Dg�F��������	<�M/,����N��zi/BJa��DU�ӡ5��y>���'�a�n��]��\�ڥt@x��o���>�S�e㽻$�n�yn��|�fEj�pa���(}Ew��gA1Ujy�bb\ⳋ��[�.-��A���h~�"WK'[y����8U �-�|�0Hl�Z�|���{j�h+�Ő�y��ko9* c����x���O-o]�\Pi��+����g��0I>�!�'��~�����W+��Ul ���}VP�7���Dh�x�@�xt���VE���0.ӈ�V	_�%��p	U�,2�T����6�h�T�KcH��F�(k���1����x��.9]�!�:��L����;���ّ�Z��
=�o�m5h��/���������DW����(7;#�e�Ѥ� ҂�H�_r �]��˂&`��*J����ξ�6I׮U�|������+Ė8��pi������m�\cA�7.���CK��~�~λ�=��x,.4�@��X_
͛�'�bJƯ''!�&˥4}P�XƳ@X6�F~a��3�R��8f+//`�(xTԴ�׭6FAĭ��}�X�^��A5�e�v��_TX�"}E��-�σ��b)}z�YWx}���F��)�ff�w�<Q .�T>��&��W�롩�Q���
܊_|�C��&��ҩ�@���6�;@�+A@�!���ͣ���G�i+��m���j9�"����r�h��Շ	iW}᭗�_#�J��[k�@��9������<!Ĵ�6��*$�����dǏ��{YQk��C��-���_9S0�'��y��AN���Y*�J�CN[��Ɛ��)�m���%W��;b���X��1!y,(���8���ִ��Q��&	�L[ �`�;[���Y�{#-z�'�G���W�z�)�a����i�[w����॑�Q�����N�`wK���`׸�(�V��9�'cE�P?�CNC4�^�l��71�h:K�g%܈^��H]�͡��l�P�2ZF����@�g��@2J��5���nZ!��a�s�	�עY�!?�OT�X���P�X[�onO��݋�zz��s��=!���T��Q��#�n� �E���аig��+X�1+4�z\���h�2���y�.��
��,vY!�z�_ ��Y�u��r�ފ��9����\d�V�����u�1pY��YB좙��=3�FN<��W��&=Só�9��8T���P�Q��UfE��oOnd��'�WXB�&@{	��P�0�/�������GC͵�'�p��-A�H ڴ��� T���2�'fh~5u8�S(�ӻW$Y>���T�˕H��b4�,�U��_�&�E�nH���A7���F������W]����WX�K�	��𢒗�I��H�%9�t2Q ���:�_Z2���Բ�Y�������|�J�(��s7�H��2���ِ:�K޶�N��0�r�iz�c(�fb�<C�[�੟���Lm�r�cLV\��߀�ퟩ$\D(˜�,���u�P01ĮT�Mm���	)j@�� �ӭ㹓Ϡgԥ�;*���\��챫����#6g��u7�Bq��h<�����?<v�7'&RVl?�ۙ|�����B�bvqf���92CaU:��
�V{=H��I�h�}�v��B�rw����0�8a�S��=�զ�:����YRd&�M`=+wz�ÝE���E��N%p�0:5���s>��ۣ����%� ;m�(��UI�+1�f�!fj'�Mei����Х�3ڮY���莻��2"�&yl3����߸��M��9�%2��u�ϧ�v�x����>��n-�:rmzx)Un����)*I#	:�/�2�^�}�� ���.���m�����ư ��w!�uU+_�(R�强(����;?�
�*]�H����:0���#^�4h��_�Ƥ��B�_I[��uc��c%��.�}� ]�[z*�1J�9��m�{ Z��u��'kJۆ���zn��矒�L&��k`��.�d@�fA�X�l�*e8������ ��J�Y7�.)��m
,��m#��g��E�VSb�qͺr%�~׽� ��ǩ1P�f�_��bbVk�}ǚL&�)��a�p2��҅5PY(w��r]V��2�H�����Ý�l�Se��8��f��61�z�����H��z�2��a�������V���P�L��v�'=�F3��t�,Q��	K0���P
��c�8�������9'�e��y�K{6��C��[j}W��s�C!�2 M(��Dum����r6
'�oMjP�Oə��%�G��)�7�4���ye����3�����ɮ%x�iP�Ys��5��B�rMȳ�)�f>��B��D���N?���n�k/[oC�P���z�Ҥ�J�e�_��m;Mwr���
��{�%%�?�|�k����_������~.�qR����f��1�����{��^N2^�bw�<}��Ms,������F��T��2��0���W�hi��Y��e��P(�?�Y��� P��)��v���`�R7�ڹ�{0�:��SΩg��Q�5�_�;dx) j�	����FID�EA����8&�?���JZ)��w{�®g�g� ���h-'ɭ�Z�
�S'	ۓ��cCP��ppP�d*`�M�����o3�Ό�ݾ|F��S��q+��!{$��J�Z/QƼ@�����)��3q>N�ŝ��W���읭�g�̈́!����1l����ĵ��7\c�2 �+�p�i���^|յ�|�����4����f	=��3�O2�l$��죍���Gzv���P��|�c�_+�é��"��S��n�|�Z#�;�*I�v�)����沎�+š��չ���8���~Tb����DR�"�yP�_W���ۋY��e$0p*�
��8�X�t[�EԻ���DM�	�Qǋ�i�7Y�xi�\����]W4�9�ɭ �"�-�1m.�i|}{�D�»1�џ���D|e�u�*�$�a"�>h��h$�H�y������B��D��7s�ǲ����y��Vb>��c�����C���:!�@.��>L���b�n�D_��{xqR&��3���0�*Rz�4ƥd�C=��J�ﴇ�7����{W��Sd��F����Z���_��I
$|.���Hj��򰙪9�_�T�$*��$ǟ�P`s���
��f�ja��0����6$�ǫ���d���
�
k�s%Y>�duНJR32mt`-��x^��񐤆�����a�Š��!�Z���	hE�ue�q����(�w�2p����.��?蕥�`*�[P[���Ȑa�of�jb-�jbu����Ucۦ��|�dy�Za*�ڽ� 4�M\���;�0_֥���E��1[T��z�1#����V/�-^��˧k���!������VP��������>zΜ`H9���d��7c6l9JkP!~����R0�l�v���1���Y��3�N����[��q�G�3���yN���ۡw;A�w�O5)w��3WB���L�"�< �3S��N�g�zQ+s}xVaz���e-��J}�i�rp�c�{P�� d����Yx�m5y2�9'BL�t���ÅR���z��=���M�Ή��O�����BP�ش���b�rq9���6d�*v�A ��z��:eǧu=�	6O1��ڻ^5��Lh�~������}�����N]����繮�� �s�b?r|�:]�g��lm��I*h=����P�9!�C��AÀ�s��9 ��y��T�I��2���c��5�}a����8��jS1c�8w*h]Y\Aj���%�t;@l?��4Kǝ1�	nZ����$3?�#D��ooB����c��s��٬E��juURUR������Kġ�6��8�^���3!���^&����DsS5DLo3bf��&}	�8S�������NZd��N��ޤ�=Gd]��˧� �:W�.X�dc�S����iǤ7���Cg�F�����.�Ħ(5�h8s�~ �D읃O����|U%�`l�����3�I���%��!w��'�	��˹����m�h{���J�$5��_����MG��t�����$���Ñn�#$�O��`{mAu��L6 �M�X�H�D��؁.C���Oa�@0r��̈́�<b��PJH#'8����Yy~�\9S��9��	h	�]-���>�H�٨`��%kCI��Z���yb�x�2_�E���G>dO���r�:-�%��B���4� �X�N�_����.���*���
E7���R�'1���F,|A�hcY��Y�s�r�#�&�A=,1a��J)���eycl#H����̛&\{V���f`<��X������w�m��1�c�M�!�L�:����EGTnV�h�Kէ�x1�#=����V��q�g��� ��Q�Dfh=�9�AB# {=�0T�~*�Q�؇��F�%L�M�Ԝ���<���i]6����� ����l��C�;�˷}[����{۝�ZϿ�l�o�Z�+b����.y;�_&rT������ �5^Ğ-*��DV�;J}8NbP�&�������������^�0İ�Ie�;��ռ8�b�S�j�yMɍ��-k�=M�kq���!��'(
�n��d�E��}�	
H"9M��|�< LڱV��M�9)4L��8��l���&8#*��LĝaH>Q�j"��W~�i����}>��?�rjt���D�R�C6�aX����Kϐ��u脽��rD��'��x���,/��)����s�����2̪.�z���p(�t���@k�
�t�a�[����	�C!g[]_"_m���˺ߚJH����|c<^��Z��5�b0Z:5i��}��4?�P����Y�pE���$���D,�X �8��F
"�s2�c��@цN��,���
��	����L������ �!�9���)+ET�K�
�F�R�X��A�B�4;b~��;^1�}x�z���d�5����=��HK�q�=�����I�+�li߶V���}I���\��`�����H6,�EQ�;�poQ��s�ػ���, ��M^d�l־��D�6a�fAfUBY��N�"$Q�-Z�74�I������4��O�C�8��A[YӪ�0N�D�������q��Q9�>�d$8(��o���r��f$��8|B< +/Z?5b��-�{_��d1=L/���Z�7�aDo~�g6��2���1r����Tr5|�̍���]�mt�,Tu�+��A�:2*�mz&E7����?8J�KN�r���[H�{8'n{su|Z�'
>���(d����}��x���5���ـ\_�]�X�`����L݇�F���c��cJMH	g�ö}�;��Ϧ^ i�Ƅﲼ��+hJ[�$>�[��y�
c�L�ht���A�9�W0��IH,o�-��A���M������� ��l M��Ϙ1�k��X�+�:�1u��,�:E�c�Qq���hC�3��}uc��M��.o#j����2��Z=����ȏ/ ���������`i�h�?�jc�<� �r����+���%؟fn��{ʊ�ī��2��7� ��uw��`p.H�^`V��w��9}�N6  ךՇ�^�p�ƀN%��o����,�9��At�D+�Tu��1��)�O��ܔz���A ^GM���E��W���������=���O�5����.Tp4�&<1�9>���4�QKa�-�&-'�n�֋�C����$JU=.j������; ��!���=zꌞ����m8�uN*�Y�m{(ˤ��B���R��"l\Pl-u�$<�(���!D��3�@%�Ǣ�#vz�n6BC�%;���u�8Vt����7�A��{��R˖��
����7�&��E��e��:d)ﭽ�du�Ή���D�����1����d&}��$�ɻ2�d8XjyOf	�s���Չ�T����"�P��5��폋��0�An�����A������iNpo	�o����0I�̴!�������F�;����-Ә��˦����Y�����C�R.D�e�lɊ��052s�Y�K�l!2��G)�ѭ��=Fo�0��,��c!s�q����/�	^Ү���EL)\�Z��,]�<�^�������b3���4��_�������������cHz7��v:��¤�
\/W���:	�̐"���p�t҅�xX��\9��CO����ͨK7�ⓝ�u�����=^��<�d��A`W�R1�e`�̹a |H����2l<LR��O%�� �瑣�	ؚw:/B�s5v7:�����x	��3�K\	"].�(��N�,�&��� �Z�<��g��,f����������2�dc#�Ҵ�e�/�p�"��mT޻Kκ	�G���R�crR�S��˂f�j�Ag던YX�Av�
ǌ5��VP������/�,�)�0���_�w)�T�k�(I`�>���㡉�1��f�]����V����G��ސ���/L�3��I���������h�n`N����i� g�ҹb���M�e�t���dW`�Q��ZOc���tOO}��V�������<G�J�����ۦ���b�h���עP/�Mgs�m���d+�L���R'6e���x�;
;��>.�$m����,��̥��wz�UF���Rx�(�/�\'�c��v�Q���=u$������]��$�'Ȩ���V* ��x�EW�$���c�V���}3J��2B��^?jAu�&U���?���}R�Ң=ʪS������zTaF9��2�eº�7�B��g��)&2��)�9*i �)ķ��`�S�����<-y��5G�<AA���X�Zk��El�h��lWH}D����f`/�0�@�:)h&/]��\6TϜU�t�Ǭ�2&�F�*m�>�yvG"�e�aÊ�8d�@=�����_X���˪�$l�Ʈ?IEM65jwZ!�����ķx)��@'�2S�=J ���P�%ݥ�5�M�Ƕ��.Λ��n�iJ��e��ƹ K���Č0�,��s��t��4���$��6�Qb����)�\��UY:� _9�;8v�����S�߿ex�k�@�m��)�����)�bp��J�AB���u:�����H4���=��)U1�m�x�w�[���0|�Q�	$f�\b��K���;B|�%�M�u67�E�EMz!�ٙ��΋k��ڙ����8c^�3����=��������!,'��d�Y�X;��-���5�o´�Ĺ�
E��%%�{i~��6�?o�7b�������E�����۳f�P�mT�����n��Wpp�vl�0ii8^)>��4���JN�2(�T�z��{F����dh3��"���ܢA)%\2~U��m�7���U�����vAO7P����A۩z�d �4+���L-D��$�p#����K�����߽���p�W7�-���V��� !�OŞu����R0l6����,�a�x��d,��1��[n�a2!���5���}��]R�5򎚱mM�zT����P�r��5S�=�*p��c���|ܒ!�Z��{�Gd��b���h��6��V�Vr��U���
�u��NR]I%h��K���z�PM����o�׍��z�S2�;T��1f����:	����yLIQHLL��g���3����KU���Q6��~ؘ�kV�7n��7�D���6
D�`3$G���S���d{ٱ�qn���e�x~�$��j��X�#�A�q,ʴ��v �ل��yy����[�|�#<P6�?b���n��Z�71�WJ�,��^9X��1��N}xӬ�&��t��槝Ty=!���<v?y�u�9q")���}k�%>q5ra�#G&�$-�����ij=jLCr Hl^LV/���--�ɥ�'(����Fh���K�����5Zڹ��hus���|�DM�8�lA1!��0"���m�F���0_8If�t~הEyaz���u�2cXa3���5�����yL~�c��b_JC�X����ox@���k��,D��'T�āӼW��-KѦ�W��n��F*���8i���~�ZA�;2Y�M\�o@��DK��z��dի.&��x��2�棵lH9�s��q�����k����fLB}�Ԝo��#U��4AĤ�gq�)��8��=���Eĉ+�~���>i���\�#]�2+�;�Y��,w���)l�������v��-0Z>����&�913�V�,�UL4����m-�3q��>����%��dP�ਏ�;OY�,�䒯&��a8݁�)��|%=8R3���/A�:����RߪR�����V�O,}�_Ě��?��G�5�朰�������["�i�P_'�{;G�ݖ'M��+IX�OMG���>V���z7˩�h� r�<�?#�u��"�q���J�99ϧwo�Xўǟ�ec�' 
ۅέ��LS���v���'o"8;D?���z�t�P�����|��5�t�%.BA�t��$ ���f{"�W9�?T��U,g	��X���2@ic_���:mi�5���)��ܧ�<'��V�se��!k��5a��ϨBD���a����6A��|'�I�Silr�`�J7X��҂�ē�a\�cT^�}�fU��,شr�&eμ>w�N��G*��(8���5�/�ub�]7g����as�
���߈Tv¡̀�Ýh0�� ���u��>�W\Oy�P.?�����<�k�\��qn�D��"�kL�i�cc~��Cj�D���k �L$J#��>�� w�/X�O�Hs����-w� Bs��n���@	4q���&kӲ�G�V��r�+ĄE^�g��Y��lZ�2VS���{�I(Il6�D_$]�S���n��&��{�YT���S{U��I�U�#Q�0)sYC��v������]����Ͱ?�sr@����l��������(�it����_���� �s!��*��K9].�T>�= 
:X����r�a_�g2tL1�<hu!������6�)Y�����֟N��!��u�C��Z�st��p�ܸ��<=�t�ި�K���Q��CE�R:μ	��\����{�����u8�1.n��9���2���U�<<X<j�j���*l5-�.���C֛�07�Ǐ�V��w��&��G���Y8P�@��/f�74�n�h��^��l�_n�I��}�d�}_܈���)�Lx"�#KJ�H�?��x���p�֏+d���-*�_ ���c'���ج&M	�73( �H�D��^9�6y%I36�ｪ72�_ێ�ߧ �?�����e�c ���Յ���o'�h?��*��9"�g�!���F�O#�8	}C}�s�4�I���ui�3�"�ɑ_��61%Y6C%��1�<t˨���r\0��}��0�Ӫ�ȣʹO�wf�Y�k�.�-��V%t�`r�6�&��O)��	��7���������0���X�{���,Fד�	@l����K�.��N��G���#��i5���S��T���B�?W�:E�Q=I��q�I����X�Z�� �@`�
�R�y�mz~0��/��J��O�em߆1�?p?�h��%�tZtƻ�H�N���3_z���X�Ң�Ki0nY_6�����̼��C>�P�{�N�ڦ�~8D��`�|�|5���g7H$�ۢ��祋HsE�o�D����3)Bn{����;�p rϬVT"�W���c_t�b����(�j��!+llp-��`��� �ab
�vlW�Փ]��;�&LL\K£�V���`U?pk�.:.`�/sy���g��Id��" �!C	���Y��>���x`���Rfr&t�C����'�Xd�g����>hO�-�Ҥ��LЁ>j��o�Q�o>C�nt_�'wC&�nV�-ߡ]�$�(*�K�Hk{���� �h�p�͐M`K��Vq'��d9h����Y�����X�9���yr���L3���0įY��f��O�Nf>�4�H�\8���,�����ȨX�;І�e*bcmi��e�ԗ$�q��_}���d�0l�6�S�[��Qb��A��,���{�����p!\c��x�k��#�v��'�x�`c��D(q���y��6Y�#w�)s�h@�X5m��aTi�'	ռ��5>N��%�������w&ֲ�<a��1Ԁ�C1s���}���R�]C뛶u��
��ߥ`�օ�  ��.�LJ.�����=7u�h�I���l>*���p�K�F�����Y�
�W��h��sTm�E��3���xxi�w���q:��g�q�Fk8��E�pz�Bl��1�d���sor�P�^9h���Dn?��J�B�	<�?Y7l�^��u�)G�d�w�vvZE�J�gӀ�!N�xX��zƱzx@D�
�� !��H�����\V	��ڜ�#���&<qn���
�$ދ��Ѷc®��r��\�&"[�!A�.��;ޞi�o7�͏bC,����q�L]�C�,�L�"J�&���>9P�InXTC7�4� D�ڲz���L��p��j
�V�|W+5E��V����T( �E��l�y�ڵ� �>�$bڱ��v�\t9����tG���c�q|�Y�L�w/9�����b����,kݓ2Gǣ8�oBx�V�w��z�P�Z��y��QԒx����6���5#Dd�,���pM�Q��E����O�ɧJjׁ���:��J�	p_����S���e$�/���mש���3:��H�;Q4}*��Co���y��nQŕ������Z�PSIB�3@l��x��>�<��֭v� �؆���Q�[�s�}�/�U�[/�G�wj�Lr�*��?����>�-V3D�a�w��ȩ�.;4�vǭ�1=]W=x�Ka_�1����R���T教
�I,909���N��$*�~^��0>��,6�9��3�C�-G��&�E�5���S���`W�Β���QD&���YB*�R�n��~7��u��̼r�A�s��Lc/c�n#���$*��/&V�h#/�wl�g����k
eG�y�ІE�c}��$���%->*;񉇃V��40�İ�[Η�k��Hz��D�%�ͫ(����z/��'�!t����$΍�r��w��Kxۘ9��{\g~�8��'�O�~;ڰ��**5K�FM=��ݝA�X�Xw(Nh�>�"�?8����v]��B>�2����2����>ϐ]t1#kb��lkr��5� �KQ�ُ� �;�WFl��Q�qZ �L�G�m�Z����[@L?z���F��@T㵪�I���~�҈�Z�k��Vk��/��ϲJ~J�r�J��0�f���?�j�m�_C��1��
u����0]>�na@�?4��ϔ���ӅuQ��ѝ�"��'���	�iN\�T�'iw�@C-� ����MT��J��~�Pv ���ύ���Xd�('�9���H���e_'n�x4�֟�pt����K�]��B�\�����b@}}Q�%���\-}A�`�'�!��a��a�j�D/���g
,����(���o�q��C�FK�>�7"�?�-��;�%����O�����E�,uF]������d�g���%�`!v%u:X��L�6��#��W�`�� ��.���tV����х�|G�L�7<��%�N��ڈig�39�����I�]�6A���v�,<I�h�9��|� ²z�D��P�����&H������@ոك��˵Fe���C�o���e�6�Hl��4�
6w����4�� 0��R|��B�eE��w"1����[����BzkK��[Dz!�hN������A����B�	��+�8;��t}���vxw�瓆�9��'������7� G�(�cW��R��Ԫ�z�;�Պd ���N�.cҼqC�S�4�I��C���<+��TԼ�K�:y��
��EzZeАM�7n	..Y]�t�q)�A04b�j�����^�4+�MJc�@���yM9UV}^�� ����p*���u��F�c�*���ZL�a�a0
�����zF�As4����Z���P1�bJlS>�
>�,�F�`����U�k0��4r�Uc+�,
���DҐKM�h@�ퟗ�x��V���YA]�N�HLo����>G��4u�Ξ� u��:pA�@�i	kB�5�Y��E�)����k��l�d(����C����}����V���R�� 6eB�"��'�2v�������]$��|N)�R>�T�/0��R oe�T���R/����X�6?`�\1RX�L��z��t/C���W��V�>2�~Ac����]{����LT��@(�}¬��.���Xɫ�)_��h�eO�H(28�C�ی^z����>�h޿�t��o�a��4�G9Y=D�wUq C��*Ƅ�����z�"�f?�[��ؕu)�<}!���C�G�x+ v��$H�rN�x���U7�KRb���*�a���Mtq{A��b^���M�XC4���c�����D}�CQ�ؓU��	��[�*�(�Y������}G�C���vz��/'���J����w Q�r8)W�'ĺ��-Q�`8�焊�9� �us3��WQ��J�J5�F�Fѝ?���3��K-�D1D\�����.LT�q|Ƀ���R��5�xh�U��i��j���L��8��W����29��G���Ŭhoͦ���9e,�/�5��S��p#�"�����z�e���f�6��;{�U�u%7�?��SݙzN�A�<�ᒀ`iɏ��YdЮ:j��WϾ:Z��g�W�
9�<�yAۑ��킾���k�����~¿��R�4H��cۻxF�����X�s���$�\]���8H�Գ>wŮ~��l���q��4Al,�����l��O~�^�6�!�ru\��%S���X�J�HTӽ�K��7r@���M�Y�U��va��*��Z�\h(4�l?/���uЖ���tFm4Y�ǋ�Il���Tf�@�<��$<]��p^��������BG���OF����]o�l��4J�G
px�Y&G!���>�Q�o�{#S�^+��B�	���M�I�U�`O�8�^X�
���dD�k���Q�S����*�S+pc6�f(NMҭ��/�b=���[P���t{7�*hJbf{B��Z}� FFK�&<��椫˒�E��Ȓ W^��B	{�i����e������% T�י���6jK����{�5t|�K�W��p�VR����F�e�u<��wk�T�9ՠ�Z���_lu����_�\���IUJ�|���,o��e����!���u�����eW���m��I�Ź�P�a���@9�u�=���l�x �A�|'�Vk���\�V�FZp��Y !2S��;��-F�X�]�y���AoI/݈Lw/t0���L{���Ǣ�$�de����<��}����!�
�1�Z&�n k�u�����/sa)��P�Yq�:^��̂XTWg��al���#��L�j1��Y���2�Bٽ$5����3�n�����2�`����}%�t&�����f~*�p�R.�I��He�B��a����5�,�����V��+�j��p�<"WI"b�v��H��T�S���Ӿ���?������9��gn+i('����F�L2Z}��w�r�@ \��>+,פ/�v��5Xzb����ό�4 ����pga�]��$6��ҳ��]����$ e��N7������kHB����,o2$��\Y:�C�uK!!��L'�c�>�}f�wD�Q���XE�N�l��͇OS��#�Y�z3l����s��R�1 ��ˣ	�D����=��1���ז�[�.l��i"��E�Z-�:�7^�p�
��>3�\l6����_��g�o�ikOc�������*V�d����[���WYct����SUAlO��T�+n����&�U�D�=��\�1k�w�%���&-a38�X�U6�Wg&d7��\_ޯ)� ߬��/�V�F���4� ��ˣ��TZ�����"	)1�-�w$���޺*��m�/���yy�o�9��R�%4���q!�g�M��nVp ��xJX<���M$Cr�o�3^j�t��7�J@+ڦb	���dj~���h)��<HY�y]�=F�����_�Ru1YR����3RT��FP�"h�)�P����3�z��ܷ�^A���'|��`s�Y�g:!����sƗ�u��IP�
IY6;����o�#]��ř$�ZWxˢ%��2KF�A*Ru�R�m��cb<�+�A�|/����o��ԙ A�Xe�Ե��҆�wt)RD��Ƕ��n�0\��x���D�`��+sށ�Oȡ��:�2�T���k��%�O���g>�+t���0����;���3�΋h�ac�~��b���XJ6�τ��A[�Y�z��)$F$��Y�����0�7�����v�E�$�6�ܻGr�	�h���>���v���a�r�� �g�a�-fs�3���.��3��F!y%� �����GUc���vr�c���/����8�j]a�	�u N�F�nn�k���@V���GE�g����7M�c���wb�k�&ǒbt��f��ޞ��������84����C�-V1����H�N׽�F��o �P�?I�RO#�*�G`״i��cE���JP���.���2+��k:-İşr)s�gY�c4u�*Sb+��h4>isp ı>�`��&����]�um�{�a�S *�����Äe��U�ų\Smm��MѴ-Y��˯�K�5���Գ��j+������#�ۉm�,trtl��P���g���[atf&�N���Y�s��`MN�0��	�J��7���=��m^�N�ݺMSf��~�tO�
��t��,Q����W��O7 <@�
؃��}�do�[S&�\@��AQ
��7��(iKD�#�M�����9�L'�C��� �KGH��TU��c(��n�aZi�e"�[��}[g���#�7.���J	S/#ԓ��� y�H��䂤��2��ŰE$司���ۣ~�s�y<@cd��jsI.�I_Y٢ڏ�7���̅-����e����65HR om������2�}�j���
^h�|�/������v@B��� ?��^I`��� ��"Rq"S�_?Pf���6`������d���;p��3-fYv����\�\�o�c�<-��i��<�l��Y6��K	DQJ�&!8(�� ���.:%�����W�t�haw8�h���/3�l\�C�'% V�#>�PB�.2�{��`e�E�.�S"]��-���wL����ٵ�u�f}�M�>�])��.�A� �^���7T��+�"���k����g�v��T��y�jK���-:I|]�N��)dD?����"�=&��P�#�L&�x�����:�Wj6@uz�������N�=�<�{�m���8��)�i2<��ੴ�����A���/���N���_�G�?w�t�PP�pi��� QI��Zsu����ީ:�ל����[���8��O@q�=Eu,�%�KY-=,7%a!�g,�|h�s�4�� �k�>�1? FM�,��"�J�S��wR-▱��4��|��+Z����| &��z�I������'�>�������(a�[��ȥoW���E>^�#��o�6�H�==á���Xĺ����kV;���7��X��$��w�{8�����(pYNU���d��SsT��%�d.�Dxח�FW�ܖI�����r2f�z╻T�eܾ��q�i�!y�⮗��g�_��9�@�M���'8qso��m�a��7��Gc�<�.�����
Adۺ��΍�����0c~��T���gh`U؃!�"u���Ŵ�0�o.w��ωr�o!$�;T��J�\����(��Sv�-k�3KG~��<��e�4�҃��m	�`͊J�AM^5 ��ք�����XPk�0v	�yg�*�$;Ev�f:���bτp�~��Lnls�"�X�8J���a^�|"�>s$/^6�\=K�F
�<��?������}ȴYHngWi��T"�#"�O���~�(�V{�ƾ���d���$����荝H��fۣ�.���m���bƑ��TW�f^>:�@">��kT�i2e�9,x%P�,x�|<�(�	$b���Ͳ ��%�(���yݬ` !R&�A|��=Z؄,�z�j!���0�Z����a�h��1�j���V��tnlw���ك�4LE� �C��\mV�)�.[|9�!��B;� l5S�9��)0Q �>6����i���:͸:�� �$���/ �Y��g݆%�����-���l�������:gtΰE��}��Y@����O˶��G���۰�W��o'�5�M�tc]�z9[��lc�-0��fh�Ta�pV4ɹm�%,Ky_����"�v��_�T�� -�|KuFS����>��&U銶�j5C�g0N�)�/�R��7��?�xJ=�fx�gFmB1�-Ig���]��f���5̵�X�s�V�4�Ɇ?���1�1��'ӨFo�<��%p����eUˍJ��N mG���}7� B����7���1����s��N:�A�c�@�1$]P��h|
�
�^���?����	L&��	�
I����'z[��$�	�ᙔ}d���;{(�̓�K��=A�� �%O]9 ���Ø:R��3\UW�L����%lN9����!/ōK�\�ۏz)��M>��h;��0���h�H���w8�]�4��"Ӏ@5�8�#
H��i/� ��a����4#.���+-d��q/V9(��k�2���ʿI�v�C������6m����)e���=���ph��+����G���'�Ü�
^Ƹb���A������k:�3�:uC�V���'��c�z����%0h��K�js[��z�y ރ�ݢz%E[�
�H&��6-��&�,6�t�>Uܨ��.]��b�e���w���݅��H^����D�
��G�_R�L Y���Nc��+p`�6i�����ZU�I(�IX�:y1�W�&�%���H��C�"����*Bݾ#��l�!瞡���
=�0���QI��JZ��U1[��J�#ϴ�5�~D�/4��V�9��`u^�W����I�q��,��&����I.*g��;?��7D�gW(�"@�Zs�?�K �$�������{3V� �aT<"���G���Bf!���T�ry��λ�X�a 6CO�c��I�{ͪD;mR^��q{~���?������]���D��~8&����q��T����yD�����?Y�`6��E!(j�h��zCb��;��׽D��j�c�4��h���h�Y�XJ/�R��(Gϟ�tz�w��2QWd�0���/,�WI�cD�-ao���Jsр����A��H'�;)l߾ϊ�	�0k�����j�^3���Pt�ڢ!�����RAG5���%vg,9Y������_-n�����,�����6�x�Kk�b �Y��4gC?Ĩv~^t[�Mz�D���:B`_�/���@�����\��b���Ah���E���:��QC�]U_�E9�Ԁ�Π���f�`֗���l�S�n5�h��u�p�H���1l݅�g�N�0�m;=0��˽C
�>X���E��� �Od߈�ɂ���"��aQŀ�=�ap�s�����JZT� �s�����t$��Z6��~���m��.$�P]����Ud��[�D�h��D�A��Y	ĩnnn��"ю[����W�>��%/|��J�[%�(���$"i����zG�%�Nd@O?7��~�Ȝ��.l�� ���(mzO��$�7�I�����g%Gu��z��~,8�d2d�"�����7�	�3�Ţ�H�k g�q�R̓�6����l�����˙Z%^+�c(��5�����Ѩ�f��z!O�TY���%�4r�4���V4.�Y%�H93û�m_��Q���6BXh
����|W=����9h"��e&�
�gޓ�$\�gS+j��������lh���	$�$}7���-0����Ǒ���\���E��\RCG�I���6=�y;�y�m��*%d~�-Dj����o�<��BA��5��<��,\
�J1D��y̎������0�e�xP�`�K��~c�4K���߃N�rX��֜	P'�)��!	���r���C�w����:{��V=:v�<�������!�o5_� ��D���q��;5#P6�rz�M�i�苙P��g"kjG�Hk��y�l�oK�	(} D�9˂J�ܳCS	(u�����yKb�o<ʰ�c�w��3s̍nȿ��u�(r�D|J�!#Ҩ���{�����d��b������8=q��S����j��e�����#,4WK=h\!�A��B!�)S���o!��hGrr��� �h���<�u��E�>��dv�i�*����5�]�L�M�`�@P]�$��P�lB|��a��_3�̉dR�ؠ?G��xٻ�o#��z��L4H���hX�N�զ&CIĻM4a�:4�����n�3�8-A��`N�<�R�g�J���n�h�6}|��Qx�6��A�1E������)E��u�I���>HL?<�
8�r��r>���y�^�ހ�dam��w�ea�4�	��3�ܣ���%�8�hjl�cM����v�;���
K�n��3f��C��%�N���t<%��#�&:�-��y�<%�[Z|2���'�C��w�tԝPD���y�C���|L�{�7]�ڻ���k�tD�$	Sr8H
;��Sb�xn2�E�#�0p� �e�������tl�C\�4�v\MO�33�i�rfOe�z}��ml�]�H�*74�fah�!!��u��a�b���v�����g�W-�ʠ�>�~UG�V*PL��拔8$�:�Uۢ��0N\J��ޏ���s]�Kt���1p�� J#]V$�%�:9��䷴���o擅xq�0�����ˉg����|�7����S���2�	� �cIg�r4r
xaK����8���2u@P6]2ŀ�ѝ�
�X�����'>UQ}�TʩN�z4#&v[����!!0�UZF��Y�<�@r�K�������k�,¹I��!Lf���Vr��L󪥀wN��@A���Y����MdC��k���s�g܋GUۙ��(�Ô괿o���]v���m݉u�t�9�X�+wl`:�;#��:��������|� �@r�:}�^�Zv��]+n�q�XNVN`PU�M}��L����x�I;�h7��ײ-�f����J�
9�!J�GE1��- �N�S�I�H�@��j��Y�`�<^���\�v,�1��%�ݷ�]r?��F�6�������c찤�����87.�g���o����<A7�9Mr�Yԃ^n���/C
��|/oj��v;�
/�a��$�dvu<o�7(�:apX��S<��X�����<Y[���hQh��41��xuv:������<
La�֬��Ӊ�Gج��4�U�95腣>����M:"=/�)faDk��a���p����Ž�Z�ֆ���� D4VHq*����
�iHFf��gPE%/��!��Y<��O�y�w�m�wؖ44�d$���+ӡ@���-���Mdp��!�vޚҒ9�ͣ劏G=������H�������f2��Ζ}��x|C��JJ�Q��Ǘ�h�|�Q�[ʒ{��Z�ݸC.E��-w��n��@�HK�w��A��,\;kh]	���݅��@";�K�̫`tNʢ�3� ��*���Ҏ
�ΰev��4K�l�+�,7����Z]$�D�֧�^��hC��bizx��>=;�����}S���x���?C�M{5�%���f$�������{�x��!��Ҳ)AXK\�-<߹���"�����dt�%�g!���][c>���⮻�/�;I�'�Fȡe�ג��?->p�
�n	���]�wa�Y6H���<�;�I���j��>����
��89����N��.��ɃKF�<"6B��,T�4�X7ߐ�vs���%�Yw1Q�ÿB�QG�f=�p9���V~BfgV�eU�V���s#�8���fX�&b�����m<����4�D�mQ$~
��I
!i(s隢�n"h�R��?�<�9�%^P
�Ӣ�z`�����3��ZD?�5T	u�Kn�����
�M�sR���0s�@�'t	���<��X�4�OO�5ޱ��+�&m�B�ԜW������G�%y��|L$��̾A:O�h����t�����q�Ɂ%I��K���߸8]����3[,9u9_��U)�� {���1綽fBLZ���!/-��ϒ��]"��
�;d�ՌiIQ������k�5�@E��e�od=�����g��2t���̱ް����`��*���H7OHV)\���Wz����ͱjhtAX8�a�ڬ�o���^�'�RR184bo+-�mI�糃�����O���̮��!Z�9ٖu�H�a��,!c�^�@-P�C�NuB�b��g��E�BsoYJҵ�,�o�C��q��Y}�Ed�hq��Pf�[s���j*( ���f���`��9X���9�/����u��X�|�Y3n��U++�dI}�D�/!D�����2���9��C�Q�Ԝ��¿���'U*���l>�fX���4L�r6���uH�>��hK��ޟ��W/4ض�5����u�դ�8@2���sKb0�AZ!t�hSܒ?|A]@�z���5��ה��w��_��&�e�F����{��Sst�'"Zp�蓨�DY����T���ձ�t˃3U�V<�z��%D��OO�5V�Uy���!�h~��\Y�	BȴnPZ�)Fz'����j�g�|FQ��V�{lF�p�R�%Ԗ͋-��uk�k�m�Q���
:Cr&[|�z��Z��ώ��]i����mވc�;g>m�_������W�����A�W�҆� �Dz�cC����侏��-W�i<�v��1P�~�����?��	$~p�Y�jj^��hNm�Z=�{_!�k1�S^��r�}Z����a�H��9S bUd�*�;�oq�_N�|)�N{9�A | �D��T�y�zڊz�=���?�:4a�(�1��ID������^�3��Z8\��c$���L�=c��h���D�lX��@���������I��-�N $�o2Q���a�E)];x������S�J��k8�����;�G��6j<!��<�͞s[�I]��膕�p��岵�����"��;u�t}p?	��Yk,�(V����g�����9o��F\g'A�z[��Z@q���L���<���<�+�ȡ���a�P݇��Z�8�A$	�s(�f��9�L�Z]zaK��p��{�IU��������S&y�wGjʮx�2��>����4`3�˨�}�-��S��x� N��J�gן���-���'�\�Z.�ɿ�?��k*Q��[N�zT�ώ��oe�e��� ���<���^t��KS����/����BS�������)���&�G�f��]�d�_[��e�C<@Yc�B �����S��5�@e|}��i�ZQ؝EuNBA��W&N���!䢰w�2��Vf�B��8)�����[8Ӽr8���M�
���I���U�BX'�a�FF�4^KL�� cM��6U#$�^>Q=a���1�y�9T	�m��0�'�؈�tɬ�ol��R�z	���:�{�����H��N�}G�!�E��X���ń/��ˤ�q��%\�j��ѭ���#r�� 6����"����ڟf'���}��-��+��Ϯ�3m5�3�r�bEM����S��QD�	nuE)��ʝ��Z�lܣ4;����@���T�B����e��yy�2�����AH��ܷp� `%W���$��Xw��⺘��6(-�W�B:`(Ji�5�9�7��ï/!Ӹ/�,b�&���q��Xh�3t��I9��>
� ,�H<V�X�Thܳ�G喳�ߊA��Ճ���Ւ��z��D?����J�k�y��Oو��&*åCO���O�ў7��N�)Ϡ4�`�.f�_>Lb}ޠKb�˄�Fh��#&�Z�Rࡗnq�"P��I�J�v�e_�*��.\7�U$������� ;�$��X����B.�lm��"��-ӆG�&Մ��>��1�8��؎���p�C��3f���IN.tҰA.ڥʝ��P+�%Ďu�1�v´<��,AoPS�s�g�;4M"ް��K��R���k8g6�p��+ |t�:��N�9�O�SQ2��缚��[��ԙA���-pwoQ��?�%}����lWE��zyc�j�$؊��d%b��$�?�i|$_�r���ʔ�����[�σڐ �KC�l�y^�{�ޜG,<���� i"���# ����#DU��U��J�B�JR퀓$���r��*�[L���8���k�R�3�sF*�60M��'��uC ��Y4Q������B�K,��.1�-|�0�`w
!�;uHX�`�'�\yI�_^��������F�F�^����M_�-�Z��g�H	�)���ضVTLX�)�`C�R~��E� ��G�a��1��#I�!�NL�,9�_NIz�Q�ʢb���6@�c_3?�2C�W�hz��N=S���Q��dL��w�"���c�4u��]�Ы��[�*�i)g�Nxp�'*^3x���~'�4�'�g��%��k�-��g�獒����;��[�  ޠ��dŗ�l�'K�֩SE��>��!���8��F�H�ߊ;�w8ּǪ�J�/��u�
AnW�s��yP���j�^��8@N�2
���,��̊�t��6)f���pIl��٥D��7�.�O۬aM�f�:��w�Ͷ�!��b^�i#G	U�g�d6�L���j���SPJ<�z$�e��F#G��[	\a����>Q����U{I�Q#��S=�����Ji�=׌��i�ZzU6@z��{����kK4��׬6pLk�������`�1J7S�yF���ԫ�-90� 9�@O���Q_L�o�,��3�5t�	�「̠��'����"T��>
?Ÿ^��!�Y?�#�o�@��G\"��,p7Tn��*��&�f�!��u\�<�����?s����?���̉�Kڮ��I��F_^�����e��f�%ꍹF��2.08��6���&#"0�ˁ�<*�ԕ�{r
2�0]gZ�fe^�Zq\�`�LN�/К������ڄН��Y��8�p���|���ݖ���UƋ�D��t��kot�KJ}u!~;~=�_x�&����٨3d\���U|�i��s��� �A�i�`��e5\��m����"u�M8����'k3+��0}!�}�-�آ�9��� �I
r3 Ȑ�2I؏�1� u����-)(��(�(�o�*�W���sp�(�|5��`Y[��i%s���+�������/`�'l�+��?D�e
�&<��_���r�P8������C��BZeJ�ƍ�f^�5K�Yk��L�AT���:��0P�L׷�1��s��ח���������Kv�*���c=wx��V���Y�c��+��ʹ4bALsH �	�U[�(�l 0��Oǡ��ᖠ�~P�ߦ(Sي� ��ܒʜnG�Z5_�h�P�y�#�RۋZ	Z�������TkSPq�k���������Զ]����8����	{�X�ʌ,%kf�P�і�����Z>5Q�Ǣ��K��4a���6��������0F�h��-�����8�޿�oEB��14�(�x(��ֱ��b�'%gs��s��G�Bdצ�;+,?uO�l�l��&��UR������%W����=~֭�z{�Ữ���<�&G�`�b";�s���i����W-9��&p�Bv	��͆�,o')�ր�4<�:������&����;��1���Aş�tB����j�tE#?b��L�8F�����'�?��6K.~V�t�����`�=�l#����W�Z'�Ⱦ�a�'�����GuF����}T{��'k�5u�i%���K
��/��K�p�$��A+�d��f<��_��+�� T�Jhk���"�i�B��78�)zNY ���Zv��v�![��� ��\br�Di�%n����O���i���:-;� �6�h��s�շP�F���7�n�}hZ^|Lcaw�;z+:���qgM��w�/;��; ^�E���gL���~�&�^�bm�� tjt������O�[_Z���JΦ�)�����az{ '��8�l���D0[b)����� �Q�z{��Z3.ѮT������Mʨ@}�1{���Ђ69������.�������/�Ѥ��K���$IG�m�	�*�th;]R�`w�r��T�:�\����G���~Ʌ{�E��0kg��UF�д/��Qɭ{����
t���(�tQ�ɵqpS��Iݴ6�)���XL�ˈ ÄFg�(�Ù�}FS8QD�3�Z;1���P,W,���<g�������h�Л�#C�tQ�^��~��n���K_�Ͷ�D�$vSkS�p�n`�m�P��e�݌��c'˚��|�vdO
4�3*��D� ������CQ/�Q��P�7�kaz������	CmDN���:�T�T���YQn��&N�<�J����L��Bi��_L���]D'�n��8��0��Ѯ�g�A�3����kdO/��C�p�:�P�Ύ|�\�"#�%&9ш�*aBD���:��4�gy���L�
�\�NR�|u��$1셋AD��J�6 rf~m��Y;qS�j0�&�w�e���xZ8��^�8B��c}�k=-O���DǇ�o�:p[�Y�^#v𴞦�9��5�'��,����S�C�\��/���~���MPӣ5�鯵��Ɉ�|�9>���h����K('�֔����E)��k�S���6OTX����}GHB�3fo�~���`��S)�������A��kl���ES>��!댻`sH�-���^mF��L]K2���x��1��?���j��q0���]Olm%r*}��^-WI���4}���hw����{;x���C91�+�O���pd���?_�Q�g��Dn�� �!P�vL����W
?������J�?�R��w�Y�iJ��<��Cu�����h
��@Eu �+�	�6��	�w$�"����"���}he�޻�rL "$_䘗:�T�;�E���`^��xޏ$q�4���sō��W(p����X�k��|�xA&�;w����"����`�H͡Tz�*U��/�{P~�	���3��pW������т#C�rVp�NP�cRޏK�(�g�2�p��_!�����z����Nu��W���]gR)C��f���*� T���~��r��J��/2%��n�z��P�8n���:��\�q����V��
����lQ9�D� ߣc1<ܖ��l>���-@領/Ň\x1��{Yn��zщ�(e�\I2:6�>�V6@�m��[;!" ?�1��8⟬{1�χ���85c����\��E���_���1���BL��� ���毸l���k�K�´.�V��ymꎄj7���F��r��xs��2f&��.���m1��~(�?OQ����$*:9�V�.K�hv�/��=�秬#����2�<*٤po!�M�[k�����ɧ0�㽻1�9MY�Yﺄ1k������&q�c���}��/�#n׾�Au���0Z����I���=�ُ���P����%W���4;[�����m��Y�j�ͪf�Ť����o�֒����Y���L�"�\ 7Kx��I���@�6�9�hN�;��6�C�T�m���6��1�j�1�^��Q�aE��s�<E�Q̇�y���f %)�,�:����jT�4��h��t�6�I^�!�H�oI
��o�{c'�:j�ن����o@n��񑐬��<���e8p��oRUܭ.�LF�B��0d������o��5���]@l䮵�K�هV?�Ӈ.V��^��L�8|}�>j���V8�c����q� G�=�K�<ր�>�*д�L��e�r��M�jZv�tIz{p�T u-~��y#��G�/�{��^���u�7w�֭��)�Fw�2��Z��hb#��������=�yYO���2��k'�&nS�ggl�� ��_n@�ģ�+L2�������s872 	*R�	��C����,���&�$D�?�f�*)1�z�y��a�K�P7�`��>0R�Rg~����	�HX��@��^�kND���#�+�a?I�t����㍙�����*�˭�}A��e��Jj1�����!�H}@����Q��$ۃ��c�$r��'1��eH �Ќ,iG��cN�l86���U
?�vBs��\�� �5�dY=P���ak����[�����")��HB4(,���i���m�Cy3�/����ŐB:�_4��o��%�U�>��r��C}T�l������@�VR�E����j$���rx�b�.3�м\2�Uu
�3�h!��n���=tK]q�h(K����:�m�x0�7/%l3w;���<�&��ѝ��f�k7����y����8��ʉ�g�q��������í�F��X;"�8�pJY@��<{=�i>� L��:c��:��l=����/���Rs6x-2eq��� �.����m��'�㹠b7�5K����jk�����\GL���n=�y���/�h����w��������7��8�=�4�[�q��BO��\��p��T6���J*��\�Q`XA�nU!�0�ƛ��.��Y����۱
���.�$�.�6H���x��B���_�Ux�V�#B������yv�wNY�$_N���+�--H8��R]�*}n�g{S�F^�lSd�»�2��~Z	ZÄ��"=�h����I�ƭ�#�W�.�<A��
Z���=�7t�I}����0����@�~4������ZyqZ��G��_+i�L�2&�?T/a1F6*ai�{�s��K��~O��T�$��(�t�&ü���D�{��:���#d�s���e��x}�O����hU귯l�Ǖ�V�{A����Gjy͠�r3N���c%�ݸd�|V �)�t���Y���mK�Y�6��Q���A�*6��Ł���Eh�h��-<�p�І����<N�2�C)w0��/l����W�(,�9ۈ��~î(Xo�I����ı�,J��,�;u<aNq���n^��>C�'�M��h�j�ӭD4�vbE6�@��^�BO�:9�G��*=����ҕMȻ�):�G��r�1�GN!bBl$Qb��5����s��V�L�6G�/��b�c���GF<�)�'�7�82�Ac�-�;��)�4_WQ}�G!�x�6��b�
c+zE?���Jͤ'z�+�|Mؽ_�1J�[��R��kY<!��EIa,���y��f˲�Σ�.�,ߢ�l��l�u+�FC��Z�ź�݊Rz���xY�e�L�"���Ö�5�ָ�0��4����c�	c�r�쯥&��m m�xP�C=D�A�*�wb���X	*�f����fu��|�xg)�f'	G��`C���\5
�{6��Co��3�M�2�_G�#���6ɩ�w��ߟ E��L���Λ��k�$���Y�t�짺�*Cv������ij�ma^;�4"`>���^8�IW`jE�¿�*�<���}�t�S�j֖�r25����ǻ�B(a��/K1nػT'��o#��߁+���1ٙBc��:2��v���v�S�8�� �;k�Y�?T$�D�(���L�	粰#.�#=u�ɾ��}�8���-�Կ�+�tE�5�i��\'&W�{�1g/�I����}�;+�X$����\��a�o���UҀ��H�� x���J�~�������C1��Jm����ض8�s�͛�=�!�DX��L�(��g����ZX����	�=�A��������#h�<��s�#����5�m]��v�5����Q�qݶ�_��UP		��f�^�IF�,#?Qi�-��Քe�q5k�u%�Ɩ�B�.W��2S��Hn�jw<���R�����Q^���@+"�:T�_jK�peΊ�y���8ߐT�B&�G��8�D�<P�F5���_ .ro�`7�x����å&�6zU����rF�0[��h�ϧ �EZ
�tᲹ5H�1~e�(܄6L���m���v8���꟫Hp������!��ri���-�K�%�k�[�O��� {����qy�8��nKnm�d��n��θ�7:���Eئe��m�q�G�P���WSWF�YKS<���U*��
�����3b�,kg��c�Za�v�w� ��3��7��gѦ^��m#���r�������h���>c�u�7u��7z�0�e����K�u���s+�o��d퉞�TN'1`g��� )4��@����s��*I� �N|��L�B��JU���t�C�[�6
���H�>L�x����n��;�E�([�t�2Ȉ�H(Ϡ�M>O5�Fa��f��v�A�Zx}���;�M'8�D�c���V�,�C�+�ݙ�ؘ'�1���XdiF[�y���U8��s���Я6ORr��F�Ŵ(�yJ��\������>�d��j��Μb�zo��,D~����Q�jGO�Tɼ��Z%��B
�����_� �����;Mt:�
 d���p�5��4֎�9��W��4��9���0����@e�����t�r&hG2Z��+T�G�����!��u,�p�b0=,�%&��m�.������8Yޔ��g:/��
��n���5��g��]��8u��½�a�^[3!���v�U$���uX���<�$E���b�*�b�X�S�?'����\x�ڋd�<4ȴ��H��rB���k)7,j6�`ҏ:����{|;�������p����rj�$�Q"�2��C� T��M���";�^������ܤ�"������� �@2���0��o�mO�\h����Gj��ؙQR����DRh
e ���Ez��M%9ͥ�k���;|�z�f�5�E <����5
�x:G���m��kp�h�:��ӀCN:��lk�Ys^O��w������6c�}�\�l�g$�-k�A�D�X,?o���|$�Ug��2C��i��)��fi�E����nBIH���A?��ˏ$�j���`��J�&�ۊ�O<�9����ԏx��i+�#�l�zAfI@��QgpUzq��b�<y��y��B�AK Fn�2Kŗ�C�S�M2������JsJ�]�����ػ�KX�j��񃫳9����&$5�;�;�A�Ƨ� ��#�<��p��0o�q0���ǃ�[�49��<k����r�)����3!ԏc�LU���w'��'��d������0��&�d4%%���!Z�8�^E���� W�6��E^�� ^�o�	���%e�
��Hu_j��M�*�K<;�0t�,;�45�%~�P��ʺE��'ؘ�e�G��m�v��M��d��ݑe�0�d�"���l0G�v��aK�-cN�I<�,�E^K�e��F�d���;��	������_h���K���p��0%mЎTJX�z�A��!��Q�
EFя�\�%�U���
*�6� f��J7�7�)s����M�9 W������n��|\�Rc���)5[]���Ec6���5��٦�$��j5jYl$�d=�2~w>8[2�.���+x���L�ϓ��xW���������&Sҳ\���[����:.9��7d�ǭ�"ޡ"��h�0�I*��öwu��m�%v7d�z��B�dV���H7���y�{�˥p=k"s�grz���ha��*�4ʊ�2 f������!g�N������ n���/I/��^�r����X�!����-;k_�VޑF)V���
��
���SVF8ul�����D��{�����Y)Mld(�IҒr�����h)��.�q��
����co�n�jI|4��q��y��(��z��ƠIp��e.�t�<�:��H]�@�]ӭ+ �٭ʇ��\�$C�,Ͳ�!�NA�߻�3,��d�}�����kON�G��(Ӥ�4~�]vY��)�P~�e7}L��N�4V�Ȩ��w3�N1��ZVtnު�ƉYƠF�[m��_anYlyb+'��W\ӈ�ú�x�Kx�Mr�U��q�!U�AɁ���b���.�z�:'uX%7�	�}�U�+#�b�]
j� ̂~�
&x0^8y�R��5?3�?�zs�I��d���ln�BG��E����gG�
I�%��qP�d~'��W�eJ���<2
�s���J]�^�Ʊd�x�3�ږüg*�7�.rx��S�%fz����zV_�4C�F�a�ٵ۬y5� ���S�-���M�4��w4Q1MH#��ހU0'�&q�?.σT�5����Atd<PR��������e�L�\�%��� �⻦�0?ri�ǷsH�H�"<T+�(d������eiϲ�eM����ѐ#k���KѦ�Z�� l;F�M� �4��E:��ǿ6t�5�Fob��x9�̣*^5�rV}�7�X�,�h5+W�6�<���+,�z*�:�ɖ���߶�H�\p���Y�K�����T�󦪣�зAB�Q��M�p��U�M��u���=l�Hb͟7��7�:]j��̻`�]9Ļ�d��c<��e7oN/�IG��^�ԃ����/Aҡ'��38">��;��׼p��[��Ȼz������3�󶭛�&�?M��CW,Lג���_ן���j �flY��\"|�����[�)��`���a�B�x�1����Bs�!�Q$�y,߭zf�О愈����$���<�=b�㩦,6����#��u���P;x�d�N��g���Fm�v����䱞&���
��o�D=�l:��vY������� ����ʶ��@�E��U��r��}E7Ά7�DӋ�%�T퇪�'�+;�|6$�1h�Y����s���_��̆�����L��S�+Y���Q�#'���t�UI�\�ю�&�IK��+��!,��C�9�_ ��7&��R~n��Z>��;�IK�T�?�R3ن�~.=��n��?I>sϴ�;@�\�Y�i�=���V!�����}� �⍑ĵY(�5�����ן����!G��̔�Y��碭���n���oGmFl��n�ĥ��j��,��2�=�VY��_��D)����^A�]�WedP�t��/�}o���gS�m�`[6&D��v+nc��x�>atD��HΓd��ɪ�<�%�������SE���+�Z�%��0��)q����\�0�=
�b�	���/{���_��!�䄝��d�>	o�S��,�Z{���s*��TO/֩�E?v��:4�c4��BX�}���9�ǡ-�0�A*2�OН��Q{��]��[Sp2��ªo�D
��\r�Û�|���l��83�+��5�㵰�i�=;����C��#��	�;/���\�\R�{"�A���<↨�c����{��?�42��M��DqYs��P��L�ȑR󟏰�	�ɛ�)� 5�i�25��O�CS�ˏ[g�c4kTˮ��H�nPb��

W���꟔����
�`^+Nq
b���aPc�N�3��c������>k���ͧ���c]�.���N�,3�7K��p��M+���M��}�u�����ioS������,�I��..Y>�Ȕ��(Y� ��֣ ߽R�8a~HS�7�zT�}m���y����`c�i�{I筣Z�o���bE��+�H2V5�f������۪�Qz�'�������p��<-.�Yi�����P1t�!���H�I���D_�y��@v�7�K=�<�"9�|Ex��䙇y$َmclR
ފMv���_ct��0��+J�cЬ�qS
ky�I����Ġ��?X�� �.e.򯅻�_q�B5@h=깘'PF^�κ]P�?����>� ڍ��/vdo~�=�2��B�+]��&A�����%���F;���_���"���M_4W���c�^r�⦣7��nɎU��F+x-�p-Na�Y|�d��F ���i���y䝠�������i6�Gwޯ��S�o��p3F�tQܮU���է�ߦ,������Ԣ��E'��+���p��M���)F^O�G���W�Еj4-T�K.�<����Wd�9NOG�M�A�:%���TV���*tq��1s�ɕP�Sѱ��,U+������� �7��Ύ6:��0]��ӝ�T��b��١�L�Ui�4=hrx)r�cŗ�κA	��̼AA��[ �|��=G7���{X�L=]~"�i��Q�y�'���&�l�u��Z.nO��M�������}m�9�65��
UG�I0R��q��P(�"���W6�l��K�m���t-��v2�V��!w���ocdO�s#KW۞z$IF<�.�]߮�Þet)�?DL����5��nt7�`>7L�͔�(&f������'�u"gyK��[K��Y���M�(�͊�U�!���{G��E�''�4[���$�8Aa�HQ�|��Ţ�G{���(�{e$C�Р��̱��2�hQ�����IP�g71�Q�����l����)��w�/]F���2��PԦ�����(9^6�������x�5��(�o��!�D�.�=�ItcBW8���W���w5r��b<�-^1�A�
|�zr��-%�>�`[�/|[���Ĩ�Jd���V.~Bbdq'�a��YnSZ��(�d��X/��$x2��0��P}x��;L��K�	e�Q37�54ƚ�����i�=A�l��XGp�	�}] 8[����7$�
���C�ѦV苢�;N9w.MB{���̖|M���C&
����PG����<<0���\����;��x�r��R��18o���]�c�V��87�;FBJ�szD��:��a��~.hP��N�=<xK��!�J�7�vL^, ��}��梽�>%)#�����腑��b�.�n�x��V�Kk�g�Uf�`��Ư�N�����x�d5��N�ο���.�N.TRp�i �V9J�[����9%��=��_���4�ڋM���&w���\uݏ$[�D@'��\��~<��k4�	���lI�X3��s\�c�4�O��B��@ux�g��5wȌ���V+v���0���.Z��YO�$6TE�I�K6�'�'k�|"�2�(w�?�6�1Ya\Jf�"�k�����d��w�k�!e���W�l�M� *��g�WAW��?��<�%�{�C9�Tl~�y�>*}�{����V�����@�k�ы�Z�f6�*� ��)�� .l����Z��.�%1m���Ӊ"���JU�7�@m�m��\j�C����m��{6����lgX�Ѡ��$�?�&M��/l,�r����w�E�o�J�I۫��H�n<���Q;\�i�� ^v�.\fz�%��Ba��(%���wR �w#�2���#��ɞ���6	|~c�ٶ:�q�6���;�պ|���@'�O!	�A��K"��	�bהV#`�q�85��
����QAw
_|1`�Ǔ4B�Όj�2��4~~�%5�хD
�9��d��ƶ�4���c��J��)���|{�s�Kd��ǡ6��SxBٲ.�Dǁ�鵊�9m�?�H/�1��i����f��($����-�l�Q�|l�A�>	?�wwY���h��f$�BG� j��ر�I����ᝤ��p���#�U<~�b�����ڏ+E���Ý��w�C�[0[�ٵ�z-�Z���=ndS꾸��D&�Ƅ��.`j�W�-��:QC33�G�?����PԒ;��*/K���]�{�#���1���Ĕ^�-�4J��W���p�҃Õ���{SP
�P1[x�61��-�'��(�8~z�+��l��hW�8:�|��s�h"!��e6����A���6�R`-3�B�y�ߟ��P=�Y�0/h[B9;�, jeOw�޶��2OBM-�1?e�>e�*	Β�g��8�s	D/��n�j�e���I�MN	j�`B:6F�(�vu��EDo�K�7�S!��i�O
�f��9�Pzy+��y�*6�0v�-���c;G�/g�̼�׻���g����Jn#r��p/��
�u�Ҥ�ulu#,���k\ޕ�e�,����)�y��I�ͭ<ȿ]|⇒؎�w����[�`Xy�W�L��=�->��&�i1�20Jk��<���#H+,LMC��9�n�S����RN|�7��������H�0�R��a��Fs���@�(����ϧt���{��q"��t���D�i9+oH�4�) N�"$!�n�6u�4�9e���p�P� ����="u�O#S���n�=y�PS�c4���	u�(����+�;j�$.Ѯ�K+p�i�sr_P<UN[�&mȰ�W�/�]FWWA�Vw���k���I�K7�D�4J����L��A�.7t�~�̎C;��'&ȧ���c�D�ė�K����i,Z� Xn6�Fo�5,�t/��)5��+s3��a��&��;�<m�����α��Ё.b��\Ɛ�K?�2�=t�H�[�9��O��=<8S���p��e�"U��V��T�LD̘���iooV�t��@sF�)=��yB{n�|A��y�58�0���]����s�4�HV��r�Y�x5joFmt�|[Ϙ��lk���+�k��':~�Q$�U�D?4l ~��A��'}���Ȱ��A4c 5+3�*�٣_Ӆ�-�} A�W��V��IbG_��������$�<���X�S�+�@\Ag�G���<�`�S°tjN Yi��4V�����𚘡�.��U��1s���w��X�U��@f�;і��d�p���e�G�/;�yuPLN���\Z������V�H�>ߞυiq�/��up�P�M���)��5-���
��t5vͨ��)�4��%�q�*-W�����h����1�ؗHd#1X�7������
+Gf��|�MP�WE]$d����;�R)E���|t����6�h�1��-��s��&N72�C�C#EqA���`/�6�
gy����5����(�	�\�m�c�}���R�rG}P�m�@�������Q jں�5UW��$#���;
��Y̅�	�0sea8(+h�����7F���/PmM�Y�E+b����!Z���|�6=�H��]���u�c|7T��[���޼��1��2�	~,��ٱ�le�P?�n���R������@�@G��Ud�g��i��yta�����|2s����Zf��Y1��x)���B�fFU�Zҹ��a�0W�Ad�J��T>��g��8��n��.lE��Z/}�ݕإ�P�k��S��q�z��"l��c�c+P&���,�P�)�M�Ja�$����NEi�U��?q�?��Μ**�J7�7�����xd�R=�Ud��HS��A�g���-�}��{j?�6V�T��%���2�]���H�$sk�M�sDTq�Q�M*,�0Bdbg��z(�XL����$W���R�u�u綌_��ew,�[���,���$�T<��G{���9�s���+���w},bA�-��S9i����ԮS`Z"�?�b՘�6S�(��w���K�%���"J��.4�˜d:��Ӛy<4��4ޞk:�D��9�������V����B��]�8�_a�'������q�!���:������
C�4������}�7��\�䏻����NE��߫���pܝ�(����U��#���������e�w�*�&�yh��L���y �S�>�Ѝ��U�U�)r���� m��-B���& I����K(:u��,��{��3��Q�O����#s�'�_�?���ja`2�n笤��og��AɊ �%�k���w�"靤*B(�ou�ԫ�����#�IJ��?�j�o�;�jTSx�}�H����Kg�`nJ:$�}��~^A������րΧ°�#�����/n���)7*�͗�p��͊���s��os�;+� �l��s3љ��:��W�u�d/�a�aB��g�A��zJ�8&,:�?��G$re�^{9�A�&	WvBJ8UH�+���L`���I����`��Tȩ���Ҝ��R�cRT�u㽸�JZ�z$�"�#:.�f��1ea��-� �=hM���2��E����C5�"��,�W�R�IK�oBC��H����0Q��[�����2n��x�䦐_��f��B���Ğ�h���p��!���/ѣ�����
h��0�'(�%���-�� �.�����}&r>}H62H㪃n�O�W�&��1�ei���yL�������,�����0W�fv�\-G���0M��!i��v �(n^�|~��%!�����*"g��4��2�Q��r����6	��Y|���r�����|F�))8�:�(#@��Ò6���=�7:�m��j>�SaF���9a�g�1�z�Z�/Fy���x�S`�r�;��������?�t�8���Y�Ŕ,�8r늺��*-?=���������8���MS�JZ���$Wh����.x�t'�I@�^�Ii��x>2���n�E��V��o���(;�뙈����2��|��v�Q�xHٛ��˓�7S�����4§�n�)�<�t��'z�$�"�5{��g�/I�HB_�H\�� /ӽv���܏2�d�Ks�Ծ��l���h8P�}1��F�o���^�y�W�����Ԗ�qB�ŷ�˕�*N]���Flhͣ�#YId�!���q7lg�җ��4Wz-��R�����9zZ�K/��6z�[d�n�ݵ���C����c�>��v./�*'��ކ�D|�: OԆ�xJ�q����1����oO�pn�����º"��Ժ��Iw�e��ydE�G�5�N�o)�gO��ߢ�n,�S�^��XD[4	�\�EG���q]�N!+B�Z5_�hS�y�+����$LטZ�]%��y4��e�)��ҕ$@�f���%˂���zن��+���knH����'(m!����v�`������f�T�`��ڢ���n�I���o��nܖҔ�CAQs�CF���u��6�x�hȸF^��;G�-x�R���;.k�T_�w|E3�Is�!m�ϊ,�پa�����s���ωͭqrE.���Rd�|$��G�i���4�u��X�Y��?)�K=�mP_m�������T��*��7�E*l-L�ٙ����U�+-0'�:����e��e�b�Z��t��1�����7�L��{�>���-Z�};�{C��p+*�j��e]�Z�1����b��#l{x�3���@����%��r_Of�|lgt6�]W�n�`�iL乕��-"(L\�8��4���9C�sC�򓾋�����l�'�~��3y!�����b�(��p�>��+^u�ȯ>��P����|�,��9S��V+���r�<0O'�aP/�3=u6�&�j�!�˅��a�[��C�AZw��L�k`�m�R,���;]:%4���LDQ:]b/W��P,��[�>,�Qb�����D��tQ5{�NI�ИZߡ�:�����P켻i ;æ V�k�|�h�5�������*�J�;�q���# �*��&�k�C<���oOl=��S��L�5��j���Է�~j���M�l9����{auc1�͜�W`�G.fQ�l���f��qK�E}b��#�r��E�#�ղ{HOT�����ˌ��������悠Wyѽ5da���t�3�kK8��#�����eG�m���f�\��|�`�c�ؒ�Wf�Ƀ��}��%#�vA��S��,�%$�a���gk�9;��9�ʖ/ 9����e^&iC� �9ȴ���.5�˒��u���-@�Lqyz9s���)g�(��{��t}?�xH��{�˧i�����h-�\0Y�*�љsN�"(?m\N�I��|���T䔛foCt%�_k	1�a��n���tj�t'U�Rra��6'���DU��Hf�]֝.����]��"���%p��Ze"�@�|�/WQH���ӝ�вi�By�g,�P��f���t��#O�t'/âɧ��Z��݆��Cn��O�H��`lA ���Б�؜K��Ĳ��rj\���s�+e�P��-�M���-�{�>1&?cP��"{�շͧa ����Y�:@���s4�������SB��܅����� ���hw�䦌p��MT��g�N����I�����t:�|Z�����lgC���P_V2��dǊ�Um����T>[L��~���޽�k4�I�3�Zߘ�R"N���fR�4Ac�}}^z���67]��P�u]�]wQ�nOב���5���J��(�g���	�6� �+~�T �x��C ��aD�Y�;�_�9�0�1j����~�JQ�A�ǞN�1m"�B��ҢE�$d��������Mz�λ1��D��	�S,	e�s�NfK�C�;U@�'�2lU�&��=�* cN'dw`M�����\R��j�z����I�CM�ׇX�1��wY���uoHU�`�VW^���sEO?��Fv��Lr'��Z*���t���������O1=��mճ�&p#��mR5C��9c�=)d�,Ї/���5��+?�����*]/���nȗ&��CsT5�5�o��A��
��$�:�>pÑ����9@N���k	1f~��8��~
"ë(��Z���\�uL�-����%��6g�l@A�	N�y�����8�,��:�����f����7ǃ'���)d�i�C�M�L�p�Tq���H���+=Q_��]����
�ǣ�W��e_f��{�Nfq����Am��H�6�bq��wEF�lp,IIi 
'��`�G8��=v�kJ%�r�����HI`3�R�0�1r�ZUA�V7��!&4?⃾�{Ӑ�˸�D���M |~_&N�'�����zv
��'��~^$�p�����S�a�q��t�24�߲���������V�c�{��∄-���_J1�^׿�q��5l��󷀺�pۈO�=�ԟ�UsCdw@�Ք�w�G�ڽEmNoY� Ĺ7�G��ef��}bCۨ�2'���@��L���O��j��,�B��N������*�E_� ���k*�FO���Dl-*߭ס$���p�{:�-�x����ü7�{��g
pO+�$|q1�O�I)����(K�l�_�?�_���)��;�i���Z,?C�[1����������m�R�)ͻ ��1�e���T�M����rnj�K����é�R�V�ؒ=[6ѧ'�iLN�5��"���L��=�`<�H�R�f��|7ߠ({�#L��Zw:%o&��ӓs+-8Uc�c�E��E5m�{�����&��D��㵼��d|�p��!8v6D��+�F�˾m�wfJb��*gF�	 ;��v'�`����Q	���đ��[�p0D��O�q�=-e���#���a���7����f���7R���4<$و��b�{�	��IeH��|�E��)��xId#L��.S'���?�/=�_�#��"Y�0QF	���>��f��O<ӯ�kԢ��'{S�?��u���d5�C�v�����!��Mj���sBuO5��(%�[�zk��O��C��RM����x� ����_�~?�$�	�}:��w)|�d1���yUִ��D�j��.[��7�,&��K!&T�J�VlA�TØ媾�1��� A�S0�^�m�x�yD3+��0�7�_��q4���.
i��D
P�Cγbȣ+Gb?�LX�����.g�Tj����QN���KAO~��0� �@�Jѧd�F`��N��y����PTJp!t6b;h���Rh��J9d����@B@qv�pQ��Y�~�73��L*�ti3KTU^ۈ������s�U�K�����|hH����x|�r�8������,p�b�U�̴!����:y���/�n>&m��#�3Pp��0M��?�:�լY78E��רּ��$n��ud̅QTP�Ue�s�J/�6R�l]�k��
����ė6��ǵ�~"�N����H����/( Z�4������7-w���<�տ�8�t~R�r �u�_�6�����8kH[�&+���(�>�7i��J�*x�n�qhU����褣%��F	N��'����n1g��A��T����	������I�[���\0���k��j.�|R_�"ПA�\$ݜOp(���U^����Z�l���-i���Z:��(��J�u*�H�
��E@�ԯF�:C�uA-�v�ʊ�Z�}����܃�Ko�k|KA�`�}X)7��B ��--,�J�!�_�sufn���,���3��#˹�M�x�v�)���{LuȻH���_>��v*��"gg,���^�(oR.8zªe�|KE�L��V����MίWL��-e��l��6K�󤹥�#m�� �ʷ�j�j�^B�H�nI;�.������yp�F����͟ƨǧ�/��ݣel��kυS�<�M�DؒB�N�)�z
"�r(i�f	$Zex9W���w�a�0�)��}C&+���� �hdQ~J/2pV��l,l�=�aR�:�+�<��f�@fK�~ű�:%<�d	��P��&eSj�p��&�EOčL�QF)�dA��jU�c(�3�JY�B �(��
�&��^j��6(`��R��(�Ԏ�g��{�a�)\�x�Qe@�$M#�?��0��1��`��9o$_���a�`S��:�_�7}���%=��kO�e�b�d3w��#$eZv/�U�g�y���?W���΁H4��ʉ�P��_|�Ƚn���B���j�~���K�w�B�g�B��L8����}Cۥ�9�o�U�)�K��Τ�0ߕ��T���^�Z�cu�B�ʑc!S2J�V&eo�+G�����Ds;'�����4��L�H����G`�=	���'�5cUHخ�f���9%ޛ�;#%J�$a�;U�D���u3Џ��*��ЎU�.0m��":F>?�Y~Q0��-�����<�hՐ��G���t̤Vk��!��	<��ɗ�+�>Te��ڸ���Z!���L���H�$����{g�B�\v�@I���rp ��w�Wbx�C�C�[�>kZe8����-����D��EX>|m��CPK���up��ߧ�U��:����Xmh_�b��>��Q@�K|;NP����"$iuĢ��|G�<���rz�1��{�ϮR�B�t�.������9=�Ί�}�as�T]Qg7�c�D����Jv��vҎ[
�_�؛k�!�1���0>�M��,%}N��2`���?�ަ��S�t	h+1�N]V?���/��cw�)`C�wp.)7�����W�i�A�*`]xAW�E���h�x�/��'n����ޔ?5�2�a��u����|�!��3�Κ��G՛"��i�s�-��h�Ɍ	/�x���:0������:��SE:���;Nm?����c�h���yWq�p�	$�i��	��?�f�*!s�T�5�S��;����i����4<VF� �� ���_��e)6D�� ����s�e�U��	2��<��W��)~�"�,�j���rP>9��S��TZ��/������M�QT���i���
��8d�v����c���%jF�`3tA��έ��d0_?u�ߒ�*U�q��{��yI�lkAh�T�X�9�DV��&�sˠ�8��AT�,TI�Iڭqlt?�$���)Hv8�*���t��7_n���<����������A�s�<8�1���K�%����u�a��U�<
/����H2��^�2�]�
ԍ6�}��o���&3���������a��26�+i��Q�/ċ2E-�㴸p�5��\�7�h�*H��֢q>9�펧s��[{TO�9�������2˖�S ���M�O#w�`a�nO��ז�	��qnrO\�ɏ9e8!i_r}��! ��m�X�:���W5����xA���i��5_���1���n��mw�(BɂG�}��8��)�D��@�[�K�:���7|��T��A�wR�W��p�$�vBZb�R��0��e9�p�yN���.CW]����4���w�Ԫ�kTc\u�՘���>#f[��gY=���v��3Ai;�<�5AIB��7N7��/g;E�ؽ#�0�6�U�<.-�r�1�8��Jf�=�T��0�Iiz-]ݼh�nա����4_,�&HHͷϰ�r1>`�ǅk��C��GEI%�Q� Q\6T�h+��Ot]�"��B��E������B�'�A���MWƓ��h�[�:��Ĳ�m�{ޗ��7��A�}�J�1�2A�|R�<����c�������xC�J?n��虪�x4�����TC`T�۞�u�G�=�E55�Yg�>I���=F�lc&[����恋A[|�M�!�K�#N���Vl�S�[;���V��Gϭ��w�8+�v�;�F�"]�B j�;�0���߳�:+�v�����Vm/��:?�����8�Ը�C��|%���?�#�U��A��[�
 v��O����z�1�1Q�:3�bbG���H�?����ܭ&yĬ�^V$jLr�����9� P��L�Ѭ��O�����9xj�D������c�04O#0�x�����m�ғ������K��c���֞�8ݣ8ZV*��>��%�_�<��J^�`����E:���p�|��pT�Tm��ET�GDB#\�,�]�l��X�Z��$� 6�d��]ca�c�۩"J@Qs�.C{����)c|1���%���}AOUe�B窋�p�:"���D6!
���̘	<�C�]2���~��/o��_\�a:��?�I�1��d8��UY��ѩ�'-���)��T�IW��;BԬ�&V*{�	Q(���S�ۿ�x^�,V�=�5 nKS�,�fp͈8G��e@h�h��2�݃Ӧ6�w^ M(�f&�3R31KٺT*���	�!��-�1J�R���� ���B��HX�7r�	�Q
��E�͎���q��#��ZH42u�_d���7��5���� ���VG jo��'�Cү�Ǟ����-
��2(3��8��HB�G�4��7
���H1�I_��_*<�$�y�T��I�{�$k��lF$�����+��H��5�>D�&���a���J�#o����OP0�@�^I��Vx�x!-��$n�Ǥ-�?�ԘS�?8�*O��R��J<DΊ��ܑ�I i(ˁK�̕j�-��������V��k�a�L�����Vo_:
�'��S;�4`R,r-ِZ�Z9�7Y)����JܩL�����VTZ2����7�CJ�<Tq� ��f���!:�+o��\NlM�gA��Z�Bz�D���G*�R@��Kٕ(�e��&x�3yf�vWi$@��b<�3af�ʋؗ�5�����Q-� � �W���� C
K��M@o����)���S���M�	��q��0HT��H
�)�u���Fr,Śl��&��9�e�t�	,��t&��`�� �o�<��5���to>�J�6E�Ke>A�#r�_2sJ�ZX�*��o�1'._�Ş���`+�Xh��0k2u&��O�7�F��v�K3�+S���O�8�N�����x]����׮�GV�npv{P�#��,�[���q���<s
�l;���/�U]V�K�����O��7��0P�`�h�J�������M�^�rqJ�qЩ��2Xu�T@a̒��q�h��r�-�u�gz�ݥ�.-]�hk�u�Cl[|�Cū����K�L�6p�R��m(��T�)�q;a]x�z��	����S�kl��^����LSh�=\��`M)���k��^IQ�(��ؕ�(E��x.J�`Ƴ�*��c��r�Ol�C�{lH�gsh��qf�O�
�F7��Lg}eٓ�j��W�K�m�O��H()5#ؗ*(CA���e�J�)���$�~� ����RVz�����lB��1R�N&�T*:r����u��M�bӇ�������1��� b��{&��OSw0�4�d>0�4~�`W�(Q�ʼa��f�s�drFΩ���baQ`X!�ѽ N�(�\���Hh}몇�F�	y4�z����>VoB������4��j� h������)A�䷙LU�0��N��T�_8;chN��B��Uh�O9-�%�ٮ<��!�G���+�]^��&qL�ʩ���1�_���n�����Pb��Q|9��v|�
�����˯G|���~����$�'�(84Y\J�m���%
�
/8_B��9y~�8Y�����;�(Hq�-��F�'���AC:A~��{Kw�с�	E�k�,��tܒ���NZ�I?��p��Jdc��E,����S,E����g�b�L��bi��C37�bxAM֐�wQt�[��8*!qvFh���.�����L9*jQ��E��v������R5LT�!�,�2a |�Fwyk���a��׸��Ƣ�G�fz�1�n.H5�9w����e��:� ��2&�B�_�9{j-�trǂ��*"8T��$�c=n������,ff�ZM�)ע"g�<��|��s�9������pT(XG�Ǳ{J�Z�\���mI'p* ?#��C�+��ë�5�E\�Rp�2Y��s�]����B�{�FL�;����'�� ����lu�a7~�/m�7�o������+�w`f�X�+?��貹�MC|Җ���4��~�,X�Ӗ�~n[�a/����JÖ%��<�O[g�Y�>��c�Й�ט��WyL���}A�����2h�2%��_0��O�����י/G�Ժ��-�8��f��e(Be�Ve�5~��s5%�F/�Nl=XN�2�m��/������N}l�Am�	G����F��>�r/U��7�
	��̵,��YH7��LS�׬�B�����t�S\�*埵��73�M}���EFd�l6�!p�/��O��6A�,8����Q�VP�0��������U�9�����=�RL���Gh���Df��=�����/�r���[��7렳G��v׹��4���? �h�x!���~�%��;Vo�9TC��-ܠ4Pև�a~���A�TMֶi�@�@h���3��C?be�u*p:�f�#�Z;ea�[G~b�wV��K�B��;k��͍�~�Y�N�EƟ
���ڲ�̉��&I�U"^�d�)Ѧ��<�q'������H�K��;�G��;/y?�y2k�-m�PM�����i���׫��ٰ�߻	�xI��[x5��a�g�?�dDWeu��-ҽOo�WC#�{��a�7g����T>�V�1i;���{MX�$���0%4�3:$�D�G��%5m���X�{�EŋW�ؒJ�5���wӆP� �^�6s��)�
���e'�Z�Z�p�y�D\q�-�F���K��-�S�`��D���Ŋa�Ai}�pR_]������2�CH._ ���_)�0������&7"�b���y�.UQ"%�m�I���X��)�$y�>�
cD�5�io����%���z��i�`�of
�m������`��Z���Xa��qk"�����B����C&�֛��C(zS����V$R����	m�2��R�x����lҹT[��4Z� 2ȼ5�,��7z�ys�E���{�k:M	<��zة��=^�9*��(�V5��+|�u>�"}���������&)���B�OH�0��m%į/TFp�M���,z�ݜ���������7R~ u��_.�~�qe�����-��Y��, ���u�5���W�<~,�w�	�����R-O�Ηx���/��K+�-��/��;0�V����5��+�X��fl2��

�ȍMpE�C�c:��}(''v�� J$6\�:"�9����3HX����L��D�s q�[�8ƭ��y�V�A�s!{�Y�g�R�rz}Z3(���p�~>3g@B�w����,���5�K����)�9~E2�3e��+\�O��_�S�hɯ'Dl^��y�P|�K(�K+�?R�o��mښ�Y$��<��w��ޝ�wO�"GqN��h��I���N�^(GC7�3�|X�Od]9�]hQ��NY�^� �o�?oh,�"^��	9	�r˓M��%MĚ^�` z~�~����_�%95W�)h��Zy^���og`g[�s��׋͕���J��#�Q�ղ�ܰ�L�W��If1u<é���zֶ�LU�F�Zzj���)ٯ)+K�c�ہ�� �4��r�����fg̎}"}��1�&��[#�WV�	=b9���x#�����֎C l1�U����n.u	�k��29{a1�D_��9��w�k�]�~W��o����@���83'��P�3.�Z��"�`�NOjEcvR�~��D�y�;�M����p�ˤt{̴�sk����t�G�n���̄�=S���S��ڮ}&�g� g��z��'O �U_6��;w'�����"��,q��:�]�@���:�P���f���t���f)UiJ�G����x�+x6{�BPy�}샔u����E`p�Hdq?r����t'R`��"�E����(7�Y/�%H���<2�(�wؿ =Ԃ�K[�/~=1=�ێ�Ʌ,���f�+��I7pzX<���=��PV��_��Ew}�S&XuH��Cא�@<�
���#-�gn~��A
^	�s����υMFJ��"��<VL��'�Oͳ��۟?�N�ו2?�O㺜��@CD#ּ�+P+��	��L�"U*o���HBtzN�>�h��Zh��o���㲭�/O�Vn��TmC������k���F5�K^<:�؛|#je�	��R�*�J��U�[�, �ؖ�ʗ*�ӟ�KH����}]��fR1唃R��K�o1�'���*��l$K�o��߃6��M?�ν�x�'|����cB���� ����y�#�#��=�PW�Y�\X�Zu�e:���u(;2�!	wn�ED���Ml�����*��yXʫ�g��>�G�`��k�^j����.�9C2HP�\��0-Jx$Rd-�Q�`"�a��B�|�;�?���h���)��5�8�E��6���"3�Ŋ.�.��J�xQ�6Urm�)��j� ��@ͼg$nW�X���a�ZG�},��Z�'��
�/���3��:6��')����-��Ms���]�A�Oζ1%����
7�`��~�khe��>H����~�yw�H�n�	��}MT��	Ȧ���%�_m7�B�5Vi,�0�ED���ˀª߳�b��\�#���e��EW��/G�t@�@�B�ꋍ��#Tx����،� �IA�, �TP&��S��� ͮ���Q�v"9�;���'M�u>r0֎������1���lꙝ8q�6F�̻i�6�~����.�:�	�Rx6Mu�ZN��mc˭"����=�MniFɏ��5�\9A;"�$�%@��E��1e���[� �RٖR"�.m*Y%8@�%I���w�ޤ>��f��b��ZR�U�$AU�i2���W��]G��g%l�8-%��i<���gΪ)+lQ����{*��W%P5D%��%���Tf�����d@2�G�=jW�,�ZLyl�k���HK2��V�lK�P�u���W*��I����Sʔ���d������J�>O0�A7n�̈́b�Q!b۔}�����ð��N '��I�C*��X~������w(��DC���_1��y���'H8���a���a������))~ڵ��f�,�ꆺ�,T is���?�mJ�1d��Ӑ�<����3YON����<�2��#�=2������"���d�h�����m��>�%W�������|�,�K�∐�M^Q|�<;'���hX��+V���i9,x�q�f��$KYzp��.��,��Q%	E,��v�1�3vɫ�-��!Yrh�3�X��V�$d0Ӕ<㣩�	K�ĕ����%�����-kWd��T�f�E7�R�a��b��@��O��Iu`�7{Q�t��Ì�:���IN[��|.B���&�Pq��Ԝ:b4����&�#)?v\�X���Q�7��C]9����w�	�^�L�r t�":�;�c8�Q���dg��uЎ<>2�zO	����@���eޔ�ׅ��1�����8]8F�_B�c|/,*������̲�\�:���`�]�2�ڿO<�>��9tZc\X��Z�
a�6�A��d�l?u����D�</O�5腝��q]R)�m-U$�>LcՌ�J�A����!�������B1x�m������(���]�[p�9�3��ʐ�k'�6�IR��9�"dtt� �;�0�+��^�":�+P�N+�#���xz1��))�& ��#7v�C4w7\��n��W�[��x,�����/lq��N*���&x��" ��Z���L�����[%�rk� �\F�ޟ�UL�<�v��3vq>���'����?�HIX�'*rL 8(}̓��2�JNL�/)#{F����m�:J�6.K�Ԅw��۠BO���өF�a,���9vcj�m�|0oq�ܥ>V�\��[�l�������=���qx�QJ���X��O$��Y�ۙ�~ʳ1�إ��ˣ����\N.r��΅j��ɼ�I�?
��o�������Ӻ�P	q�z���)� ���ɳ;�**Q7�C}ĦJY�'9��SS��W����nϥm�H�FRo����*�ea_hRn8j�߭�f��o�@!oQv�}�,�b)t�r��&��$J�F$�uS�+ҚO7�I���^|{�l�'7�sϾj�݂�!��o���#�]��KS�S6�'�8a�C~�$W?1�w�<����".p@�����M�{a����������K���6�.7�fl�W&}��G��Y�ǫ�ʁV<-p�ԥ���%�\Xu �c�Ȏ�î��%7(*���B(kLv�V -�J��J}�z��M�����7��H��"nFOS%�4��oM�8�lJ�xzU�<	��f�0�)�V�ov�:�P��bJZ�@�ܝb�H�4�]�>����ý(�uЏ�bl(� �í}b)���2��͓`�A=0v1�)#ٱyX�Ĝ�蝔B�:�F��Z�jN"p0����͢\���ڸ�K���ty������r��M���fN]t�}Tp���?�p��I�g��lAٰ���"�QlL�[x���d�a'g���ې�&i�٤:�N췅0u-�k���wW٢t UZ��ѱL���	������<`U1 �*)�w���;�x%D�5�gfb��HL����ۂ��7��W��1bf*�$�g��,j����x�t��ִ�7GD�>�"�O�T׽%�����X�"I�t��{��J�h6s�G�1�a)����s��	oTH��WY��X�^MR�T�#'�Q�Ja�ޜ��m9@���5��a\�,�����ډ�09$���j)�f^�+ =t�/��h��N��x�^$I��ل�nh�nZ�J0��}l(m�m���yqO�F�&c?h~���֨2X���ʁ�R�PE������z~�
¨+J{�ī�// �Me�B���"�^Ԝ�T*�8JxL洮�7�=�DUd�����K�JL�����.���鏲�1M�U��b�4>�f�zOy�J� ��O�x�e����hi�7�4���BhD�.)�W�2���8P�#�Z�`�zX>�
ƅ`�+�G���
��j�I\=�$W|����*�U�b����A�T�;�̑|���Ӣ�4{�V��I���V�/�<�Q8�jmN�<)����Y[��:���+�~�ң!�%S���J-i���-�2 5���{#h�]�(H�_�H���K�֜�֋IK;����	h�*�C�e��A���C�mj����0Ė��*۾���5�R���������hBƏ�R���BJ�g��B���c����Ax�C�_O����b̜S�����r?J�����<l������ ����P��LǙA�,�!�t|�?��Ң�S~M��"�J��F �f�-T*nR��f����z���}�Rǎ �T~��.*W���x�QS�����Cy�����o���i~�hlWo�I��b�O""������O���h��øHoS0�@��xqr��@��) G!�S�,j��3]��[� �H7��z�ݶ�<�oLw�*�(���[���G�	���E+��!ZaԵ:��	��V�n*�N���/�1�~C�zc_>�M��UΙ6]�!�(N�a��C+%P��QjG8�1v�m��U��l� ̦�^ ��2�>�}��+�����e	�ی= کvb-�4?����$� ����'a~2޲��MNl>�F!��$���\�z1/��xie4,�K�U�0�z#}b���jo�J��/�6��m ���(.@�U�3��qԭ����pQ���J]3I����)m]td>m���M�S����vm;�ۑ�{��lK���d#a�6�.`B��HQ)���i�&�~���W����ޡ���b�ᑜE�
װC^L�4?9��p���~�9*Y_�o���okA��_r����B14�`�u9��!�PyJrQp���)�]'I�Yƙ��6�{9�,�q��5U�V��V�qo�R~�rw�ג�xRt�^�FKd�7�:6^U�aD�ȟk���p�l4���4���8[M��GL��J���ٚ[�X�s��^^���e�h�`uz��²a���h��>��F(̛�ޡ�����gZ�\��e�}���Ft�'b�h	�6A�,��*� {m�I��<^���}ĕˏK����Mr5��7�F&pO)�E]����\�N�B"<�Cݽ�J�����jE 9�40�Ψ'*ZVҝ 0�{+�����x���x�D�H2�y�_��<�T�a(0�7
%�v;�ۅ	i���4����b/�ݎm�#�Vu>�.�Pot�$y���V�WE��4�_#Xy$k��@8�=V�SdyhSm�V������=�Ĕԡ��N�����_������:�~�hA�s����R�C��S3���w����U���,�]D<T�&���Kj��F�t�s9C>5������+}�]m���7D[��4ŏ���������%�������_<���kXr��L�}�4��kg�`!��T</��YF�]�"��N`7��.�;/���	O���|�dN8�tB�>HH�����fB%*�/U��K�R�K�y��@(��W�Ǿ��dq��t$����f<�T���=^iW�}O&�̇�/HhW�s���p�r]�\bcc��K�ln�e7Է���w�E>Al��u|��F YQ,� 7|<+;g��w�hyQ¿�9�A��j5���~���"���� ��l��o��^1ܧIbbR�E��5Ε� R�	E@���ڽ�ّ�{��ơd&����E�)�]�i����z�Mzz��4#h��w2����Zm�_�����Z�p�\��5D@�0�^v��!�z_�,��M!�I�Z�/��}]V5��P{&u�;�z��k�@W���[c1�pY9>'�~;��r!����X�
���y�w^تp�-D��;��3a�J3��Poc	#L�[�'m�H�U~Ccġ�/�(�����	��7=�u;����_L��Lf�C�
3�x�˔�����P�@��$|?�����_?��Tr��7��O����F%̅[稭��� ������2��L�����q[�a����~p�h���;�k����hx!j�G����d�������C�ĊI'ٴ�1|Du �ۏ�}y�� �LޥH��K����:��I�h�A�{L�����"t�������M�O蜲/�����z�DaIHs$8Yg�V��:4�-��J7jM�a��=f�,�����W�3y#q�c���"X�,���G�`wA�||?<3���vV���L_��E8���:znP���H�A'��G�=�}���M�dTn���9��D��PzIvf/U���]ғ�w�1��.��ePOx:��Z�L3fe��R�L��3��Ŀ���>.�l��x���<�jؤ�ԫ / �wbM����li{|�WE:�z���&t�AOK?�\A���/o���⹯��-�A��j���`U(�����G��lt�h?���e4�g���4Ko\m["�^�7�p�9��:�/i^*�}��Pꃣ�QȈ)N6/�
�<��ň8y}<���N���
xP�2Ĵ��r���
�͂ɱ?G�	 ��6?���![�on8�5a��f�xPǓ�B��uT����d��:�WW���8QV�L�,1�٫I��V�r�˳��9zXwk�'ym��F.�z�h��8���[�1�����������}(������96�|��Q�N��ɠ��I��<�]VR�2���x��Cx�)B��������@#����e8�u�^QԶ�~���땧4�wD4i��U[�Q*ª<,�}�U�D�r���t��v�L����|B����fCC�����`��jc��X�������Ys������e
~��)��:��
�l�w����F/vӯґ��_�iV�%b��\�C(�Q��$kc$�3l�{k�7��F�#���ؽr|p�Z�,ش��['�*u�D+�-%j�V���rU��C�z��/�N0;fE��]�^YfA�	�]��bU�0��6����wR��c9@�hsSU�_ c�W�S�
\�����ʟTh9MW������"����A@�d
���F���.53���7�k�R�r�0���-�L��{�G���O�U��3�V�2 '�%m&O�(���xE��"PHnނW1��bń�o�z���ea�+�I��x)��������NB�._YV���bMۘ�i��7|�>��7^�+������!/��u�A���𣣗�b�� 	�p�7WJQ�������d�ˑ9�����S�;/c�4���`Ϋ��UIv��c�ug_氏��vؿf� {q0ď�9E��U�tUj������v{f�����k��{򕪵� }dq�E*�ä��}��������V�xyɑ���"�ջ����"��ȍ���I��[6��o���R"ueP'��X�#�&���a��vl�8f?���Qs&c;�� ��Λ����J?���OGoL)�S�`�a���[��~7G|�p:�'j��x�r�hn{��ؖ��M�H~ޯм���<s��'/"����r��������(�3k���4L(�]�G�iT���"4��F��a;���V|�ǽ��| �P����ωv��e%���\t���Y?(��������ñjJ�vm���*�(�_����!-|�	X��!�I 
���4ƣ#�a���4/B����6FY�oA�B&E��z�w�����a����i�Iv��i`���]����[��-N\/f��bШ�S��6!V\�IR��<�l�w�|!�2`�n��|W��2�@$�҃(A�A�}��j��Kn�&���d 7}��k�t���gnjߔ��cb�||$�z�l���L�Hi��y�b���d�v�j��Ȧ���fhsb���O�n�di�#)u^�nx���\�[P��u���i��)���zQ��+Lx￣��=xJ]��VY(��R-��CZ(�r���Ȣ�-��G�N9k�K���p�xܒ�0�1���NTY�1�@X�'(�F1��%��\��f�5o[%i���n�Ԓ�F����l�$+M� u{�ņ/~�VY*�ݗ/����m�wt��J��,��b�l`u�N�V�OӬx�9������	`k_]bc�J�����A|l���dR�p�Y�����&&'�n*m�������8)��ɍv��}�j�;�3��Y��᠁h�+�h�� ��A���Oo3��L�W���
�]Ϫo�V�ˌ�[�����\ښjwIi�����k�6�z�$��C�J�4v����k5L@��lm�j$�̂)�L�±��H]�&R�V<R�#ef��[�;L��eLH��͟d�z�UO��ieUw���09��1Wl9Q�_����g�ۿcS�U`j��-���ޙ��(���Ҝ�̪��Q���4���ɟ3�ȃ�p�'b�1�Oa��F`C������X�"��������0鶄��)�~Ǖ�5����g�	�o94\P7�-(ҪVs�Jߢ�&�Pk��`Q��nT�z���s&�AMs���
��/�{����a���\�3��(eC&*�EI�COJ8n��X��Y�������ʗ������F8M�SD�(�H)��	U�ٳ��P~]������o���)��G�Q�D~VSpD��1�$��ŀ,O
��0�RNE]��.5�>�3���u���5�{�"��0��S!Ň�����:W�:]��L��>~���]��	q'�E��m��㨍��T+�#a������y�.4��JZ6�֏]��'��(��i#>�h�D8<�8�\��Q�%b*u�a b n#^f��!��4(j�����`߁1�CԹ�T��ete?��]H��I�{����~��f��ꋮ� x����y	���@�#��%nѾ�n�*��>�)d�k��������J9�����M��N��4�6��!�/�8�$���F�`���i���	���"9	:Dm����"j��	͡�Wm�DH�H$�����Sn��D
� z�+�[\��~��ʰ0uB���7�
��0yW�_���V��p���:���)��J��x{T�n�} .���>ۆp?D��H��տs_�"�dsѴ�kv5��՛��ͧG�٣#�ɹWG�TlgZ�f�����z0��^��e����b��|��i�w�P�=�g����Q�֯����@�R�>Y�N���M�`r��=[�{[����v�����H ���9N���}�^Qh��٫����V��s�����~)�Gy�ɠ�OK��g�����W8S��;.���P���t4�Nۮ<Aا��J��z��|V!ݚ�	a"7��M���1k9������2U�MG�Sh�"PV�jqT��CM%,gt� �6S}��"�x�uRo����8���I�!dHp�E�^�iB�q���(��$6�|�4�����K��O���}.[�>m�<I7�)*�Z�)�D�X׽�E�K���!����{Z��񫸿������)���QJG6M�(�%&Y0�e�2����G�=c=}�̕QyT���tڵ_+Q��8���l�4�Ư�6�v�8�����s���e����C��8�p&>bA)�T22_�����P���^@C��=��cF>���>�7ǄCH2�n�@;/:���|��R�Z���<F=���E�ϝ�ًz��}�������|�hJx�1p�4�A~��[���~�B'����y��) U��386F׆�-A���CNh�~F1�pr@oDf�l��$�<���q��V��6������|P 
g�PN�<�'Ryî\���z�Q�O^��' 3�8��0Q6hD�RWƪ/�C���N�}H?�}k;��z�Ɲ΅�'���n*���x�b�@^��7=�!�v���C}p�4A\�0Rt��<�����h|u��Y4HJ&syO����e�t�¾�%�B�#���[#�f>�d��I���<��ޢ[��@QW�Ҳ�����[+�Q��&��8$]V�h0�5����F�ګ�'k��H�t.�U�d��@���Bv�3I�٩p9[�@Ҫ)���`"��W�3�XI�mMӦ2-!㗭F�F#�F�M�Q���]���g\2J���-+w!��������&Ig��;z�D[_� �[d������i*
�H�鋢j���-���j�g�L�C|o�"R�`ד�|�+tL(M�l�}�����N���eE���`
�ob2��'���t� @�Sî��js`�V����W M57g�QTS��&W��EԜ�Ts�_�
2�W^(��i�g����-]���x�X�5V��+���B�����1�Ƌ./�c�U��b4s�6*��c���6��D|��2F0��=p���0�vmI�Ǖ
�}n��)�4�x^�x�Iu#  ����l�^���t���g��BRۋ��6�LIu�tzg$K�n��Y��	��R�7mo� ���d���np���z�f���5��u�\?��w��DO1b?�t��iz��b��1f�������	ĞJ��S4���8mS׋����kd]�Qi����q���ߌ�" 1���qr3&;|��{W�;��^Yd5E�KI%�F�)>8�ه�'��W��,|�ؾ�6}7����LZ���دܡ�j8{����c��lm�����$�R NIk�V�ʎո� ]D�A��Ta�=]�����;��0y�)=��wnPW��=���\W�� �1\�N��q�5���P�Tob�֪�:����tp����)��'�^c����F�y�B����X7 �*�jb$D�K��(���Nno�%��=�dD5���0�A�|}�ݼ�E �ݴm��f�+Z7u���}jhI�;n�u�k��E
[���P1֪����K�T�ͺevJ���
�x�۔Rj�ث0oDDL�h��&��9j���I�YIB'a�lEơҬ�Y�6f�A��'}��k��](�|˷��`�b��GY�7�[|k�\��ܓ��ULd	�LoCty��չk�ʊA�����ș��2wu����#�ơ���Ȃ�ٔ�0���g)��f��e����������I��>��b�|&��/�a��e����b]�����2��2v��&���4�^�����)��V��wS�f5�I�
S/h�5$�@A�� ���SK�'���LQ ΅�+�d �6v�n/���1���k:R�O��DL�=��l�L%/�o*g=�g�3ş��&{�C�t��:��;����R�1Jl��&���>��6U�0H�����q�7�G�����K�!m��4I�sB�v�!H|����#� �=�8:�W��FeN���{
=hiY��)}�2���6{O�h�M*�����FX��6v {���۶�YSHz�K�7��y^]1��3�
N;�V�Q�H���F���?j���"+s��NuDekcmPO�%��Zڏ��gϾ�*�)V�鲽I
zѓ�˔N`,G�;5�K�����d$d��������2K�4>�/�F���*��f:+M����pYӀ �-���wEr�LH4��p�b��gX(�tX�Ǉ�Ŵ�͑R4xb�K��E?�Ԧf�?`#A���n��_��zh~.4{���r&P]4�~���V}R��mW> �}%��� F�%s�����,�������2�S�Ph�1iOx�/U��<E����|����`�0�4�1?ᘷ���	�[.H�=�=�����F�L�":�Z�]o0fܛ�|��}���l��TuVd��M۱SUxd�,���&����gŚ�41�݀��j.���h	|X<45��D�|0���y�a��n�e�]�ꆋ5ቑJ�(u���{C�)���m�#��/�A���!�M�r.a��K5}$㙛�Z��=��@�;�k=H4���QR���|W�� ;B��bṲ���0xͼM�׃3�ڶGZL9 w��]�(	�Lݏwئg$���I]	��"#"�P�Q���SǼ�k�~ ���8<�g����~:
����IH`��`�8�`���m��)V�Z���PF�CJ̱4qVK�E*8��MH��hyUD�Wf���g��\SשP�E�~�B����ժ����g��}R�`�x4�6����N"��{Z\o�$�WYu��ۗj,뢿١be�Tyw��r@b���+���A ��O��1��k��)�o�q��0х&��թ�;�jE�S�H[J���� �(�ʉL.����KՄ�\q��"���u}!��g*�1�>�^=cJ�<mKǛj���*6��|a�
st� V���o�|��tw+�,�W+�
�����'�d/+Kf
�i�M��Upܽ�~$4;2o��ާ��F{ź�V�D�����3�ߵ�Q�e�����9����ˁ��e��̠��܇�l�)Κ�l�H SX�I7���I͎��P����U�R��巉Ɓ��w�T���u���u ����s��	��em:�km{�6����F��v�w��[���/�͗g��)Gr�ky�"Ex�6t'���߆F���U�L<�������$i.�ʹ)�`m]b'��O��j�x�1m�o��\���y	�9׉kQu$C�fQ��_�	z�ҩ���]��3;�agM�����H�!��C�S"��WF������p2���dY�^碌�G�F�@V}�9�)j�P��P	 �	]d���nR��9�0�#����H�ds?�xj]	��O�?qLҠ�E���>|�{~�Ϛ�y��3��L;=<�$@.��B�0� ͟lE�i���!� �{�<#��N+�2�j�Y��m��A�M� ��z���NV�\YȼY����;M`[{�]�������#�:�h��uӦ���?\\�Z�
��Ws?GA��b���O�F� }p+��T���p����ˮ�1��go�r�҃��`�݀� ���M�>g'��vLy&� ���J���b�t}��	r�|
��^1�X�a�uw'BK�C�s�y���ta?��hyۖvm���@$w>�Eb�����Z�͑]�W�t��������Si�M���+U�8�{���9pu660�8G���]�4k��
���(E��@�����r�ۼ �NK�¯v����)6)�������^���v��r6�A�|�q3/��H�OaQ��Y��3K���B�:C]}@���)�\��WJO�$/��`�(*ʄ'X������8�@��0co��`���ŧ�H��BJ����TI��e�`Xy��8��D���H'��|�s.6m4����"ƃ�Z$U�y�J�G��f�dD���π�ǋ?�� ����LZ�������jz3�kCvB�-9�+�P0���&�8��He�{��=f��
-C�Ey������z�R��:v39֖����<hją��D�%!�a�Eq��T_K�or��&��I:���'ऱ8�h�3��?C.K��Py��ϔ���d�������IqH��i������q���R5*.�XW�nC�W�H6����壊���������peBfu��oj�������^�0�3�?�@�µ���Ez&�t�`f��%��\��@mI��WS��BtYژ�.�o��Y��b� ��e]^䥶0�����*)O1I�m.�`�l��~0Уt��Ly�t.�Kd�n�0ӭ���cN縨\������Y�P��Á�Pa @�@:��Z*	�r�.�6M�rHB3)p7�f1�������'���*�ou�"�R�k~�x8c�k�ៃ���hΪOh+"�!)�]!9_����F)t��_�P<>����I�,W���b�#��bS)�+"�wj�n
jH�;9B���_@�^��y�֦VT���]$��(���vx�&��G�'�����栉J�",qt9nL8b��������J-�BvK�q��5^&�=焽��H��Vj#`��?�u�B.��� z���,�9�B�˸��hs��b�ڄ�X��$�����"��W�Gx�?�#�)���98�P$���(E��ދ� �D��DP�ŀx��"z���e,��z8/����PR��$��{���]��6��E�I�"b�:L+��/�a�y�����)�a�%�!D�"�u=�@#X��F�|�$-�wj~ll��޾��*X�P�Ǥ�>hY�hƾbm����U�ZߚI�qȌ<������6H,���V@�Ef%K�CC���z����7Qyӣ�$��=f�Y	u�C^;ǭ�l��q�����p�9Edt�լ�_X�����	á���"�/��Lm+E��7y�K>�k�FMw�e���{�$��X�W���'Iר/ K���O��;\�D���$Y���B�Q�G�{b��4�"t�f��b��V_ܲ����h���&/.�PN�U��m+sq��B���~,z�p��fϬ2���خ����Ǟ`eθm|�d��V��%3[�l�Sl&�YCj��B"��G�m�Cq
���˟$W}|���L��|��/v�)EN��/2�kK�GQ	h��G,z�����E_�s2�T� <6�qtM7j1��Dˉ�2H|�W-oؒc��&��z�ˬ�Be�J�[�vm_�I(�kM�6�'M���tʷ�))���--�*
���FbN1d�� ��ٿ��<n�<Z#\����z�r�� 3c�~�Ja4�+�N��T�(���+sFo.�xCa���.�<��!�9��l�����d���d����+t�9z��KZ%�P
kV�+���/�A�%'�?��t�	�ѿ�} ���z`�U�����������+��
K��;G���B�
ˌ>�O_)��52f��2�w���e |j�nĸ֭K��eˈ�	=Q�0�HU�Z�W�~�GA���<�F���pZ�6�R�B���3��q���t��Aͱ�JF5#��ϐX .�t� ��E4�?MM��)Y0�	�.��k�V��7���o��m*�DbP�#O�������k�fݧյ"_�!��1�� [Ȩ���F6l��$�a;��UZ�E����F��v`�D�ѸE;n;}o��`��̾��u��ג�d�ɼ�agH����k�hP-,��EP��SzoP�iKZrx�NLHg�&\�ff�6/�=\ɒ(����HeUfҫ��7��I�X�W������Ϊ&�	H5���`�Q�gȉh�?9б9�Q�iҥ�ۮ��_�~Aq����[C6� g|�e�Tk�/�љ��? ��2��S�oG��J�q��{�x�~]N:2��{�'Eė�P�b��:-��/n�/q(1���ȟ�420d9e�[akП�x8*��2=钜�W^e�Ԗ+M�q���^�|����%��^x�PNl�JKH�@y�C�w:K�*�����$�t�/Y�M�dA�E�L�'�o^gQzC����˻���@�%���؏��$T�[�����v�Xpӫ�k���5lr�"�L�N#m��'��r�R���ea>q��6�1m��Ŋ'[�%�ԟ
��ff>�3���4��J����V9�噃2Kt�H�-�nm�xd��B�;���^�V�&J�R�uR�,wP� U�w�A,mᓽ<e[��ޗ��2�n6B�1$ �UK�����Ij ��F���de�IN��d;rȥ����=<�T�����X0���z�,][,�m3�~���u(c�(]hG�X~#�����93F�C�Q�~��m��o�R1��>� a�:�����*��]yIP���E*��CB~<͊�ۮ��8���	��*��:ױbúס���fM�+/�`4O2`��Ye9�1b�JG-~�������"��JCQ�dC�G����6;LH������}���:�P����p�͸�<Sp/���[�L'xP���G��QtaI	�BB�3j��@cF�(��=\�A3(�w~� �"~ݡZ��&����X�V��;�7˾)�-�+-<,<�mt[�IH��Ճ|Y0"��5�9��E��'S����A-�+�ۤ}�J]C	NO��/�����1�_Dm����ֶ7���@�Uj|��l����/�b��L���V�,�B��d7�-��.�v��~����ޗ-Ī�{Bo���[~�bN�v��п}+$S�^�E�S���VuX�U�i��r���{o,�oT�����yN���k1U�hB{QRd��AA�,s�Ib�&��wJ7{FkL!h��
��!�]�ц�6����J�����5�8�H��^M�9�H)$�b�>c�=��NB���\,��11A�}����7I������5s�7ܗ���]#��ݘ��mg���|ۃ0�:6���㵍�p"�%}D����$4ఈ��.�뽋J��,PG����Z��H6����1q�4{[Ȇթ�"Ik�Z|gJ<ّ�DVp�|�_��V`�8 �oEd���5���֋%`�/~�l�H�}}2�c�����,��ѿ��WX�mo=S��4�$�Ho�(��P'�`�_��SxȨ��X{�oF���ٸ�^����XU�o2zl�nܥ��K��o3N��|�O��thM�k��h�:�s�������\�f�G�"$IZ���������*����\�_�$u������abK 8��тt���b�M�b��ڭ5Β��Ŧ���j��:H瘖��K%�0@���9	ce���>Ã�֍���p��Hz$�u5��-�:>O%._C��r{t��"�5m���>RH�s��#�Z׃���
u5��(5�C��i�/�A|i~�+B"v�@���|��ˀ��s <0��R��@�8��3�,XuAd�تvZI�5YC���V��yt�35��6d)$o�,��NOI��|"9���o���0F�k8�G����Wv���*J����1���� `�� �A6�57���.����I���ٞ���d!'fk�B�������6]�ˤ��CSŕl��d���l������.�R���r�ŷ��@h�UV�����f��,�.�U��&���@ЕX��y��ۭ�j	B��2�̔��Dz��!Z���6�p=}�����wAD����	�	w���]��(4>H+�Td�%���#��tx�Al�&*V#��� ��.WJ��eQ�a#6�뿐%۩��힁��es9D�k�p��4�~'=="ò�clV�f�*�?���+0�������F��٢�����%���b;:����/���ʱ�sR�F6��+H�C�j�}�CB�..�#�/�������i��ez�(wL�.�s�R(��%��`�5,gՕ%NV~aEF��,h6ܓ�M-+���&�l���A�.E��/|��e_̞M�q����,IG�~[����n뙇�;0g��3\+=I*�}�}}���]��l�W��ԢҠ��ݨ ��sL��_�!����4��׎I���֎���G��D�jcG����gO�:N��n�d<Q�1_����F���������V�����Q��%p��Mʟ/��������t��,C���A8O�����}�R�f�����ʺ��M�X�����a/y�B�S.�_�aZ	�γO�F!N�>�O|��a�q����WA���u�v~�:���K��=�'	
�h4z�?�o����vd��
tNnBS���r�&Ț�n�@���6�л�O�BZ�'8�4��[O�I��ıw�H����ȲȿW�	�:��5� ��Ѥ�����z��'��؟�W۫�+B�����Ap=Y��}�S���6��p��*�̩��Ai�;��CC=���ޚ!�t�zH?p�S2������q˼ v��ֿ˷��Yw��{�L����@�X-QA��$����͍�3$2I;���=�0�-�$7վ��`yK�W<�c��Fȑ���>R�E�;��R�1@�^b:=��̆*T�X����l�r՚��w岨D@")hZsJk%>b�p"��]e5q�n۪<__.��&V�d��My���뉵�;ӊ	��Y�c�����1��Q�yM/ڍ�~[�o�I�O���J��������+O�p�w�|�[r��+����k��"V�Z��zfO��k�ɘ���}v��w�u_��k���ߒ�@�8��tj �A�zNr��A�5sM��ԛ�狐@��F'�}܅����_R�� x�o�\`��,�N0?��S��^�-^x�G.x�+��
�w+�n��/ق�+�{�wΉ��Vx�EC
�I)O�z����	d�79gm�XT�}}�����wo`%�x�G.�������k��C��$�r�I�ok�%��6s��חv��<�19#h�J ��n�Z��G�O�"Y����W"�.i�w���tT��I9�1P�>�(�x�t�F�XR)Q��q����`(}/=�$�ݝ�������]�sZ*_����zt|�
�p<_?4~���^��<�S�%_�Y�x�,f��1+���Cf�#=��t.�?�c������F��r�v�۞~IL���CU:e��o�=��~�.��������}��=���[�9��I�׮�T�4���@���y��n��Nb��o��\0Rs*�>zV�'�?�]7�\��Lfr�ɪGćڗ�`���M�u��ӗP��>��Kߥ"�ap�{H괶����à�v����^�bORn��,��COĒC�S�;b�|z���`�m�`Ne^?���Ũ�rnS�ot{�vLM C�j�薕`��&x��R��x�!}^�8Fw�c�Zyύjc�v_C��� ��z�~�˫�p,	��Q���]�˚Q�/��[� ��w%y�2UtRƃHd��47�B!M�jU�f�j��2���oރʟ�%+����M@ǅ���vH?c݃�o�,�w2E����8b�V���$��w���x,,�m�KJ	�%ݘ8�ڳ��F:F���%�x:�,*^�����%��qՊ�2iԎN�W~��I�Ҋs;T�WPh��[0��<s���0��GJ�@��+��E�b�2c�,:r�,(Z�]�sR)�:')~���*|��w�i�䲖�j$t1��#KU߀�*Sg�d���(�xE9�Vb�8sm�����,�GPS��6�w���'���.l�1I{��lF�"�v�f�OR�í�"�e|ê9�"�Q�Vۄ(����i�-Aiȱ�W���-��?�O_�b7?���[��zໍȏ��j2긑����IF��feQ�|����[^8w�3�/�n�C`|�{9���;����-�����&�V�R����R���`�7X<[� �|�;e�ƃ��P�'�Q�5XTͩ9Nm_@�Sx�_<�N)�.4 3��B�+U�þ���-o.M�h��㿃�d�0�W���le!����z�OQ��̒�+�j��B�@�d�o�uc;�h4ޓQ�ֵݱ��0�J��wk�#�*��.�Ą��i*���*�X�"j��V)sg�a93}L�f���>uqº�=<��2�~�k:B�e�L����zs�j:[B�s�,K�!�����2�Ր"����my�!N�q6�mk�A ь�\ �,���\_
��\\JJ��R����N�����6��$:�Dy��Lŧ�<�e]5Y�Z+C86�_j��4��7�a�-[k����<���6Ӷo#ӽ<<�
e8�'?d�{f��/���qB�A5TX�$�.��˥�칥������w�r�O5���N��f������r\}@�f���*0G�h}��=�Kƭ8TT̑�C?������iƹ��O�>n�{E�]��3Q���}:rOk����c|K�-ٵ����}��")��oU0�ݭ/	xbˆ�*�Ӣ�bg)�(/蛙=#H.�A�2{�h|����-�?�k���D�8�Y^�,���b�k�?�������Œy���7���(J��� J��]��PAB�L��EG���O��ԥ���(|�����o
mE�t-�m a!�y|�3"�Mg�g��k?"=Q�(���K�^�M��f�ν"H�q��L6b�W�{?&E����}���F���T$��P"ڬQ�ٍ��y=�0ܯi�\!�n!(![|.��x͍����&���M�N2/��0��T�G�Y��+#�<�S@s��< l�~]���Ӂ1hb��;W�;[���?��d�|�R& �ʹ�n���=|��jc�����"F�5*���� R��F��}�9W��"ER^XZ�b�h�k'�_%u��
f0��EX7�K���z7BT%$�D~yـ������>�v#w�`V�����5��<a�L]JG�G 5Tvוּ�.�
���O����JKh��/BY�C5��$�l?�������:!����lGm��>6�$@����H���`U׬�+���aP����{צ:gţ���3m$�(����7���� ��"��
}.􍁌l�������=�����dS��Z��d�v၅�&���h��+�$�-��g��.�x��
�^��;��`�1M
�?�n4��/�-d�#�K��l�;��[�� ��Z�Ojo�\V�U`*�>���ݭ�����\����Ė?�C�����N���Щ�[Q�X�Gf��A�R�ϽW:ȍp�v���Kr����U�݃�˻U�ѹ�y��D�/���A�m���-%V�����y�1g���]�2�<�ڎoo��T�(�����՟�dS�\��Q"�mϽ����銞��M�{i�-g���G�yT�K��^#��1} h�W4/uePB��b��s���p�0��oFϑ(�>*�����1�d���0�ӝ��kvQ�L^���`X�~�b��!F��Ɯ�.������a�4�n �%Eek�%K�eYJ�3H�t]V���D�$\��������DJ� ���������o����m!!�0`�&��|�D�ך�ťz�����h3\i?WX̪'Β���cT�R��m�q.�)�'�_�ݞ���� ���Hh��K�kBڅz��ۑ�σ�_���d-|ՍH�o.�{8?_�*�6��\�ͯ�mL(�0�W�"j�+!��d�z`�`IG��,&w��D[Lf;���4�p0�Z"t��^#�=6~�-���`2���a�E���_��yJE��C���kg�ʲ�1O��Ae��/�"��D�"�e�B| R�I-E&�X��D{���'�sF�.�p�ҙ�.��0�;m(��0ʉ=@���&\�)���i���bn�/r��lS��swk�p0��`k��C�ǖ�TB�ʑ���_TU�q��7�o44*^��"��R�TbƢs�BSAU����^��������y!x�a��=���r5�b^�������� ��,(�L�&S���q�F�b��'M3�KH"$��Vk:?�4������6���T�<ڋ@v����d0bŁ�Z�����1~{[�߃��8ՄN!2!� k-�CQr��F`A��	v�c��:~}ˢN-� ��%O��*i�:I�-SSm��_��n[}�Ks��]��.��.jit���ry���c�s9�^�i�4�q��Pz��ѧmoV�!�*�p'#Yʞ�:U���o��i��S��7�:Y��</e10ut����W	��t׼��m�7�W�N���x�:WA��6��7����-�A������*��jf��$�E.E�?�i53<��`sk�+�1C���a��N W��Ă>B�
����ͻ�˜R$��*��/�Y���H���u֟��q놿iN��͏�w4~iT�������Q�L�Vу�Y���ώzt[,�ds]�@$T���w����*t����B7��2��NKg
���c~�UM'};t�����M�Lc���;-o���4���7��
3���$x�!s�P�}x#��o�ّe��'^�L��*|߬�L7��� �A���EFp��M�X������,��A ���Zwju ����?L�v1�'��R�B�2N�+�^q�d���X�G��t�h50���W�\ōL�oH�w�f`!�0hվW�U�QX��j[��I��:��p�����C�S�
���Y$�'�t�q�)�A�E���}~YF���0���ﳐ��U��cS �^���m/n8c5��T?�*G:��?�hR9c,{���~�vT�xC�))'�r۽X@5-��g�?�υ}�V|��56&�i?5���:u�Rc$^�q����eG�>������O�e⥣N��*��i�w�C�i��,{5\3��Y�<n�
Էh�%*XŎ�n�x���ZsS�x�i;]g���NQ�q߽ׯ-�Ma�y��%��e�Ĭ��1�j%-�y>��_�vrO��re�2��Z�앖��`5�^=�
�?������Mn;�tf�՟�$~��Pǘ>}�v��Q4OM�Qz��(�>��Q׷�Œ'X� 4���,F��_ ��[]���G��\	�6�yv���~Ǝj�BF������/]�:Pv��z�18�}��ʠs�?>����V��|�_�_��gxO{����I#,a>!��@�F�{mK%�I�w:&�=km�N�mt��t��7�>*��4�n{�ed��:b��k�`�m��R���A�uŇ����n&Ȋ�/�W�ށ٧qq��fӺLΌ�0�ll����f�W��Z����p�F��eo���0��f�u �[���ؽ�D�6�57��T�rz��4%��S^*mw��/q�䁊dg��@�
��L�Y���8a���3��l��/P蘝�gߢÏ#S}�2xͳ}�*��j9��.�z>D�@@Ҷ�,%�AR�:����7�%S#|I�U\W)����_ef��09Lv�efk�q%`{l� �U��ı����\h�2���B��q���m=^QlH�L[Z8�9�lGGM@��V��\e�@M��x&J�_�;]���kwt\GS=ջL�؎Z��#RÛ�iX`���3c���O6=�Q��u�5a6$�(�)b9kD�����S��m����ƀA7���!� ��� �DG�|��a���o��"�NZ���#3{;���#��vB���o?s��9h�4!m�悯�	=�ݣ<���:,3V��h��^��:���Ə[���<(��lR���]�͌r���@�a��6��8�U�J��&���+�-�ABE���P=b(6�u�@1MB�o�䓶2�0����-^+u׿�xf��h�Ӛ�jؽ�R�� u�p*�Cpy��ПK�IC�ED�OO�B������R��	��0 B�7�AA��	Yp�&� �,T�U����y�]�bTd�}B�� �2� w"��dE����lSIɲ��6�<�aRX	!�I�mM�'��q�S�+߰������c�Լ
NS-��J)�4�$�z��1���׋<§�����_3Zv{g�{7�~H-�a/�v���S�Tb0Sd��{ Z���:2��/Q�C�DJ�V1�}�2?9`���zj��>)�o�U����v.��#Ò��C~���g�|�F� �����*w�_!��]�b��x�P��h�P��.\I�CՐz���^~�`��*���:���_�,�a@�c4�3���o�<t�/�&A�b�߅B�g�?�4�pg�{[��<:0;�#�P˒��UV�"����r���ӬK���~M��:�f�+��D�B��s<�^��PH\��u���� �������4��t��g����L�$S5��	�v֒��Z��,�:tY�}�ԧ�И�BE���b��1\娙X��1�AA��r�L�]-���C�(�1qJ�R��}/3cz���.}�]��S��8��Cl����9π_UbՏ���e᥃�S�\M|������9����y�?��Y�ƣ�� ��kje��M����&����,j5����{���^W����D����-ݝ!���yq���}ջ�V�r���s��3��Z0ht��\�4��F8�\AQ�҂��>d����lgyN1��w�t) ���������E|��6Ӵ-lX!�����	0�!���ܳ�`���x�3,="`3�b��3��f�
��H>���E�����&���,�H�*b��~�H�Vp�)i)�ڻ]z
���G�3�Z�|U�vN�拘:��.}}��[�f���ǵ��֩�E��S�dT�åX�Ӛ�r�WJ����:�A��L���I=����5~b�v��@���v$}DJ�m郎�%��~'������3�R�Z�bnrb ��o��'��sI4�<���-�'��9�t?����;G�F��t	���j����~ �#������b���y]e�1܎f�U�]E>/05q���`M�A�P?����x���c<ٖk�}��Y�G�V$�#�~�0���
�SzMX��)\�?�^��{�x>L�e���<*dk�_x���%�W'v�~ipLi���Z˔	�O-�3�.J���Ft���GI)�z�r^�˓3ʭQ{Hz��^7鐊3k�3�G��̬$�;?ǆ���Sj�	�*����TFG��d�=�]m�A�b����.T��un�}�[	)�Y	p�˫��ԭ9�����5n���f�b�8��[��v9����P��J���y�u��7#�MM�z����lG�K帇�����wh[��'��q�1s�>n�и+��z�M��m׸Tӓgb�}6
�HEg������V��IE�mY�}�����#���e�W�Q'��v���y�гX���b.;�Fa������|�@� �4�ݦz'������b���i�LWi�	!h�*FFv�ͷf��6Z����]x;�.��Oj9�E�Oɉ�a
<�}h�����'�x*�]oN�И�9/�Ov�HR/#����G+5;�\��D��vy+w�U�\���p�gt�%�-�UK�Яn?y9��5�!s�&~;i�[��X%�=�1�a} 7���+G3��d��U�ʑ���۩�L�D%��tr�Ό�
;~3����F�	�m/��v�&�"����G,�GƺQ���A`l���*�S��Ѹ^�!˧�̍�d��F��	�{#��ծDR��<���l����Qk,o���	̹���E�zb
�3��ب�T=�f�o%ͮ��U����~<�@�|4��E�����@�����?�/�^�-�,2\�5}�#��u����P�b���%��x����9�W!��m=w��l�^xl�����s�'���]D`I��;N��l$��~�?<Ʒ��'	_��Ȝ�v-�T�vv�r�����1D
�� �� �I��ǳ��3G%��M{=�_D���O�i��sk)��I�Ssm\V��#�P�������Ԫ������ܿ )x�܉�f�z
���?"�|��1kã��~�>�z��;k�^�2��ĥ�l�]^��� 4�il3O����f�$QΓ8V5����\��S�#��\	�t�~��?)�);{1[/���ZlyA����\1�; d����u�7k4zY)C��t�X�Eij�7����I���Ȱ�hq�z��G���$#�OAA[�!n����U~�.�&�di.{z���ccÜ�O5(R���뵀S[���1�|�@?9�W�@!IR�c�j��
�T �~\���������Z5�J�wgSJ���~�t���dF��M31�v��^�B2�(S�S`���|���u�u��'='�.�J���!Fϱ�'���N�4�b�L���+2<8gɌ���K�t )�����?�C��>J$�Ϩ�K��R�썖
��ׂ���n�a���iQ'6����5'趼9��L[$�9�nYyV����ᘷj���E����*���|m�kc��\1N���`�g���ٮpa�NN�h7h�SɱG Uo*�Ǔ��#�}�񒴝!��2��1�5ɰ���9c�맘w�W�z�}
�k�'z{Y;�p9�ve>G%��:��vi��粵&k*�VR`b)$Y.����\��ϯ�o�˹��Y?���wl�����`����Ee4*�!2<��d��ƿro+3QG�~�&\U�v\/����&�1�2OF�vQbZޮ+מ���l��д��&m�CznuP&4+v���c�i�L ��ǖ�8ܓ�������y�	p�6	A���ABj4Af��J�����Iݠ,����$��Qn<��ٯ��gEQ�z�������v4z��VY!E�Nߤ0ַ�8�� { ���A�#�ڿ��}<l2�:�Ui�NڙO���Լ��n�T������z8 �'BָQ���\X?u$�Ѷ��Z]Q�$/<��ځ�����K��\ޡ���?z�7y�G�+�k���Y6�#G��E����(�d1WM���8pZ�ʺ��[�8�Mܦ�����!�kg�V�MY�-�f�� ���y�ltǴv9�?N��  T�v`0p��L��~�	%
:tv$?�T"'e2b�Vo�؎^u�aC^K���ֈ�ݿ����]:��ü&E]����X�TU��6/�ٴvkN�_��s��ɾ��\�@��whF�㣰)k�)�h��-�!#��z_x��FG�JC
b2�	ؒL��h>P�	��v�ҍl#�*��(ؘ�	�eM&�t���z�C������z���F4��Y� �|-`#����ک��*!ݹ_�fw��C3�7O��6�:��ڷJ��f")t��V3�]V�h�6:�P��V''�k�0����L�(V��|�[A��&9G�<��K�h�ȍ�/4��}�
e%�\�ň��K�Ň��T���c�a�Z�Hwu9?�T��Q�}n��h��/m ��hb�V6	�J���k!q�M7��f�N�\�5�Q�(�����G��:�e�z���˷�������#@�/��3��D�Z�8f�5�K��:�.�8k��BZ��`Ѭ��_���."�]�����)&�6���R�Hk�����-��2u}A�9������P��
p�S=CU��8����]C|�u���,����~�1=ؘA���"G��#4c�B),��Q쪚l�}ȩ���13�P7Ԉ���	������`�bl�=�8����zj�U��Ʀ�Ĳ�6Я���iүb�Q<4\`�G�?pI֚Jρиd��+P�r��rtߡ����o���s�����Q����upPrf�C9�E��WT�_0����XwU�Z�~7>�@���J����'�����>�~W�97L�;�k���- �0s�.���ڞ+i�5&�Fہd�n==�!(��V ��,��~��	�_�>N�Iq������s'	
��8���P��`j�B��D5�Hf���|�KX���l��p��79J�7c�B���3�r�J�^~��"{ղ�6�������a�*���V<2lE��-M�JG��5˝]�tfq�"5����zJ[g�q�%u��)Ʋ�[�Uj�B:=.��ͱ�?��$�<��p�v��f����GO�3��pa�X#����ٝ�[��ph�F�ҵ��c�>�T�&	����r���n@��W�����Ъ�����ėT8!�F~��'ئH�M�_h�t��&I{c���n�K�br)�O����ko�3�N��_��}�����G�!���{����l<�Fz��h��%�����'�w�%�L��X)baԎ3Xr1~Y�P8��9�k�le��f�ph;�T]=0�4��3���ȑ7#�7�<������O���EsANx��[}�-z�k�U;�|��!�{l�f��d�πm�6[����ڹh��΀c����r�1�z/���o��̇�*�@J^נ�+�T
	c�]�7g
v\�~��aq%^�9��'����!��SM�i�
�OC�1����h�����l�?:C���*	���VYmq��̢�}�1���i��(L�t��11�=��{��<����Zi��3���xBz�z��C�	���Ԙ�b}i��/댏�	��e�W��e�uO:x;�9r<'��K���T�2>(�F W�>�m-���R�$���E�_��˩-����rM��Lh�)Vy�+�ד]�"M�,�%���f"	�����\�{��&��Z�o�=T3E����b]yt��T���[��{=��\{l���K-iN�K� "6���[D�*��|����R�&$���F���|0Z7��)Ľ��V��}�&�}�2X�0�4$y��Ӂʩl��c!�#��Z^�l*=����Rj,��
�hᮇ�	� �����_;��]h31�8��R�}&��K�d���['x��GUF.K�.��wM�TZSmyw�"d�Ay��'�%��c5�G(�#�}��r�?�n��e�]$k+�<�P�ħw�U�?\�CT�_���� �̉����و�������	ύP��E%"0����Vh!�n��+���~�C�l���K���`��~>���ũ'��c��W�0z�l.�ڡP�a��v��[�,��y�X��,�,�r� ���)�d&��Z����+G�?�ݯ�q,1g�#���/Zf�Z���q��C���+�,7��W�*Z���O���*�6@��S�����ӦCˆ��D����4q"����m�F`t֡�U��W��ubL6-��	x?4�� \U���ڧ��}kC�_�9�@g�L�MD+8۶��7�8��I�� ��>bH[/8
<X��?�J�,����dI�>���Ꮎ���QA,��	��
T瑍���ѰS�8=tJX�#�)��K���@r�m�$	�J*-��(<J��IyP�1 ������B�P�kߨ�tI�נ� ����� �cu[��C(!cdwqo��1^�# ;ͫw�eu5���t��U�_g۔��J�٭`�|�d�)�3h�	��fN@��'w!�a"J=:��ޡi���@w:�P���Xk��=�2�N팶J~�D=6n�>�a�y�}B�3������_�):5�V!�<���}��V�1�G�����	%
��I<d$�H���_Lk���i�q�v��4�s�Lq���FBvsF�_�g�q���lH-��sU��(ʺ ~�\Q\Y-f���՛	FZ�#G��+]^�.�A�x�7��s;�#�;�[O� �����<5����$~��nT[�BN���:_)�k���3S�z��G6;mx���C�Y󜍏��̰|B(EJ����L�x��Ǧb���ClV�#g����7����T�ŏ�Q��0�x2"L�.�Ma-�cd?R�7��E�dH؜4�(ò�L�L�x��(�)К����'��h�kG	��@�P��:�����ڡٗX��{�,�-=b���݁ ��T���+t�϶��Ey
��?����f{�	X#�po&\�_��۰��0�ɒ��6 ��JK8�t�eH����
i�*���YJ�:�n�GO罬��d��ҫ5��pDq�9֨�J��R������������G	���戤��N��k��L�}�tY��|!��s�3ጢj���Pߟ��!���迩\Lɪ��qB��獵
:��=��ez����n͇.R��7r�ˉ1?������SZN�Z�t���ݵ�K��'s5��0x�j^n�W�h�UP|�?��ڔ�s����!,X^���k�5� \�J_��\ޞ(+vȱ�.� ��(��'KG���f�8�SX��ਗ਼�ُ}��e���K���aE�}4K���'�,ځ��Sh�jU8Nc�A��zlb#������n�r@��Z8�C�Lv�*o��
���j�5����
j����p.Չm��ܚ��e4�[�D�=�x�	wp�zz�&��d�g� ��v1U���z)���]R�HSN��GH�EJ� �E6P}�h�"��2���]���e
q�P���Y����"D4JUD�]��N��4Y�=m,T�G~|+�|b���Z��	*�5ЗW��.8@ƶ��r O%�is��`j��@���^E\SCC%���@${0��7;��x)�ޣ'/h�7 n��>K��,d�
pfj�ť<���C��xJ��n�{r)ԯ�j��WS� hԮp�4�:j��۲�8R�c�yE�{D;���bQ�죕�w� >a�?��7Y�Pv�	�I�����mkP*`��e�b���}}h��"8X��)'��eX&O���Kb�q�QZq��jp�2�ќ���C����%4�ra��@cCQÿ��0�>�OJ,����o�@�����T���<��%w�Ȓ�zk��i|Z���0`��P��	[vX:���ǹ":�vۗ#��η��Ї����y.p�5y_]�ZgC%S7�c�%*��Պh⡞�&	�r6/[2�.�N�x��kpmI
8Z���kT�{���4o.\sQ72�		W�NO�����+�ں��iP{wfO�3�f	~[��ܑK�>`�^4�*%�*�|�
�x-�wo��LZ�wl/�u��z��7�,ϯ?��=�?���ڜ96���1ݍ�'!�����c�������;�UM?,@ޒի�����w�5Ō�BY�4S���|h���د��y��)�[x@�.~�vb��~Ё�&�"�E�Å��rdK���R�~X]�����Db��t#ċ短��T�X���Zک8��3���/��D��q�q�E��綢� 8�a�.#~q0NT���+v3M	,�j�� I/wj�ތ�k!;�ϻ�SĖ���䴵b�C�ߣ���Ƶ#۬�/��s�yW��=��џ�n4�0�Jr�,�'Bߏ �$Ϛz���q(%�E��x���0�5����q;� �.�+������ j&�	��R����v�62,N�����K)dw�u9��G/t�����OP�C�0��x�����Yh���~�S/7�_��D�`1�;�jz|��y����ܥ��S��%b��GP�穪R�r�����`'vs.����Z�����Tg[���@�0g3R���D�#�6�j��Sm���>l"�f����gάm]�I�cjS��Yk�������{k�֡=��2��R�}lR�46��c_.�K^��#��>'��Ė,m���j��V�l=�6����U踉j`70z�Y�]��*��r�3z`B�W�k�i��Pq[3X�b�I���G��m�!�'���e5RJĻpn<�}ᔌ�A�>Cd0u,vԕB���QVk-��o�(�b
:��y���Z5`c���n�]�|�SEl���N�6<��,@L����>�	
E�s8^���qw���[��Nn�\#�'�4�r1��4=M�5����:���HDmm!��${77hg��̛�4�el� �?��;��0��y�u��V���i�$l�f�;n�^itHS.�g2�j�T��NSp׹�͂�\��U����p*;8%x��M�Pzs�t��C��&/N�)��y����SD['�}��X�t��"���贯:�,����kx�,?�VOi��y!B4��\i�4}�Υ�Gm�+���c0� ��k��J�sw���A�&m"cGX���w�3z���[�xQ����hb���D�'����g���͸>70Ï(k�B��x���جO��|yP����i�&,rM����1y\�����R7\�H�':EY�/�'�� �d}���s��L9�k��z��0�OC������~QuqQ��+�xހ����Kí�}X�bv��U�ƪ��E�b�9M� �J
+�J��h�[��e��ջN=��X�1�gw2�OX�m��*�dE��Y%Z]\����uLO�n�@�*R��@���3l���I����?�m�L]��rE5�V�8a�2d�NB�A�&��ڛ.���KC݂�5������o,�	0{r`�D�N�z )�^Et���2�4��FLA��%�##�,�mz6-�#C������u�\���AfpƖ��ʆ�� 3~5�e�,��|6�q%��x���ǰ�_r0��-/���6�z<�f�.@yt�շ���i�'�\*�v�X����j�����!�91����Q<��`|:��C�Xd�h���]�A��M>r�����\��t%��7
�����C�	�𛴴��?�N)U2ϛ��JKΪ&�$]�Kq����qs�0�1�>��N��j�Y�����4�L?5��i�2�'@�fQ5�n�-m�f:B�^���T�T� �C3tE��0w.��b脄�;�S#��]\�"k��\f}��`k�;���ˁ�As\&�e��ݻ;7Ix��뎍���̱�g)�x{p��Xuy�>]�A6,{Z��#��ݍg�,��
�Q�.�j�vN��`5�����]#�8���b�oc��C@�P����)�
rt�-��v�znIԠ=����Q5�R�$Ji��	Fx�s���8��@���/2bd�9�!k�
xc"V�J" s��CP��������q(Sm�{�b�j��5媅�jy��H��ͲN{���7�����$�Kg��3Ǵ{0�"u�ݷ�y��W��*�a�LU�P����9���ƾv�
]�r]�hp�<{7Kp�,�v�X���[zY�?�|f�'*��5������F{�n��e����xL��)jSLi�\��K�f�!�2�����#�b��Y�N���|�r+ ���"=J��sy%"��R��V^&�E�b>%g��"mC��/ժ{���(�(VrB媒� �j�yYan%�k��}t��%_��.�feRz�ъ`�S��T.G[$�C4&1q���bA���Jp�\�ɶ�Ȍ�WaT%�wtC�	�64��Z!�[���$y�|�����Fp]I�#}qi���8 ���gة`�7���Y�ݞ2��R�� J\(pQ%�� !�i/����j�3��cʘ��q\�=�#Fe��F�[�p����$���F/v��p��7�J�Z�eL ��%�k��)�Q�R��5_5k��+hV��l�7�"�)�_W[�3`�ix3�YGn��������1���|D<� {vO��NVה��|��x��5I�>��SCE����g:���F�Ў�����t<-�؍&�&sRMB<|K�;.�F+��3-�����&+�����/����ha�;~u��!�Fv��8�7C
�H8�0�:&���]�o�K�Y���ѓD��@cP��=��,ʤVp�K��	��ߟ�q>�����z�Է�=l?v�U��B0�~ ܎KOI��)��#h90y==p4��>9 �ܵ�b���33����gi&�+�j'����6�`��q���4g����^S��q���D�2�gƖ�O-�]��wb�8�g�w���! )��5Qgl���|?�"R}�����R��h��e���$���.��S��ZkhSj�,?�G�b{s�G�,�ځ�Һ��iνU�yC�ik�i=7�tx	�s����YK����!zT��� ���h8�&���3cq�ݪ��x~әu�$^\7�{�<�	��8�"����D�J��/{��&�趍AV7g�7��9��-R�b��E
��1�YC�?[��L5�\�2�����bJ���Q��s���!NJ��������Z�B�-���bݿ?aL�k<�)u�:{�-+Qbm��p��&�:ĐRXX�	}Z?���
�YVK�6L�l�&pA|�Y}n߄W�z�3@��\��m�?�)ҿ�C�g�����4��Ao�FԽ�Wȝ�#���ڲEs4�+�S����b��d�x]*�omϩ��-����v6�M}ȔDK����rf���^���2�@���/�X�/m�c��(�ٵi�5������9��z��$}�$z��O��� ���6y��
�=@_[$k^i�7*|��i�� S�
,��g�e��2�qmVЃ,Oc5�C��'Y��<�*e=	9!r]���
�vܺ�Η��c��R�Pd+�{b� ~��`/��]�~O��<�c��<�Yr�)�Xs�Z�$���@Oo�랪}&bt|>�"<@`��U��볜/t�J���}�OZ����H�Ya3ǖ�Hb4j��o�i��,_X�n@�X�{��/|:-\��M�,!����k�:���XD�t+���`���ױ�;Uչ�����(�3��ޠ�4E%�OC�E�q��TNM�y���Ȍo�Ak���B�!/L^Ά�➞~C��ȸ�~��Y����6U\��������X����%��B[d@`���p���h�<8'F�Ud������)�_�W�[�7���+D\xu���(�Ú!w�U�Ε_׬��:��D�ZTx�z�N53�.j�������/2���f�������}i��������əK1�w�y����ff �-�a�R��2IZ�Q	).T�	�s�j�k-~W<�ƉG�!�섗��S7�.u�h���K�t�J� �ܷ��Ī"�I��D]d��HU��b��{�Ϧc��� � ���]>b�	�
8�I�1�������zPL�E�]�ţ�6! �)�7G�hҴk턐-%Gd�O�4W��6ֈ�����uʦ7sv;���N�\m��@��V$��ΙL��k��C]��"�����k�m��4꒥kr��GnX�(*��'��{��_�n^��e��J`�����^t壧չA[���I�
ua��؆:���+���Î�� *������d�A��,0��1��q�6���M�LR�F���?>�V�|�}����[��F��������˒y�B�F����3T�܏�{l�j\�m�X	������3���f��e2S�B�4��p��<0�п��ة)*]�=w��zjhX%�r���,�[��xr��Wo���"����;���7�z����{�����A���7���w|=�nR��z�����s��)��M��0y�5�������>���L�:S��6�$ALr{��D�+K��$�ӹ�{�a�?:�0��til�"2�v� �Iؒ��{@&���|�1σ;!�>M����u�HE���h&�H�t����C� Uqk �?.`��E8ҪDA(���)I#��-U	XW�ho���� 촗�$�쩋�sv�����~|�n�,��[�j�2֪��B�;���&,F诖���;�i�q�Eլ\�af����R�I�_�l�D±'��� �'r�A�|�携���QLf��L}���n�9n�{�z̓����tB�`*zzwÿx9�f݉���x��m�R�ؖ� w�g)m�$���t)�A�fD��0F�H�;)��M��4��U�Ϡ��m�.�F$N���3��������l@�d�^��Q�<��TQ.��4�^���?X�
tz{�k,��^Eɒ�N�v�M��>7R�/utDHu(=�R��\������{ԓ3d�D*����$^V���7�|Z��uk���:�p����!$-���+Y�︟�[Ԥ� �y�m�0����z8
7��5P��b1��ԟ�n|ߨ���שa���3��I(����F��Ү1��'��_�`vʛt�A���ifm;e��s�1�0���O���l9�PY �����NÊ�o���ͮU�^����"�&
�`&��j��*7�K_�h���ZF&!�J̮���b(���x!�_�8�!���R�V�'����(����(t?�E}k
�7�6�V߆Z�3I��x}�[}���<�x�XR�u��&���؇���}L���y�/L�
�M'�r����D�� �K��L�xe��T��'�@$kLʝ1p��Ǘ-v3�9�b���!g��-�&�[�u�W��`,pzx�x����8*|�/�^��T�m�}�OT~'�*bK�>����p���f���
V��Lش����;�N`Kؖ!/dg�k�����y�#���ig�}�/߫#�jT�k��.��1��/҃9����M~ur
4;���3)h�ѵҵ�&)��}�pq�.{�,;�
%�[�ӄ�VS�����r�]��(q��/,y�d����sZ��.TU���M�Bo��Y�[e.!���!g�>��N�����6�V�?�q��g�r��w��]�_�b5�$l�t�gi~�8Q^:���R��<FC�h�oy���g���4(�k��-���Ty|/̇H� ���9x�|�c*您�׋�����܍d�x��d��=�z�kƒ��^��=0Ǵ��C���L�d�cס�����S�'W�\ޡ�^V�0���g���,0�]�C������C�5��pF,QM	�'�xZ8����	��)�G������[bg�j�G�z#Ӫ����@C�Mǧ׉F��*� ��~�\+)U��]�Z���8ۈ]^�������k�l�[װAj��[��j�	~אxhZ�*J���6)�m�o�%��I�!��w��W�qR���w!�����gl+�Lv|[�z&I/�F�nηg���*�����Z��_�̓�!.$�&ό�C#J��co��!�~��ʄ���}�f1��m��I�Y'G^[�i&�pȘ%X�:Z�~��)�tn97`�Ĕs�[�Y�_�V��;�3��Y��T���t�V8���q?�Q@P�n�,5���+/���-ᘋ�!��O5��,��#��T�����Q]؂�I�%�t�/Nk:��E؆��:22��c5�c��xCy�o�(��$v(���$&�?|�GO3��zyy�a2�-K��_�Z5&�bƘP)����8V�D��Ԑ:o�68ݺݙʜ܀�����o���m���+�e򱍥6>%�RŰ�f~�N��H��>M��ڪ`Fɯ�} �ݧ����ʵ���\�6�3q��X��)������=�꼹�0�dP$���o��e�(GP��2xm����D���\����ըC�p9���(*G�[��$x�Ux@s�V^���&��?F4�eײ�����=�.���VG�B4�6�~ol�ޫ�f?�Rr9L��u��q�ܬ#4!'*�@6"\yv@#����x�5��@p�̸�1�o)66��#ʬ��W{�V�Hy�a^����v
�+7���ݹ`�w7�@�6��b�@���8�9?MEr��w�}1��6�XH5���L����L��9�R��C7P��k=�6T��ʪ�yB�V�*�+Y��ʥ=%cw^�fE��P�Z���	fR�Ѭ�����Q�P�P�3���Ү��sb�n��CZ]P�8�^���*�	��)��e��\cz�D��_}���J������s���'l�*p���Je���_�t�p�P3�G��YEm�1Xr��p"p��z�1�1�#cB�Q��=|&��4�^u�@�6�1O��	o��Ti��]d�������q[d^���ɟ 2���(�ת̛���{��ϮX��?2($�N���վ�~���%`�ZV\�G��ׯ)�d|�Ig�����u��	��NG'c���Lg�#<�(m�@9��ae�O�T�ɉΈ,0����j� ;8!�c|��XU�a�2�d@�~�j1��s�Cc�?[��t��u2C��z�>���9a�=�[C��a���GBbS� ��N0���#ᕕ
���I/��Po�)g<ޭ�b<u��7ȣ����(�X�~!���.^jT>9�4�H��H^�#��@�	��;?�/��tL9gͲ�P�,~�|���3�~ҥ�CX��SL��&�z>�O���~�r=S��S����,��ƭ!1���\̌��D=�<���*��nb��l�����ʖ�>|�-uz��{�C;jpJ�l�T�X�fa;;X�B8�>#�$M��ϛj7�>�M�C��s��7x50l�j��u��O�3�@���� gŹ~���B	��c�]�}ݪ�����F��6 5�9.
���BR�񐙃���E�D�wo?����ֿ�]D��	�m]��S�X�ñ	��UK�X��?lWr��q�EA�t	�=���$�}Y���(�p�\��a����&϶b;�u�YM�'��P/�zx���zi�اF$�S� k�+�fw��f�T�j`�S�R���it7/�3�]|)�5��n�yg�����J�^�u�H=K���[���-�>n���w��s_M�����ʨ����O�}�����"4h��0e�����G#�����b���뷾~��)3;�}�?�K�d��ػ�{��B�[�T��֔��T
������oqa�_�8ec�� aY�Y��e���t��K��ܵ�e� L.�z���.8k̙ݹ-��ʲ�*��B���E�.�J�������M\x&�(C=
B�G���5_'KCW�'>��y�fи�N��!MR��<��_�k�V�i!3͆�7܍�Bn�z�;��"�8|
4�x뼱@A���}��3�W�X��T/+fSX.CP5�=��+mۦsJ6��スP���i���S]�.�;����eF�e^�N��_�G�'�C+�J>G�Ɋ;�
VF�xX�nO�� H�����M�w��� ��"O>�E1���L�N�_wCe�	M�Oq��K�A6��s��~��5��A ��cf�.�a�j;|A���;�5�0�r�,=��e��V��(�� G��Ad���z�44��`�j�{��X��|t4�鿚�.<�-��[�=��w1sÜ�$��p���D4��p�'M�9!h��-�nc��,C�l7$�L���)�h�3��2�n#���O98��5k����hH�2`zZC1Z!õ 3o�j"�lh���J�V��%��9��"u*t�F�X)�*q�/?��4	D�6pĖ����rkavv}+�1m.R1���0�P�_Ӑ!��]*v�S=9���u�]�@Y8�����8�U��8�Ԙ�b�%p��#���D��BыO[��ך4��+�>.�:%A��3e߼��8�����i�L�z�Kq1���m�$ה�n��Q$��"xI�؝w��@�(T���ܾ�%�h1�]��B����>��i������ �:�
�TT}���s���C���8�-�\8t�õ�WBo���҄K<i{f\��1��36d40�ݼ�NM$ƹT����aۄ	�A���!�_hФ߉^�x��;�ՇS2]���Pߕ�1=v����񄍷�(X�"��wt�}a�p�4��}�ʐ�}���GVܓ�Ty����I��V{i�$��		��i?���K,A�'�/%AS�Ή%�p��AA
�s=�TA��^5.㼚�mY��R�h3dl���gt6�'R6FE�F��t+l�����u���(��[{b`�/	�֨`�kGpj�����c7��Õ���X�b�Y�!�$�>^��ϕ7���L~��	3�\$(V�\��\��c<%���vl��Dm
���ӭ(D<���O�Pĉ�����d&)x�����z��|L�Bk�� ��kɢ�p^�Q:+�h|[v*��{E��;Ͻ�$ ���4A�"�&�t��sd�*e��7����sL:1Hs���:a-�ۍӄ�p��g�m4Bo��B�X)`@����Qz|O)��]�&z��Ċ�aˁ̰̟�x�G�]��ð���M�;���C�Zh%����<|����29>�����;4;'�������O���ӣ{���BP>ӗ��΋�럾ȕ��T��d�Ĩ2��lF��O膎ˏw��^qG7�����ָ��,bҴ���4��O9��YSh6�ݾ�\�k�r�ES4}^����ѭ)f7:������ɔa��=}���-��8ѻ�ҕ�G���W��M 뾗)`,��˅�wFn)G�h$鵒���b�b<����� v\t�L\8�!��~KFr�_~�!Y���BJ��+�Zh�;cJ!�<)$%�gSBޒx�Kf�7��I�`J�ra���N^k�N⺙~ez��VWaO(�k@kj�ڜa��C>���%��r�C�lL�K#��U�f���� 2�0��*;մ�Ju�mP���F��Aۋk|�h��a�2�����WZ(��6��Ɨ������\U�u�d2��זbKe��A����Ğ���w?2�BT�z�[��"�^�˱b�:7Oޮ'X[��[׆"ŧ�M!ZDL�f	�z�w��д���)D��L��N�qn��%�n�;GM�4];�3��v��O�%E���T�dN�%#���Ǡ'o�%�j���=Q�@3J��)�]���ƥ�{u�d���Z���";����?RV���.nL�0�Ph�j���P<	�{��'M7ѹ�{���������q�!}|s8ۮ/l�fO�����n�E$B����j��p�Ɂ5�5�
�MR��L���-�]i��\P<��H�G���)��R��w��l�R�P����JO4x]��v]l��w���QF�ƜD�grF���!W)c�c-�7����r��K��Q<��	��F��ʫjk9���}�%�m|���u�y�}�e��b��N�΢u�=��ӃP�������˾������?��">�ˋ�=Pɮ�Ӎ��Èhk,<�(��g�<��M�g�q��E)C#J>jC^�^~��ݺ�Z�H����	q��'��z2��������ɖ�렁�[�I��hi&\�5��o9���G�uddQ9«��t)�^�i�4�W�Ay��@�{�1�o��B�|�u�ض偘�r}�gw�ӎEk����8�Ӽ �Վ?��ٰ;D��V<�X�HN@f��,>�ʧ)��������|��|��u����n!":�dK5�DΤ�^��L^8��#�ģ�������X6&l�
��|R	h��L���Ӷ�/�Ҟ޲��-8�I�{F���CSm���6�g�T{�> ��p���7V9ڟ�:UoA��_��{��d2��h�` G�_Wy���Z��w��>!L������_��}m��3�`��7*\��^v��V�J�=�nu���g=f�L.vX�ߟ�_����n��?�A��_!��ɈP9iMJɟ{~&�C�#�7K{���R�H0m!C��j��<�̌wVl� �;�29RrsUіo�N�0���j43V��_{�r�v�xz!���YJ�*�C`���}�7`(+?�Q"��N��W� ߳�~.v9�=W��kUDh���J��`"#�N7�f�y"�l��m~�<�yn6��6Y�׊G.�r�_;i?���o���_�`��Sw�%ʉ�jW�-�M�<���Lc�&��n���u��C^a�*ka�ҫR��i�5 8W$�����L.bLt���cG&��iI6�����~f�:D��,�5��g7���L$�<n0Ϧ)o�-���[28�!�e�#�	����ɇ�nl��O����\�F���Ao\R�0Y�e��(X��WF�F�e��4�ǱTQ�BE{�%���K�Y������QZd��꨼/� ��{�A�]�%��/sv�	jvaA��4���x�E��b�L�-QX�F	��K�����~�,�b���._�2m�5س��(�e�os���iZ/�i�zl���[̚���++��m] �䏗m��}6Z�&V�M0 {��?��4����T9�o�s��"c�߿�n�'Y��I�D���s��Z�3	�5r�a��/(��b��� �E�$E���٠�D��QZ��(�s��C�r�Qbr4�t�Ǒ�^I�AR����*��D�1E��|���;Y���
��
5HԴZ!�-��X�X,�Ċi��9���C,��e{C�K�3z�$��|���7%NhQ�Õ;T�s�O���˥FX,
@=�|C�_�!b��>8W�$)��,P+xnn \���6�IӴ�d4ԙ;i}P�>�EJUq�_�ƿ��Ur0
ы��C$Y4�k���}�����pTF)�,NJ+���K)�yb�N��9��g���qW��=>u�R�<x�_k�Ҽ͂ˇp��7��6Ń��"4�Y���$�tO��]3�զ�H�!�8A5�����W���ȹPwaN�����ƙ����r@��W^��Ѱ�'�Cv��5�wE��Ԯ�T��"�e<�uB�����u]�>�D�T�$=�(ꏠ�iE�`o��'��޸/������Vv0�=�6��&-3�B��@,|�,�ʠcizr�KvU�z��|��)�G�1�/E6
j��"�a�p��Y��O9�
U�T�b3�x�����Wt�ru��%��,���w��b�O@����)��gҊ�+�9���]ζ�S��ف�k�Q-�n5A����l��1򮛘�yCA9�BDZ�ҹ��|���������VR���z5���f��� ���x������U�2�5Z0��#&hh� &\f:��Mcf_R\4)O���^�Z*����=����H����A�ំ������a�"1шo�zZ��z�i,`�e-���`��~%ʫs@=�{MDy;ff�`W� +s\�#�����d����a�~�B�튱}�n��ҫ%k˦7��ܣ7ҜVGȮN0�`�бK }e-	���Ү������6�0�j�^�Z�51)��{?M��#e~��ǉ{>%��lx\^���{c�{��A��r��i��� i%�������r��@8�z7s��!4$�%,��av[�,(R�3��M2�I�7�J�!Ei�JϘ�bC=�&!%"}Y�(�)�VE��B�(!<�=+�9t� '���\���G��cE���v�$���I�ڶ:U��Uj����T�e�V����(�!�z�UoMX4>���r�X��M�Ƴ-,5�K�o\Y�6��{Di�^���g���h	�զ�������Kʍ[�v|��j[c����r��z\��"h�G���eZ劮�'F4�W?�6����"������q��+������
�G������ui�!M��3	�:3�G�~�l;�p��j����T
H	Bn�"�h+%�:V�\�H��Pu?^�_z|*��O23�L�j�����iNO�1鏒d���.ÒoE���1'A��Vy�(lͪ�#VD?�)�wڕΎ@#K4L{ �/ꤜ�F�Q=��Cg6vS�ð<j��� ��%jkK���w�9�By�l��>=�[j��Հ��#��ʿz4���MH&�K�%AD���~�䕌-�N��@dr+al3����F��U���0�";/���ץ�ݥ%H���P�P��orI$D�k����"Ѐ;��%��v%C��ٮ�>�UӘ!��&�I@U:߫%����k2'<�9�N��`;��{��a!X��zV��d����b;�)�5���.�fa?W������L5-�')�sQ�Z�XX9K�҂@�XJ!�!V�`�͏�bJ��4�?�~ݷ|�,�.�d����o8�n5�{)oN��q��V�V�o���+�ODז9g�҂���]��q��ptLo�Ո_�:JS�Xs���\�Z;l9)��\��Pu�1��+�ϩ"���Ε���Ꟈ�Q��!�lA��5�`��(�����	�Xs�GʱU�w��Sk�U_Ӽ����#�X ��x��"�Ln�sR�KyhVYV�u2�.ikﻏ�>��UHby����<�v�ڥ�}�ʳk�&U���7q*<�K�Wc�C�V(/�K4 ^�#��Ҁ�4���$T���yJi�Z�)A+�L��2�	A�����&�U�V#"[�I1�wdD�۱��
�w:*�&�yE[� : I�:�F1(h���=׺��.k^��3�2�H�\!�J�Ry�*�C��+g�9��?��!z��|��?S�������"mAH�0�����njV�#����N������Q��FJ�N��[���WP��o���Kf%:��Ć� kM����'�x
B�����[ޠ��=R�O?B3���m�I����coțs��}�
�]s��.&6��)x.���_4n	��Cg���������v��αA���Y�Y'=(4y�ѳ��]�����r��>ު#S�#:;�u@ڕ��#19�*L�����ؾ�x�����h�)�-p a���� g�I�mj�pP6/���@�(Έ�r"cK��Oȏ�{�7R�kۉ��|ᷧD�I�@U������k�������4�mR0b4p&�"��ۃ79w��Hԇ%8���%�Lt���Gր13|��#h8 ��U%����1��2NI����rE�c�Ӻ������XG2����y}�6��;�jN4(���_�ʈL4��	�C�{�h�!�y�`W���O�?�0�dP�s��y�O�S`7Ð�Qᘰ�;��uy�I��m���UKit�D��뺇��M@�sD�UF��P�!�*�}Q`�c���v�fV�2PO��4���y�5$+�}x}r�,Bx��*��J��LRa��x��:��n��z�xj>�%*c	�T"�k��A�x����a�r^�_�_�]ob��L��B��k��]�VD1���J��Q��p�}"
H�/�HHc�e5���HA�!�Y4�]ﻞ�!�p�(���׬r��q ��dVНդmȣ�]�֟G=[�:.ܽϨ�ҒT�[n��m���ȏ� �'dElQ�^7;�w��l���õ�#���Պ�F���L`/�V�4�����e9�K��������t�2b<`��v:#��wQ@Rʲz}0c��Q~/�?�J��G|\bV޶%V&x
I�N&��f�X�"��5i9
��� }����&^��^-����v�T�S���O(C��1y�o�M0���;���&MqO�r::�W\io�%���"�����~5	�kL�<%7&.FL���Jn�i�f�t��L�Ϧͭ��@x��1��wr�;��Z��q��e3'D[B���&`=]ըɔX���8 d���}s�7X�Vw��?kʿk��dw_��7hDމ��)4J�T��G`J�GڡK��NM��T��i�L�����4;�� �jU.�����Ů3+��e:Y[�ī���iG�x攁T�z�!I@��� �*��Cw��3bΒTC���X���D(P��j@����������<r��@����e�K�X�;�W �M^gS((+u�w2H}�>вG��R�)"��)"�O(;��*����p�lW�=]��ʝ�ˌs6O����=ʷf���`D]G�y��iRA�'�ߘ�a^�O�v�ƾ�I�_�����,h��I��A� H޷p�M��5����a�>��t��r����w]ސQ��[z�ޝy�h
�UW��;\^��蟥wm�7�!Zh�
����@�w�~W�ll�7��M�>I�)���g�(/�w�V�	+��hACjΓ���\=G{DU7��>h�m��UG���
��v��+HZ5E���'�v��*�@Y� L,
;%�R��i\�eQsY�!6��+�{w�_�F�������I'�-�b��{�F�<����j_쇣v�ߛ�i�DH�lX�J��4w��2�����[���1�&Z3�P��h�����Nk�6���!X]u�6��޵��;.y1��$���>o�~�I�B�N>7}'�p���nn�6�p�?HZ)(�˟7D��|��m妃@�k������x���\=n�JX��/ �ݞ���)�����>��B������5��<������XsbT,�~2�pwF���
�b�]E���a��±N���X�s�w��RY���M8�>�"�4ԧ��<Ù�i@����J7�|��c�=�U%d��lh$��s�Azy�~V�K=��I{8�U\Q�X~�62i�z�YJ0ô�a#����Cc_zfχİ÷u���s�j�+Ut5=�&���3���m���y%��TF�3ӠB���_��N^_�x�8x�?ď��c�(�Y�
�C��y����#���q�=z���֯R����9�I'&��`(� �P4L��Kmf�ŋe�ȉ�_~�,+h$:�����Ƙ~\���qi����:lT�'�4�J���6h�W���Y�ӫ���B�[�������;�Po+f]��Z�q=�R�@Y�tI�ݯ��2 ^��I*���s�I�j�4.Q�1D�(�ڠ=�7!za���#���'���� ��\��#!��2N�\+������4��M�I: @��s`1a&�6�74�
�"�W�O�wD>��&^�m"�w�>���y:�,�G)dp�};YV�2�j8:q�˷;�<�Y�B%���~!��=.}��X�rn���Ot���g,���������ͅh�!��QMD2C���V�)MH:A�� ^����*�`F!���<�X���zzܗ:�e�O��F��Yg�*u � ?W��� 
/u��Z�2QYxPTu�G	�.5�Xǘ��{R�m�yRU��ݎ�U���#��t�l�> m<����V�@�c@oM��b��I�.B'�a��֡W�UK �>1}xZ���s_�$���0�N�2���I�_��4C��P�p��#>�M�Toѷ;�S*u�Z�'�U�'��>����Bf(��ǋCfn��V���c�(��Z�2�7
��e����f�w�@�M:7�s����&1+dM���h���1(�HF�Q��������Z����@?�&rX7i�3��FТ��1�� J�ݣVL��P�����dvEq�94�>��]A:Υ�%!���P��|�鍒���dg	I,0���tBҬw�PFUK�&�ټm�"=�0P�4����q� ?�擈	p��f��	���s����܅WQ��$����2����'*�T���k6���Y�#�v�V�Aq]BΎ8E��;�ˉB�AkT�@T������pZ�tP�t�Wi�
��|������� ��['��{���n��ʕG�B*P�2#xT�yt%o��.��"I�(�[��[�/լG�@�vj�9�|c�5�qӔ���N����n�,ډ��r�K2��>`�[����݀?zPN���t1�EI�z(ˈ�
����*V�;~ϲ�Q��'�ô=�"�e�����j�H�XT���"n��x.)B��xi����Mν!��DN g�ݥL蜷&�����L��JX�OC����l��a����q3�t��g<8�pN~31�~]'ѿ�\���u�T�/L�:yY[A�Q�����j�1���v*��+AM�L�r	�V�d3p�m�\[-�󤳼��s�ʹ��e�p�\��
<>���t��{��#s�#%��Ե$�rM��͆�S*���j�w~���&�"z��;~�{쨑��>���/����Q��kS�&����T91�2�{�t	�0�U�J� �(�ρ.����nb�g<=i6Dd�vk�6��(�ʴ�s��������m�'$.xpbL��[ܘ��՗Xc+�̎�rKO�p��k������ �G-T77[8��+�]�1������OS9��B��?�e�D{�v-G�l�������V��Γ�r�o����pv��k��d��׈�K#{le
[	_��_Q��UI�08��/��3�hݸa� <��A4��.�UIՎ�w���� ��fL�iz��֓Q�}��2Ԇ�;+��@��B���_��Hї���:����?w?�H��s����!/�23���0�V��U>��?D;8l��Gmk+뇪r� +�K��e2�P�����E��>�5�{�ZD^@��K�a'P����/�$��������z�)���z��ޘ�Tܼ������?Ր'*�j�괊P�Ѡ��bF:V2-aKΙ�B-|P����&�H���k:���>Ơ��ʟ���R��5��{絟���Z��k��V�7����,���z9
���f���;���Y^�iْ�|)�"���}���=���A(���>p�	,���~�m��m'��|�op=�{��M��{1�: �����~�A�r}���,)��t�/�L��ȸe�=�w�v�Zzd�p����)N�*g��lZAN��/��"٫���C�V��|:�'�;�A,T�_p�'`����%��u}��Z$���R����۫�c	 �o���t�m7A�
e��朽����\�����T��[1,�à�"ʞ��}�Q#����Jtʮ��-�\�{�D��#<4?c@��NB+Шɸ4�߷��8U�K�0�˚q��f6@3r%P�tx [���2��4:�?$� n��>G�x-� ��̞Ĉ.
6<3JZv�?q+�D�'���r���g��&6��Zci���MU�4�����~���,3�-�E>NV�~�����j���
uN�I�ܳ�_�]9�0����؁������8'߬��0[B�H��,���K��?~C�82��2r�8��\�������f_ab	�n���>���!��'������V�l�'��7-k�|������r@��al��A�ԷƸ�^�CA���m�垪\<(��N�*P�ZUp�^~,1;��b~��f�o��QZ�J��,\s��{�t_�GOa�+��uGE��^��B�89v�.SN�_��^�=6CM�kn\�r�U�C��;&p������H�=��Ï�F]����q��r�ԲR�h�c�y�P���/��Q�B,�fQ����*��?��ab�¢�L���kK�&�u���y�a5�VRsT&g���(��֎v��,. ��o<-!��Z-�H� rE�K��IJ�ZO���_�-��Q��u�-��1 �QQx=�z���_cf̬U�w����˵�|DS`+\�����*�.�h��5�*�Y ����A4��ˎ��	��@Y��$���M��%W򝐯j�����q�`��L[�(���W3����}ka�kۇo%��lhĪ4d��נ����W#���c�a��l�y��ھ@�%P'�+��Rd����<�fa;"�i�chY�b�Aw��ۉ�O�
��P7hU	[i��
4�S~F���o���cȀ������"�fy����S��`D ����~���N�7yW�����ɻ-�����X�!���#ީN�dZ8�U�����#M���VxG+XR�'��r�����m����m�V�w٘�a���v�_��yWz��D���:�;k��HY����RK�W��H�M�l���jF�H4D�Wy�k�D��̵&Y��tjN�:'W�3?[��t�����j�T����5.抎Q���恫�ZwW@�|�
�G�2�A���'��Jd��e+���ݩ\&�³7-G(>��*R��v��E���Z�G!��6�������vӃ��o�[*��#e벏�Y�v�&lXXy�4D�^إrWO�\�w\b�P��+i�'��t�4�<��6�������sEK���f��dZ&9^᫈��?�,  ��6_*��4���-D�NP�8�^�$[�[�H/%�zz��	J+���(��C)W�Y^W���*���������L��`$qA5�L�,��ŝ{R��ي�C�ϒ�@����tg8��+�]k��V��oj���V�)2�y[�-��IDTc��Z���R�g�����hܮ�^a�]�s=}�E�5ƥ��,kN
�W��^a�@\i�rt���=���Dg$�JL��͉�����µ��Tݑ�3��h�}�.��~�)�� .#F�?��ʏrcd����[H�'�����c�04�#�\�u������񋘫�(⺍h�:�gT�qB1x�m�x6�����兤F��s�G��'vb	De{0J��{�J�|s'y¬)�A�%-�尠u����@�ș�zJ��%p���:��$�F��n��9�-���I��G�X��"�ع����[;�G��y�v�x��V�ښ����s�];�s�bp�j�Гu�i��_Cz����h��*6�el�@J�OV{5��kB�|TMd��x��aH�8�fdnTB��u!!�d�а%J.'�
nva���� Ԉ̯�ъk|'>V���"����U�HGj#��+!�+���\��c����&��6E�Q`�)j���FGN����:��;'��;�I��b"{��2�콵!0��
K�o�Gra�g�m�� ��u���w����:������b'��̨�r�m6�<�i!)�G����Yޫᡨ��7H��>?����*H�M�5��C*�C@�!N�c��\���Y�h �&X�Xf7������<�ڼ��gJ���?e��$��$��O��]��?X�n[��~��<��ǡa�7S!{w@{f�j�$z�[�y
�4e5�ܒ�w���7fО��A��Mb���pc�=�3�N7CT��@��_c���GS���ΐ!����)�$�^JJ5��Y1;�㓃�~�J��h 3����"o tW��CC��m]�uݷ����Q��J�٪C,�i���y}|�����,��ui�0F"ܑ��`+\�4v��>aף��h�+z���(�E��+
�e��0T"�كKsճ��0��N�@p0G5�[����5�YfO��`�,�L<����p�P ����l����-dr݀c��/IX;zpe�H�S��h��5��*}w��m�c�k�f2X������0�^��%�����`u�O�{��<�������jU�
h������jƫ�?���&��#u��f0�"��8��z���֎����Z�kr�T�>���R���s�^w/ p��Í��?�c{G!�3�^��Y�	��2s�͕�۾V�� ����QLo{������,��^|M5��)��₿��_fQe"<��P.��-�r��;�!z18�y����7� ��A�F�`�i�3������q���dAJJo<u��7��9+�<�+k^6}���Ky [���t�U�.��;C�����������^�+H�L�sUd[R�������
�fB�q��QZ(��wn-�݀n=��h8{L�

͛f��k�"���J�+ت���t�7i�X�
�@��2��^bV5�v<���@4N����j1ER�-�I�m/D/�v(�$nF)�"�ʸ]�l�n�J"H#-bZ�ZcH���,v�F���P��2��.$K���齰���rB��ΪU�6L�?c�ɼ���&���u�����/�S"��Sq����'�Bk�TL.�1a�,�u�����.��6{L�6L�>��2�N�g:��݃�T�-��9����<�Kǿ�����0�uݬ��T�>��p��uL(�����3P ��p^�����߽����#g�v��j5A�*ѻ~K5�u� ��x�<֦�;S��U�)���8��#��<F�`��7�!p��=/��a"Z�D��Q���KL�V׋�-��fZ��9�����=1��
�[�).���5��{�ә�j=x��!6�uRԭ��G��Ǐ��kX�0�*�E�+7#�J���{ŗ~Щ�!���G	Ȝ�f��u��~S�;YL|�ڴ!�^C�p^4�	�!��$	�zY��"wD��G~ <���ӫ�d�I��bCdG��>��}�L�n�FN�D�\��l���`��kL��BCp�)�e�!�_�OM��pà���)��d,�Bkk���)�%%P��T�`���ƌ�-Xi�����aht��7�6�,��h�av�ʆ���n�t�ݞ�r������ٺv����8�/�6��ou������:Y����(��S��6#�c�m���	�27�OV�c?��J)<~���k����;�����I��6J�C�<�L�%��g�'ϝ��`!qw��D�T�� nÃ9��4#��d�<�q�fy�V���x�G��.x|�=�6�;y��vYe�x\��X�:���ސ�u�Ԫ�-���qYx���5U���͉��J��8�>�
����V)�(�`�e^6̅���غ�{���e�m�;�t��iE������OY��F�M1U��q�L�!Wt�6 ������NH�&[��'�u^;����\`]$�.E���A��{�L��s���x�������{:�pܩ /1�"áÅ��v�{�����Ň{�ѭg���$�[��4�/�t��Z'�x��닡G�4?�������N��A��h�sp$��u�0ns��������_�4FK�B�ʸ�j�+?�'c�dc�Mh,ʑ	#d�}��֫���<�ɲ1aeێ�A�IWÑ7Z�si2�a#�$p��������'�z�io�3]�L��Ơ��HS���/�r��
�p�S�/�Λ,�~��kq�X��!Ab3��:y�C�~0�u��cM'��U��� �~Lw��ib��{{eD6�k�e�qɓ9ʢ��1f��? )�����:�<ʍ���Q���H��r���k>�[]�W�).�]D�^���2�R��ѥ)�g�d�z��9߾�~��H߳�9��]��Bbޑ*�?�V���9�	�j�z֍�����>�����1�P�H|$mp;�� �k���KFD�y����x!�fw��׆�!t���9�
���e���qg���p���7��p���{�Z��5�|���W�=\���t#�v���0�m���_ڋ^�J��e�:�nb\̀��h4�++R8OP��$U����~�f2	�%d��t3#iڨ<,������p �a�.CR?(��~��:]x��|*X�l��U�+����(i�%�B��Nٶw/���ޓNV9�%:��\Kd�|��|�>�̿KѬ��}(�c�%�nXѨ,��|��*n�D�.*��/�@D��l��K���t�����T��@��� zJ;l���7<� �>`ڽu�(ęԛ��:�v�>��c�U�%��Zb�]&�K/����U��Dp���5�Mm+��!E�~]���m�#�a���PX	�z���ת�~��"�vԩ.���J��#�~��&���p�@]0�&�s���c���~Gm��m?�`?�w=��O�A��舣�oG&?!�aI��+�a	�E&hbxױ拝�~n��z����� 	m�!���������K�ʥ�g+~O���`��Է3��G#�2;��:�������EE���w���:鹛�1�f���o6R��ֆ��@���ӌ����3+���#�m���.�M�1V����e��X�$��q0�^D�;\��/���0Oe�L�+��~Y�
׽�
B"�Y��W�d�XH8��xU؇�Y���oH�0�0�ܾ���^��s�>����>�@}�re�gZE6�������6��i���?�A�∖�@A F�a�>�..Q$h�V�W@�`,�Q��^]ɃE���B���'������_�����f�y��!>��Ҟ=�zI��u�v�i*JE�0Us?�����'W�5��E��ϏK�2O��F��v�j���e�C����h��j\��iKn7�4��-����D�V՜���f�}4�Њ�i
4�m�6a�߰)T���D�^���=��R&w�"�Mf@Y	�Y����B�LbcL�cJ1���Z�ښ#~eH@^��5[3��[5WN<Q~߃o�e20�q�W}��Xņ�/�4q{�$;�������ĕ0>j�����C��VP�F�G�3T�u�����q��O,vk�f_�s����tn�	�fF��ᜰi��3i�!��hJ�Y^a���B�~�a��P*a���d��%8G76�l��]/8Q�Us�hC�7�o3)\�S��	�{"H��R=�Dh���5$b�j����Ÿ�Zq��CmY��4(����V�id��� m��dT\�"�[.BT1�0�4�{.5�e��	�0����W� �xb���.8>WӸnU�h��Fx�� ��	+��"fʴJ�'�R|M:�r���MH��ņ	u�"�v����Aϯ�p����N!�:T-��%��ʈ��l�����JxV:P��..;��Mc��{ibB<��=��&%Z�&�+�F��������]ar�rO�nɂ`?X�݆$�����<U5jQ��<�>W>�+¬$����ک+	R�;��]�ʗ��3<t�+�ǳ���y:�Y�8��M�j�w~�g��C�_��4�������X���=�f?�)P ����M���M��}��#PA�)߬�;޹�� ����_%<}�I墸��X�<ړӀL�.wz��2��I�<�¼n� �W"�����Oxi��{� r�|T��.ٳ9��0����v���������;]�$��|_я��
ɀ�!$�����{Q�<l��\*�b
��q6�'�@%�#B>r̤46Af�fW(��{ڜH�[�\G�~�%�$�C;��W>��캊W���u�%��"�S�Lǐ�?��@�֐��f��O_��: +'P�5V-��^��S��D�thd<�, ��TX˷H��N����K��d�q�hj�ɸ��k���}NMK(�:�B��!$��������`2��Մn�U��t�8��6κ@�G�[Js�g��G�����	[��%�N�^�@G�r;sz�]�.�DIG�x�AvIR���6���-h[�{L����}�J�u����#���F����[�5�#,µu�`v��I�Y��u�9��Y���B����h���5ԕ)�ӻY��'Rd[�b���Ũ��5��R}�x�&�`P�����������F�k��6�6}�dis}[���y�}B�</�MxH9m�Su��r<�ۮ�,˫ĥ�����Fm�8h4�8
j����a�@�IqF�Ц�Rd����{ֹ� �*�~5����O�N%������h	�5?��5�כ+&��,`<��F,#U�ݞ��n+�R���f�0���T%���<�G<(�8�
���H�Wf�x��!c�MnhK�ñ�e�b<Ÿ�r'}��\�@=�I�)�"K,�N����8lD��o������5l��� +&~�)���Z�3���Q�fV���6'J�$�&2�3)+���<	��߈�+b{h>��cĆ���O�ݽ 2+���ֳ
LX�����Z�{�p��ERN�~������b·I�lb�����Ⱥ�^��}�H��{�gW��P4P9�H�6��U©�O.���L4��8q%5�j!ʉ��9br�z��4�N3�W?��n��׃h=�t0��-7|��P�=ɧ�e��r\[�w��-ee@��������۟萆�c��w�� 7Z�Giͥ���Z2~\;쎭��F�~�����R��<�L�d�͢�QT#�Ew��#����ĜS���T�G�Lc�R���)�I����Z$D�s�qRs�lYx(���ط-c-f!��
��U�]�;m��`�6�Eh�ҿ-1Լ�{h�(�^��{3�ѩg�\��N�8\��$vw��O�d��!S��/�q�:��ˊ�� �0[�d����{tg�v�M3��Yi��8����:7�ˤӗ;�Et噢B�G��ܻPC��I�H����$���գ��
 o�z �p&�}V�t�m�0��|�·*b����/�l�_�����-ۂ~���V7������<��\��H.�f��<VE��yݜv�+����VD[�pt�gF�s����ȍ�Jh�~RZ��gɃ�����f�b�%�����{Z�[�Ы�܆?S'�AM
�}j�u���<Q!xC٧�5ݺe<��U���O0�}�(v����x������)��ZЅ��̾�2��zV���jm�%u�Q.a3Q�X��������є~Px����Vy�t��?��>��ސ�����!t��HS��� e���Y��}�)���:m���Ю��QtVXFA�v����e�<K��fM� g�q��ԏ�X�L�����&�����G9V������Y!���qRl���bh}O�����YR6FLo�~!��\��w���PK�.�[Z���_�?S�{����A�E�~�6|W�����N�Y����+I���N(@b:^�e��,?����ëNQ��l������Y�	�D��`6��6�v�az�+-���xE@nI�gT���|F�3}��\ͅκ$I���Ϋ���~�{4n��O4X4���}vІP�d�e5P����i��	I���elX�)���G�Fi�ㄅ
A�6��
!�����Q�E���zK�
����v�v"�V0���҅ �RG�6����
ֵ�i��f���\EM���xRg�fW*v��ϔZ���@ZX�V& �2��h'����yQmަs�a�t���a�2�H/�zu8U�L1i� �ƔG�B4k�L&ޱ�՚Qmb�+֡\�0�9M��
�;��ԔY���i|%X���.c�\���\���<?�Xm8�*n��<NzZ�.�n���������?T7b�	F��1�n�e��>u��J�h1���Cy�R��xD�^��.�k�> vb-�Z�7���Ȗ亠)�8NI
̝�U����.�' �|��-�AD��:�����O�����^y��a���(�q*�oS�ܕ��/ҝr�����Xñ�Z���:CC������M���C�s�	V�}��<[:�!;�1�n���4܏"�T5��S�e�T1������>����h�w紊�̏��gf�Ґ��;t j��XRmķ��x���;��SL�vAD@���S��;�>���p}g~�����NŐ_�2u��>���/�T�&v�pE�.uƞј0�hlp�8ڸ��9N���t��[�c�rf�BmApy��B�[W���7�
�p��W;����b�.��P�f��#�S4áeJr���F�QZ>�I���&	���`Q�C�\�Q(����Ȭ,��ƪ�X vz��<��8����V����\5�6K�i��ex���Q��e�"�1��P?�2��2kl�����kZn1��TI]~��ﷆ>ۅ	�牘��o�52����n(�����Ga&�S;A��Q"�}���
��NZC�����#%�D�u�Lw����#y ��L�P�5P4�m����\~.��,�1� �ͯ,�	�2w�h��1iϸ
�,�!&�We��F="	#/	�nT�#�#͉xK��B��ȿ@Cu�s`���o�8~r`��*|?����V�'W���	��s����j��Ij�WՇ�yX�y�C�?N������������g��A]��מ\���fT�J��9��e��$����*e6���F�O���2Z��6@�sc x�^A�7Eݟ��Vݧ��u�[M�	A��E������\|b@n��B�܁�G]!j�i��{�b)Z6��N�a�̏���8��E���0�/fp��Y�`UmEQz�%����p��tW�K��'g��{t�A�m�Ʀs(
�r�\Ή�M�l�1����l'���8�%T�k���G��$c3����z�µ�,�D,���?�Ϩ����}�#M�+����Kn����|P5Ɏ�c�7�d�����ƨ�,��N��]��Tg<��
?6[�k#�I�u ��U�;�"Q�83@�7:@#X+�t�k��oى?o�J�hܒJ?���"�J�mٛڪ�n���j�.U�~����?7LE�C�@��y�l��{r
�����q�1=�R��!���`Ӧ�\���놞bG���*���Q�c�g�$�tFR#�Q�2��:�"�d����']�)�C/6 �u�e���ojܿ��Xb��cBk�J��d��w#�-��cjsq���yt���wƏ��v�Z?$5PO���F���b�Ș�	��$!�)�?:v����G�3Ʀ�ڙ�Ef�-���^��sǳ�3k�UE��p�
<&���t�	m����x�����J띯��x�F�Ue=:��|	�A�I�-,�!<Jd�nZ�6.$z�N��Q��u�(�J���{81�Ok.�<��[X��4� O��"{)��9���U��x����Z��.5
#d;��j�|pp�(�a�SW]ڹ�XX9���%�vw节'Z#&U���g$�A����UN���LY�\���β�2;>�nۇ+�*�׫N=	X�}�~v�r#��θ�9g2�H�u{�Vљ�g�5�aZ*$����o���@_��/���̑��6����&��5)����Z4N�&�D��k���]���ds��魥��m�ߝ�sk3nC5{4����C��7vo�ȻR`�ӧ�kRA���&�K�g�������=�{f9P>F(\H	@}c��H�}ؑ��D~�Ѥ�	���<�7��iF���:i��	�^�Y6YBڨ���(��>��=�o,��Rw�zC�~Xu�l�>"Vux\���3�g�е���������fBC>������0�:)�C�\g���j��{�{fV����ٛ^rc��A���JC�N"�z�����B�3D��$�K���Rw��G�y������=.�G�$7 Mv�q˼�U�un�$TV��X��X^?�ez�ی��'t��g��-��P0�:�~Z�{��t�9\z祳��Q�CR�0F!>����4�&-]�mAQno�����BR>-�A���*������D�p܇�מ��@���2�!Յ��`�gA�D;�t�WI������K(y����If�na�{YF��2e�!����vSf�]s�2ږ	Y���È�+qW@�� ��Zk��r�����w�W��R�c�o�L�Q�뺣�~+b��趶�����FV�Ct�Ĕf�����<�c���%f��m��Ir,M��g�{��I��[�$ g�ز���J�������ԙ���Yf��·�0��ro����n	�����ɽ�oc��*B+ǉi	�s�~e�]�bڂ�Z�G����Mb�s�Ʀ������+�;`_b$�#�W	���􌇯��~O2�0v�ӯ$躉���[�
B��$�4P��|�!��W�Uф��οO�i���{�����)6ȄU"��4,[�w�q�{,3�m��9�G��*z<G�@�/�a<4��G��ģҸ����Q�����H����hRǀ4�,��-�M3�7Y���^կ�� �n�����XٿZ�:{�?!���X.��^����A���[Tڊy�V���4��_�����G�­��:i�.�9�	/_颧AJ,Xˋ�,���d�@"�\�� ��%�W%�%ߝx��}��_7)��;�����륉�g"����k�E���va<�b��#d�}E�y#C�!C��l�O�I����|��.J����?] ��L�Z�l�ݞ2�H�&>���J��w�Iy�볘Q[�pB�7�>3�4����3�vE��~&B|x�
Hl�E��`�,�P�e����_�)� �0���x��Ӳ��Ԭ��$ׅ�Ӽ��vm���߫0ӱ�:����
�A�(�ߵ�.Ѣ�* �;��v���X�w����bM�R�D�O��.�<�)���xp��o(�ff���-�M��@3���x�}�=�XMQ���>ڲ�3���ģ3�S�Y)в|��֭&9����1.H�+ �N���$(|� I���Z�\AR�d���v�1�,��]��{��/jxp+�q����)*A=��9�?
B:4�蒖�����h�Y�ڊz"�hl�r� �b�_[�'��E0�N^�M���*>/��
퓕�Z��N���{������՛j�D�O��>�����>�0�b���'�R����B@(���4����PuZT�qnzԬ�Z�� c��@��ɜP����gHB�i�
�]@L� ��s�#!��3#��ގq�U�ja_"1��GY�xW0'�_����.�<�p�$�6oXu����b��LGS��!F;���d�r�N�F�o#}<c�]$���馉�O"�O!`)����T��?O��S���g��7l�~/��cA��Z��{-8NbWy�b���Y��
�(���L~^�2a,�-�����s^�ч��Z]�QVG��t���� *c�f�;�lB]A�O���m�Ƅ ;i ���"��#|4N��{�48�[:覐��n�B���xM>b��M�Z�O�7nBR@�i>F�`����T1�-F����P�|��v{��ŏ��x&���!���+�'�z�커��5<�sP�R�"�O�i���%���t�[d9|�|:�̏�8�KqPͧ}v1�>���I�8�|���2H�7a����.�/�&���ܦ��{�7�c���&�
=�9����`��m�A�B�n9C`{"A��;��U���z.H�>j��I�e~;��o����i�L/˓��G�Z+�dr1+���h�*����"�y�A��K>��d���g7W�?�)+`�?RLn! ��"���%55�9aӰP����!Un��?��:٪4���@F5���"☝a8�H�VХ2E�+�VE��Q���|V��R�l�0��73�i~�tk4×	|8�� �$v�)��1�ŏَ�5���/y8��[�b���Sm1��\�Ң<��w7"�t�;u���ao�̶����c�� �Y��O��0��Z�Վ���E�z���T6͕6� :ц��� ��Mk7T5�z%�<�����}�n��ߡ��p�:Y�L�I�"#��04��$0[ѨvO�t�\����l�<0w�Ґ���	Rn37Z�گf�An�sS�����u۩8�H�9�<;z���M;F g�x�)!�W@^�؞���l�Fñ�����Jd<���!�oսn!�S�-&j��B�	��T�AfH�9�H�}>g�n�3�+^�X8]���ٽ��?�fR7��]�֪Q&uh��x����ut�)�p�8�h������k����%S���"�@H�ȐDo�?5���B4^�ۘ��Oya����+��/�$V���1��4I��^e/# �`1�ۑ��L��4�(�mPkn� �L�iC�P�Bh�c��E� H.o�.�v�5�������Լ�iҶ/��R��)�2�q��#(*,�U�1\>M����i�չ��3�_���O���Xj��ݢ��;�(����y�z�G~R�B�ϳڳ�I1��.�կ\��bH�<��%2p�����YԴ��;��P���*�\���¡Uh�Z1kt6�_�n?�6FM�'�"T>o*ޮr�<p��b��a5��n
g�A�m����HZ�����Ԯ����>t��Y�������a���&�w���9:/��K�٫�!�8��$�~&����g�X�R�*X��e5OLCZGL��5Ik�&��C��o��@[=�)�گq�z���ŇZ����Џ�KyI� I�d���>���j�z��ir+���*��=��O��� ��Q�Z���q{����O��c�M��sa���S|Mr)�}�{{����,`�K���M��]��P�t�ɗ`�r�S���_(���9��b���[[�&@���	�Cȴ�b�.�	�׮�|i��Ҷ�D���гSF5@�0��~��3Ig�c�o��K%��r?Q��U����_󅮷�U����g6VZG̹�'�#��
�.��b��*s���ջ�Jꪧ���r:���A�\�:��fHk�+	$?����
�Z�L���}��#f������g4E�5�5��?3P�u�2��Y�S)��(�]HK�g�F�ܟ�����k[��,�&���WG4����F$�Q	g� +��=�ò���kŒ[���y��~;u��=b<�s2��3(%P��^Z����y-��\��@����߽���մ���X~/n��l$�D�\�9�
���RZ������P�N�]^G1�$zc9�ՁJE~�ш^˅�b�A�"�`���̬�?���;�óԥ��+a��	5�J2좶f�^ƿ��6	�(d/p�)
,g�T�؄�]Qd�q��SY[�bi�����k83���WF��$=,r�n�@$D�yUd�9l�b'�$&��,��
{cR$���{gV��;^^2�8��A����1-�F�`�&öڡ��, ��\���k�J�5lC�,��.9;���E��,��uA�7^*a�֖e߁f_�������� n �1r����	��i�����&��������2]Z�|ʀ����Enq2ѣ�O���q��ރ$�'�V7-������G�$J��߂@2�F��F��,(�_ak�L��++8�g<KB֛�f���+4c��Ր��#簊�}�4����b�� �7��E*X=�^;D��ra0�
��
q�n{O���dBc=m��1������ֿ�\�6��DUɐemaAGIE#d��a~B�ٰ���ڌ����Q����@�s ܵޟ� G ,�vj졝�xϓl�Q'����<9S���T��W���a������,��*�٦?�߉Vºd���YIڀE�H0�^�Z���R���3�1��o7�|�bߋT�c/�����ulX�%\�˃Ycɰ�p��V�:��7�c'O�
q��/�T���I��}��6���qP����*P�6�V� ���1����}k�cq$�
QX�R;�O��O�ĥ7�� LI[��SE���=����x>���]�j�덼��̶�7�wpu�DŃ����{%,����;��]�1�-��x���$u6E��6��Wt�ʺ�K��eֹ�6�	U}�h�%Q��^l2���2vg"�����DMr���3�	��ֺ24�-�XF�LZ���X�h�ф[ w|������Ά���5�#������`�v���2܁jC��Ώv�g+`��']����y[ݐ� ��e�1Q����4�m� i*���}�Ú���ך�W�}$�U]��y�c,���|>1yz9 6c��A�3!K:�ı8�H��`�Y���H�����բPl�zdH�1mJ���0#Sz݉��ŋ�=� �y�����Q|��G�ǅ82+�MPJ��#�h��Gi[�o>�a�m��'Ԇ�I0��p��O������+�ʵ �O�C�'^���V8���M?�i���S��-��F&*�򱙸T��.�p�Rг, �~�yd���'q��C-���D�6mNۙ#��?�ќg���q��Mc@?$ѽ�����#� �HsDՇ|�Ū4��-��hf����y�4c�Q1_G��a���M�B�ȻO��^#ƶ��(X��gjf.��^��쵢�^����_"�
�����3WF$�y���tz��,3Y���.^Z��#��T!F��ȹV�B�񴠨hz Ǌw~��X�S_�\C/M��V�M��y�u�	#pV���I@��E�b¥�I����@�V��6uI5�B�3!_��;b��|T�T�����2G��*f�O�6ك}1�\���G�Y�6�-�oI�׻�cfv묍3�%���:�Q�:��%	W�����m�J�J�b�!�w��h�b$$x��@���ʋ�V!4�Rc�3�9h�4��z����,LI���������s&p���x��F_�?k�tD҇U@�5/:>�Y8��Ο��Ԁ&��̍�ɽ��$:l��UB	^0P+H�`���};[iN������E �Yh�����}�%�,15$�<��4n�ɔh�~�zs��:Vs�Z"���D�f�,r��jd7a"j��X��,<�bڕ��74m�H�ۄ�4������az��4���2������fL���3L'� ԴeO(>O^ՠ�e���=�����w�_�O�4.�\&Ҋ�x�,ƨl-�������K���=^�4��w�x�C���p���xwV|F+�X���.��^��ي�I�Dl�ڃ�W����I���j谍����L��`����!��/�������>>a�	��p �yߣW2��+S��*��\KV�DH�`�+&���JC\؉�M�ی�_��R7/��ϵy�a�(�KN����J�@IE%�A�� in�׀S�@�;g��� �������Rٯ+�����)9���}��r�X�׼���
����&r�c] �Ui�A�]�����;u�3��*����4�E>/�H�s"���4 ��xO0tc�6ۛ��)��n薯��Ý�y�+OYpk�]���6HS'1��CӉ�.gn#����i�!�/A���n4��p�+S/
��J���K2"����ΧZ���{̃�T4!�0�� /k2p���rø0�	gyN3���m�'u.9U	�]����v���lR������� 3`�e�"0��+��J�c$�o�������Ϟq��\���
{�h�u�;'4I�y1"�Vl*q�:�W��/��'cf-a�I�b, �v��{��n���M��|�
��0(i�{n�r�ͥ_�{��+�Z�n����.�����3���p��:�>}����䟐���ݝ��H��B���n����B�h���^��EA	(s?�� �!E c9Lv�ۅ*$D���ěG�8�f\��a�����غJʠ�D �+�u�d����Ix�E�n� ^�B8��Wv�.W��
s�۸���iK���� �cV�	�:bM4�w�=�a�s&�)�]�/�ވ��^�=K%7F�lѴ]S-
sN�Q����,̜�SV�B�ꑅZ�WR�K��ʗ��0��ve�����y����r0�@��W~���/6#z�'2I;��@���t ~��Էߴ�J��V01l��J �r>U=�4Z�Ο\����5�L�mYK_U֓y;�;���ݢ �7O�9�R}���N�!cT[�9����Kŏ���c��\ts&��A$���	��o�^� ���ڊ�+�G~�=;�>�@���Ͼ�ۭS��M}%�#���ng�'�S��Z_�y9ﻀ]祽vxa�TtX���qVFN��uKn����4ē.��}�/"�M0`���(�i�_	w�_L�|��6�in������4#����Q�k���M���$�oGH>Y����9o^���WT4>��o&P���S`�QJ�@"������f�O����S�3A!���R���\� ��8����GUr劵z�n~���B�++��"[�9�,�����A��OFO+�,�t���WSվ�AQ�0����HMn�ԃ!7� @c�A�)�+�(��t��1d�g�݈�3��[���^ԍ�!s̗/�w�sޱ�ɻ_�C�?۠j8L�Z��D��-�����j��޻�U%��ժy�w^�����Es�[b	��\W�������+TS�v���l���i!.D+����@�q�\@q$}��G�K)QSq04�=��tꐸ���+�Qj�\�5�7,L$���C�� �,���n��3PU��`4S���v!�v�ik�/���/1N�%�3�'��d	YDj�ܳ
\G�bA(b-�ʗ�%�p6Vy�c��8��D�Hd��� �J��h�R(�s��0���Oi��(mkD�'�#��Hq�j�fk��E1��D�_�w֍c�h��0�n��޺z_g�e ���7J� �� ��D{=��<�)A��d�%���M�Bs-�$I�K�zj����
\,T�)��318�
��K��5R����t���z���(M�@���'�69:Z���km�@z��'�ăF�	� N_�p�X��⁀�X����]؉V��D+���WӴ4�>�	R��V��̄�7�'�A2ae�Nu<�f�^���H0�j��r�[�:���07fܖ���+��;�6]�WX�I�ՀY� ?�*/�jx�](:����� Z���V��k7��lF)[��!��qav�Hjw�р2����0�H����Т��.���R} ��h�UFG�����+π&(��cP���+ |a��Շ�<������l�(�w�v�"��ӽ�p+x3��?qN��'�\f�胩PEG�N:gh���w=���NUKb,��,�[���s8d� (�$$�20�����kpe���h�o�����q[a	�꣩~�w$�����u�c�m(���`�����,sF�3��I�,�@t�0��Pf���"���P��r�6�����Z{5��Vz�,HF*�/���,�u�Q�)�+�ݣ��~E`�0�}Ns3!����?-�E�;�@�����/3�4$�|k���ח��^E���x�p���PS銣�}����)����7�h}@E.��c���Bܒ7kF�("�ʘm�c�v�n6��{��ߖ�Lː��Av��ח��OY���G��h�*ψc ����������Ŗ����{�'��G�EI�B�e�^;x�����
!s�^b���`6V�6��
8�:^���G\"����"i���tVJ��5"|���.���Atf��A�K�N j?��ݔZQ��8�I�Բ��x����ߧj�m��^���bO��� T�@ $�}�.��B���>�@��+�R߻&"�|�F��8��
c�[�+c0<2o�yf_2v���Yl�ǡ}ݫ�tp���͏���x�n�˽5�rb�8��u���q���L/$�8AդF;�ct��φ��26<X*K}��_vjo��4� �|u�7�4G���ڑj�a����;u��4�*a�V�	 �������Q_�i��>��*]�>��T\�#����������tKd�T����Y���x�x+�`qu���Kz�1'B{ϐ��A#�Tq�^����-�S݀,��C
���ְJ(�Ż�Wu�zDn~��*���>$z�lyZV���l�r�� x���a'AT�X�����TMa|�~�$Gp��&�|U��������Ȣokr ��nM��f�TkX�q�&�T�w���@c�Gb�F�UZ���7��{'����'�H�%r����޿�5u���Fr�e*�/>\[l5�|T:iwqm�<��ż���c�z��#�z����7������G��~��F��bL�����{C���4��g5�Խ��`g$�~}'7,������qv'׺��|��!k�~R���>�U��}�/^l�ۋO�N�#�q�y�e�U�ɖ��
�Q��S�H5
�i�a��>fꦠHFa�M���ҁ�� �;V7̣� ú�����d���kxUH�����j�g�>[��f�?�Ռ�D�K��8���C!��l觱�
���AA�@y�G�"�2����L4�x�M��wq<	��=��!�c˼
��m��ӣ b2�D�+h�b���#`@N!�nm��)a� �JR�D	ͨ��R������Mu�dd�i����c3Vk[m����$@�4v�*u�dG�|mj��y��Y�#� �7���`�Q������73���L�G�=����l�j��a~ADR���߼A��1�Z�R��V�7�`Sp�Ч�j�D5c�q��$�"_��c���Zo�4�d�;^ޒ����HIE_���j�Z?����4�S�d��00���+�>����<}�4��d�GIEi(��.ґ���?������y�D~�ܨ�WI?U6��q.�� 4�3�P[i���e��4���5�ǩ��O��jah;��5x�`S��bX8	G�Q��K�&N�5ְ������F�VO{1��-%>�nkZmv�"����4u�؃��m�\���4��7of1�8�!�˅�px�2����c�����2��{�g���V+��^�^s;�K�)ق�Hg�O�mD�� ���ftVA�"��j8�llf��[(�`��ZK6Ʋ��W�
������������o�Vvy ���:����	:�J�9���N{m��Mٓ�\y�iI#�PfLU@s(}j���࠭vm����Wֵ	�G*�����k�{Ǒ���]<|hL����(�F�#��g�]ГV����k��6/l���eK,��fƜ��^����ssL��u(���DШ��K�>���F�?�	���?�4"� >�.Y͊���b�7�����;@q ��`&� L��2���	�w�j��Coٳ(�\�= Uj�k�����Ĉ�L�c�D�"���s��4�8d��}�Bl�Ý����Yi7�"��I�L��-HݚUiLO�V�oa[�z� 2{�W(�j��/��P����� �m�\���[bx8҅�O�#̊s��(��x�3U �:^ڿ��{�hT��r:Y�F�����M>6���������}k���T�(|��j�f$����ap.-`8��{�Y��x��>.2 [���D�)��F��� ���D�.�'��fu�J�:K&�X�m3O�)��o�`��Mn�P=���Nk���`�
�����Ժۭ֧��	�yy�i'K��6Q>�����jQsH޻�^1Vc����[XU�S���Ģ	�C�*|�����2�WNr�)�	7r�Xd��q�Hb�cF|"��2�A
Ie|R%��۷w=T�6\á��s��r�XWG�6�B+|�����B�ܷgV)t��h�����W_f�tK�A��w��כ����ߝ��F��G�����$��T��D_4���]���+ڡT�m��8w����P �w�V���o%K(�l:�p�\
��8JM�ڤG� ��\��	���	����k�(�# ������j�0���G��S�����⥅��h�v����/"@0�wh�VQ�x9�,�(��P��B�H;Y��e�q�Y���|ؠ�~�S/��>5H��'�jk���X]zW�P�bPs?o�Ev�:ݍǋ�\���q&/f~1�B'�
`�X��>�����oD��p�(��)̼_�� �$�����x������Q98�|!|?�3�lz[:ZC�fݤ���J��F����Zg�x����o�C�ŀ�a�p43������o�c�n�H��������7D]��3��o���6Z��g����*���5?b��dcѦ�9���fU���������L
So��0�{�=�Ԕ�=K'j��5��#�.iOh��"Cw��N�R�l4�Oҥx�n����Tti�]�n����~�݁���u�'��%��g�X�k���ܔEB�J%c�?0c�����;k�"� ��J�1�,X�aփ��<�f��y�S)��>c���	w	J�	�6��A6�\Xe����i��k��Z���xLT ��N��m�ݍo���5�CTF_��䇟� ����f 9��i��f��	�uaM��L�LFX��d��Ag��Q�X������%9�a��7,aK�q_�v�(���NY�~��̡�|7�{�lB`鱐�Ͼ:d��-Ͷ��[b�]}E+�5L׭����~�W��m�M�c�_���B��Q�yd��L�]���ᶷ;߱'zI_7r�s�7� �?��h�Yh���#y����=2t��
"��w��P�]�ݖ�.�hVW�\��i�ڒ���9FӸ>T�{�k�5�Ū�5�h���s��A��m���;���^�+k�w�h�)8�: �<� [��"��M���������p��s�y�gվ��εYͻ?*�I�	^k��wb9W�G�
L�r�2��d}�C�/��@zXۨe)4C�1��F*X��� ��&��&Wu�X\��Y�����oٓ5K�<M1I����Dу@�Pnu�lM3�Ju��K�ꇒ\�O�@��s�V���S��+L �޷n K�
�}��>^R5�*�Ɗ=~��a�,fr+�EMz���3�C,G���zj��EU�<��ۤ�U���m/M��5XRhxf,�R`9*nX��h-u��/��5�u��J5"ƒ���"��8�Ԡ�z��_�������T��S"x��t}mZ�т:���yYu��1��9�o1��/AC�f(����Z$���߀Jt>��<�w=�U.�$���kD����(��Ӕ��2� ���z��j5�͎0\*��	g
z���K��&����_�U:���!Y�&��-,Փd�,�_y6l�u�o����J-�����1?m��r�3gj#�$b���粍G k�y�hHP�/�!���KE�-�S�I3̃���r�A�x
^�u�[	Yvz
B��B�U[���Y��ќ�D\o��1����p	`�<C-F��Q_H�:,�e ��t6Ġ���a�B�4���S#Ymy]c�TS���jn�.�?�ECة��h'��̫x�u���*"����\C�10��XFB���/Ύ��������oG����l �jd��ߧ{+S�>2�,���Y�d"@��Е�K
����^NW��0��������M��<�!��ίӻ�Q2��FbogF#b�B�h�+S����¼� ��	���h1�CY��D3�)iŻ��D��;���(�]��*Q����[�A�H-d63����!�O�O��'����z$�t�mpA��=��j.
7�6Ǻ��G�E�H5�3�?ZVW'��a���=�6��ޒJ�g�����L�$��=t�EN2�; ́s[�@��|��������]��[�ƅ�� w汽E�7���M^�*���H�
3�Q�N��~� ��P�t�!�V�^�
20qːX^�u�Z)eK}Kq���TZ�B/�ܠ��P���0�BU:�p��g�"�5Ȃ�o�������[M\��+��ԉ>r�v�����j�qo$�nU=�����4"e�v�c��% Ь��%5��]Z�2
��{�9�r�-eѺ�F['�U��}Ms�UAı�HK	�,�N}�*b^${9	����������l;/²x�� �5�ɍ��{�۵ɨ�[$hl8Mވ33�g&�'7�-{�56�@@2��wqTǖ�>�C��K��}p�K�n���+n����,b��s��1UX�^/���,��z��nO/����cuޜD�o��(�U�]\�\�����}����!��jJj��ϩjUKN�������g��J�8|���(��Vrɢ�ۧGx��wK�ͤ����v�i�#b���
囉��`r;Naj��/�E�H�C��i�hg��Z-sC]����E'����DO��=�%�����uȁ�~� �0�CK�,ZͼT���j���i��X/�M�@�i7�T�O=d.�u��p���uZ@��Pl��w6#)"j6|j����q�>���������n�++���R\����&�Nx���:��7/�����+,�~�b,BjK�p�Y��l����A���|c���}&c�VgW��Ň�iP�U~�y��To_ ak��֓V%��q��w���PBӐ�%N6�����3�	�,"Z��	���W����^űE@,-*�A���WsZ���C7����ZR�b�.<���F�����4���s����r�i�8��,��&�[`H՜U��a{�Sŋ����V%�m���c��Är����i�:f5��ЦY��|������q�vJd��7�����e��?V�Z�s�X:�o���yLi
  bƋ%m�96<v�\�\���S�	��Q�$�@b]T9��1��2]�CG�U*g�$�N��gU˴$%|������^�XbJ7>�6�����l��-y���2
z��"�&��5FĎݷ�� �Q{q�N����6�>Q��\E��Q�[�<�@L~ >OqwZ�k�fɰ:A�A�k�'��\��cX
��=���+�gl�� �&�p�|K�y���o~])[:��x�g�����h�]�N�~�T��dN��0�MZ@=c���*|bļ��vW��������Q�g�7K�%���Re�Je���9�A�v�MP�"�$��j��
O�zn�CNg~w��p�x�7��u-.��z�X�a�'�d��eR�5��#�(�cA����W���Jx���F5]2�d�e(a�5¡؂N��\���N�!����}J_����X㏎I)�#plf���8�ݍs<��U�f����lԆ�e�w�~�.�+��>�nC�������* ^Law�����'�l���d5��\�zkT���>���q�����l��	�@̷6g@�ӑu��K������?�'����(.�J�;[�	�$�㻉"d�C1�:(5D�n��|�&����7��1�?�BVj��Z�"e�����%vI'_���-n(��寄yȊzU�͞���V��>�Gnek��L��ۀ1[b�ݥh�Ha�*�[&?�[	�^���c���k�^���"�O3"����s3΋�b3hЖO=�� 7x�t�y�`�LK�<̖2�k�{T�&�������S�R{�Ǫ��|���߂���:�`g0�N����K;š�0�,!�vr.�G��Af$���V�e��_$�����Z���6��咡�t؏u�r}�E�E(�f߂��'a�Ejp4>g@ɖʹʇ�z�R�	rE,F#e��׍�.\^�e�Q���"s6����un�Mآ0�m+�^���`��Ҫ��	t_����R����t��L��q�,�}0�ưx�z�j��tS]���Y�^(d�uIջ�Ĩ+}�
�-t�no�
:������ �pb�ػhF�c������(I���}�E=QO�=R$j� -�՜�@0Ϡٲ�'����|F��m����姆����*��5��}#�����t��Ħ��r��K^l6AL��E���ˍ�og/��{��*2/���a�D=���BCD�mlH=��ksGI������/ نۇ��?���&�;�vn�+��)�(c��/�w֝�C�$[C����)�	�-)���n��LFn�{�,�C!>w{�~[4_��d�7�׭���j����X�(��SӝΦ>O'�-��f�$��ǜ'0V��]ʝ�P�(��h�m\�o/�Tag�:�h���d��cb]��������bQD-VO1N� �pX*S4����h��0���xS�Όg��ŉp��"t��ő��C�D�����PL����*�W�ЯMn�"�(���&��x���E7���q���/g�ٚ�,�8�43��8�|8��u#� �!QCB)A�ߞ�	:�P��oS��\�x�y�(��ȹ:��ئ�t�p�п����!��H/�k��zyB���N�Bw�{@�&� ��Hl��V��Y|7`1H�#B>������!,������P��;��o��
X�T��9 �Q�^�+��W�Xh��N���)�=O�����bf.� �-�SZ�!{����V��GP������ ."��h=��������c���l�eQ��AA�X8�����rO3:+�Yx7���MV�V��7�0�&��Y�9x���
�ش�H�G"�v_�,w���+9WBρT(#'�x"��Tǻ����w��vd��!B����B�8dA8%.�*��BM�O�����o��"��� 2�~�2C��X�jN�<6������ؐC5%a�U.��˗m�5A���fz$g�x�����.M�k��M�1X@���E���`�a�	��]��"�>h_�d��f�p?-���±�l����>V��T�I��*B�����o��z�5K��E��3�0�¬Y�H2rv�$5�&Ye.Th���q��~w0R����;:��Z7�ee���$\k��#��F֯dsp&���j����<r��5�,�3��\�:ҟ�;^Dn�S>��/�o�C!�e��M0��a���w���(EY_�$3�
H� �f8�yK���i��M.T�P]p��ka�bBM�@
;��1C���f��&��X9��}1iP
����3�p� RE<�>;f�HΜD�7[��e�xx$�H��u)�X�<�GeI"+�H����z{��HPO.O��*�)�#>�?���T��3x����8���q^+�^1L�U���?-�l��N��4čGj|Ƭ;��J�̣ٙ&�\�%���3OX����kn
WA����FO�x�ϴ�Q����N+X��W
}�Ƕ�SΪ���M�FĮ��z��o���p3%�J���VG�G󳊍�6�ps�;Fb���7�1���X����s�ͱ;KZ´6蝸O�V���i��o�g~�9�f����#�z%o���T 蘵P�۴��!��-�~�̆]����o���;��=�A�ȟ�;�ܢa*U��&6}T�i(�cl[uW��n��-e���L��+�dۯ;���>�h\]:tL\KE������n�ٲ�<��IB>1��%|h���gֽ�����a4�/�v#@��W���U|U��p�t�#9t(���v��mt~ W�9���6�������pu½Ě>�7ptň�b��B��͋�����A҃-/��g9CUd�ZԞD�����3 �i�K�2��u~^�(����0Qm�����NP:�"����=��]5˄a�S�?q�d�ㆎ���u,�Z�z� �TTI���s��V�M[�a�X�TƴFP�/��4�N{��)�P�b���*ZL���*M�F.�智^%��?
�����+P0��d��Uhȱ���R�tʹ�Q��n��~�D�\�"�K��y�_����!��?��#��������H,IjA�쏁�q�=x�\��5 ���4�˱c�:C!�p�G�2��AV���poC훇��"�"7�G�UJL��z+���<ʗ����W�
=�i9*�0As��Z�xt,�r�7��Q|۱����Z��`�1�����v�f!ҞM5^���k�L%}��"QXiy�ːgB>1E�sC��b,W�N���)������r��#���B�P[	�7�@ƨ�7L7%��;~/D�n���&�#� �,IE��L-���[,�Y��l��̇
H�?�U1�{��w�9�I�x����B��5)���������Ц�(ǭٴ�u-��Ȱ�XV�8wo1ì:�@H�ݘ���e(�GȏPE��DT���oL�|8^3'?�:��P�!�zZ�O�.�H�m�}#�m��Ny��\�\�
��9�vD���!ҽ�"ME׻��w�(g�k��ٖl��6���o��I\;N!`s͑��u&6��( �5�9�>s��߾���\�u�e�qg�d��繟��� (�m���	��}��}��)�@b[<�$[l囈ᙕk�©p2�<&2���$�p��#q�^�P\�C��8rn@��p���9�/}�v��v��*�i�G�Q�Ð�U	cc��� 1�/�H���0�9�T��)V�:����
��	
w��od�u*���Sԏ� O3;+�k�i�̴I��5�Fa�F�S��ͽ�"!.G��#0�Z5=�h�5Ct�$x��t =�Bpq8��5�k��ϫ.�9�o��٫��5
wvy٥�|����(����4-z��_����
5��*�-����"���wU����+���4�LNB��*#��M������vm#ͱ��i_/L�����G)/G5�@�Y/_���:�����#�#}���w�*!��3'
`\c��	��>�" %W��1�&�K��Q{���|]a�
E�C�=ܚʪ'��f�ȿR�nْ+qSS-�#����#ǆ~���&�c�2r��&G�Y.`�'��N���-��z�ёh�+���0���?�����
�={�X��I2Ѫ}��Ďw��UR�-n���UX�����ⰾ��;�ElM��O�#����B>�������5<���)�,�fl�0x4�L��-q������ L���<�������=�u6o�m'�7->��a7�	~�K��$��;	A�j`�R�����_�bx5���yXu{��i�t~No~1^,�0�;���3=u�Ti��E�VD�C�0pX\1�w��mS�;�5f��z��h�(�%'�}Z|Ǫ�kg&���xȊ�D!T`06z��X>N�0�/h����<ˉe4m�J�F��N�%��D��)h�7z)����$� �-j�Cٲ��pc�i�i`��\�6����c���B�I׽��ӵԑ�-WW�RU(e��zk��a*i���_�����@t�>�b/�צ�sy��f!E�h���)�ٗ��,T��k�du��b�2m{K�j8ʨ�]Sk!69�J+����}x��XЄ�#�2��+� ��5�S�I-�c>�t>ҙ4���@ca7)x�����e�À������ ���nh��wc����BQ�I�Փ�����g�EV60�
B���0���{�p���~n��v��M�7|�4!: 7��K�Q�Ԩ�������N�>f��T.����9g��ŹU���vlM(�p@k'��*~�9�܏��%/{�tQ�4u@-���i!�~zħsi�a��ʴ���jx��l�b��i��)�����-��7<������Q9����e�.�}� j�t}/��p0�߼������e������-q��Bp�Xj��M���!u�8ʾ���t�����_x
����)t�C��'H��3o��GI����O�E�O²�r���xh�{j���Lkn�G�Э6��3<^ӛn��X�ӆ�~r���wi���/���S�*x���̏Q�[w��62!bq�e:"I��s5rO�Z�홖 ������h#z��cQ=�o ��HT�����>��=�*
ƱcxJC���p�����|V�����/�m4�wZ���\p�c�Һ��!bH�^�:�r�<��~B�W�/G1x��j������x���J����?�p|�����n����D�	ь��hD,T��Q�"]�P���Nr��_(g[����]��	�F�c=���c7"��@���֘���H6����Qρ��H�#V-�yj���a��|∸�чI�#O8�ְn�v�h��[OD��A��i�[iL#�ˊ��0����Q������?��Z��6�X�T�u��"@�߹,$�����J�o��B�%���2M���u�|���I1UV��&@��g��J�`}�J� �dR�.7T�B/E1[GfY��܆�)�d�!J�U�+,�C��0��t�i���5D燐sE=eL$&�Mz)��U<;��4T��$���&3��*���æSR��j�b,3�͊D�8�����u9�o�I����k���F�r��1�1PSt���I����Ec#���͓�n��1O��e�����۲)��'�:4|B�6;Un��qج�a4*R�(�
9�����;k2nBqp����̘��
f��}m ����Վ��,᭷���̤�.(ܯ�	������Is�~ffSq�c
��V��%�JZ{��+�Z[sU&�_��l�|b��c�cW8eOz�Y��>�r8���!A��/���HZ��a�(}����/`e�le�,�3̠��bh��|��xc��;"����!7I?�J�j!`�)�.� �ߵ�fv�="Z/G���C��_�$�L2.�$Xe�1�knR6�6Z�RG{�c �"�܋*��ea#�����ף�Z!;1'�u٥o�O{�����U�j�r�ǚ+��A���q��;6�-���~&�x�3o�,��uT�ezׁ��A���=D݀�s����r��ϕP�6�zt!�3݉���7��r��S��-��УK3g*�Y̗#�x���-��Ns�i�[˚]�,A�#��L2t��� t�с� �O*��v��H��e[e\� �Y�9N���z�B��,�I3� B��$�B�ٿ���p�Ѵw)� u�)3C�V�؅�ߧ�-��|`���k{�Ѕ��%^�7"{���ME��UU�q
�O-��O���&4��Э;��PS�.aw�I�˱ocɠ�_n�õ�0�߈B�V���9¼	���O��n~,+Q�֙=��+w?�3��J�н�{��[(��so��'�� �S�ur��40zy"Å�)2����#.�D�~�;�=���57PG�~��5F��d��C�^t�J�3�a-��E��y�6F;��*G'�&;@նI����>ci��i��]�Z��XX�Q��}��|)�v�<�yDi�`�M�q�8
=��=䑙a���5u����`H���TM�i3�R����(E�5K��GȚ2|O[nz���GǛ ��:��!���Yu�'�?��̟�����' v����Y���#E�T�>si�fY��a,Ԝ%5��^�A��A�J�4`�i��G�������O�v� G D��5#f�g;����"D=j<R�0E�.�`��kExB���Q�S6?~ǝ��5d��.���)��W�~����^J������Ͳ�7��>���Pi�JJ����Vt�X�_a|��'�_~󒥹���Y�T{G����3�ǥ���eh�%���~����o���;SH�O�A�'�/�^Ɔ�>,$�{P���A=�J�]1�-t���՜�B,��A	�~P�ut��cr�;�*���\_��-t�����n	��@�ܲ�� �Wk_{��q��(��Wtb�D���C�Į��Y��:C"�w�Leِ�l��X������>o�o��!)����T\̘d��hn�$J�y0x�P���k�V���k���ѿ6� �~Rُ��h����4�a���UWԧf
'�a"#t��(�@-Ŏ�[��Y�4V8�B�}�y�S�{���+ǾO/�
��wR�D0���sI�֗�?�@^?�u��Zx{�����K0��,�j�{�萵����cd7n���]��������e��ik����	@��ʹ���	6#̐v��c�ϔ�Ԋ�x�d��ڳ��+M༄x���v���%"tD8�z�:x��=a	b��:娷�4k��aEX�����7+���FJe����=x�Q��υދ,~�/�6��S��R.�,���.t�n㯇Y��񉿩oVM�QP����k�ְ	�a�̛�uї�����W,[���p ��#���j�7��� 00���o��@�`�е�>I~.txd���hZ �(n����Q�R� '�~���v4 o����ꁶS�%/0���E�/��\� )�M���E/�H��c���k�MY��ɬ�A��`h��EI1�� ��D����8�����%����)����������LYZ�6
��AeT-=�X������}pm���#BSx*�S�죯�!)7�h�����]��j���
��`�jD!�M)K�a���ə�A>C/uk-��Y߈��)���K�Zs�6Zvh�7��둞n{�Ό;10U�6��6=����L;&�A۸@s!����Z�*�j̶������*�{�]�53T����gO+=�;^4eIZ-�D�L�y���|a�&��1�[�܋��u`� c�!g��O�b��H��<��)�T//�����^@�l�"�ȱ��t~v��T�e��M�B�r�ݔO���cն��-/9W�)ԯ둷�m��?E����X�϶[uHĮЕ��������c�y���Ŵ1��M/a_��r�b9�\}����m����#T�&H�h+\�
�jU]�"�ߍ���Oƪ��� �'c�Wć	> s������@�z�V)Hw�H[
!�05?Ek{�B��' ����I0{����H��J����N�ڀIWH\�\�i�_s�����:�uD^����!�Rw�R�_�[K|N6��?\Պ�\�Rjucl=vzQ�;������=Iv��o�t��x�wK���i�3IeB%a����o�;bq�6��F� /�K�a��{{!�gOԠ�}[}M��T���b2��ݼ�H� �L��y��R$�H7%L�LaԺ$P��G�? ���<()nՆ�6�x7�Ko���|Bm�r]��y��Ap�m~zy��;N�8,YK0j{Pk�Ĩ�6�N8w�M;����Q{�e๟aPޜQ���Vǳ�Ba�¯ó ��1�X�ޝå�Aↈ�~ꘔ2�}���qۊ5�d�7fP��2Ċ6,�nP;���Ǥpn�wTY҆o��+ ���P�҆NXM���Lj߻֞vpM5��7��V�c!7��t�g��y�F�D�?-��4�Kr�]-��r�k���3N�w��*�J�(?g�|rߒWX�g���ծ��(#0�����`�;b�j#�p�.zjl ����1>��՗��Zu���>��8��a���d����XS� ��o�W��.��=�V��ZT�h~~�F�/��S�gZ�I� /}����S(��Y���u{�* `��B.>��!�D��n�J���v��QRp	Rǳ�>'���kq� S�M��|@�������L�fs�z���U��!�ۮ���Ӣ�����=T��-ρ�q{8��eөG����Ϫ���%W�9T �m��|��������i썝�t����!%
�L~�L_�i�����gq��+�
����>;�fTA��o/�����8S��J�!�4���3��m����xF(�1�>�'��)�a5$��}TT=5Ȳ�������-��(�2V�pKG0.t��cT�e�N�`}��E�!�V4D��V�*lz��>����w0;�;_듿5���E(v��x�����v�l"�5�"qp��C�[��- �P��;u�n��DBKY,J�]�	�p�B�4&g��ơ<��s��򠩹��ifH�vO�>�� �_�dA�o���h�Y��o��,���R
��n[��t�;�A�#�W�2B�Ǽ�[�և ?��;�o�I����7��.�m򡖛b'�a��.��� �[F ��݆V5a�l�����Q3=��R9Q���y��mt�#�U�}[X��ɓ��?5��?lT����O����W����Rh��̓�0��q�0e��CT��Q��D�6�Q�?�h7�h ��%Nb�;�����J�L���Ue��.�F�L�������_r��O�6�<GFmp#�{3�o��)�k@."SDK�j��sil�����M�� ����`t>SׂV�ʽ�m��ZVy�
�k� �AUב��Lݣ����o����c�93�(�6�Fk?Q�i>zu�1�4-&� ��A����B�0be)��\��������/0���fOݼUEݧj%�nv:k��l}��H.��l��Z8�/T��Ѷ�IoS�?�!ي.!��mq0�/�;�����4#UW'!�S� Rk�˒���$,�3f<u7]n;+w��æe$����(��$�MTЍS�gk������p+�H�,ߤ��4�����RV$]	'j���?�
�`�ڒ4YVF�Q��	s�6��x�oP���1c��<�,N�<�0��n�;�*������~������hC�@��M+"�Y�y��w���g�< "��ͤ��n�A�r3���Jދ�*l��%��W�sڡ� ��gJ*@g���^"�b���_q��W�!B���Fv�������;���(b�F:��ϕ��k�}�Sb}��P�\�-H>��S'�D�ʨw%iH��;=�'��G�ne�Տ%��0T�OH��O�I���X�DL��<ѡ&����J#�!���Ֆ�"}���/5l�67�[)�c]h8�\���W_�r6-
��.��y�mrk\JGS
 {C���gkg�)��V�D�;��J��2^����%oYIZ����*��C(|v�9��d���q0�P4[���&"��--5 )�i��H�"m�jw4E|M����b�o6�h~�ŀ�����o1��p��hv^4��M���A��1]�o�*-k�-C���mY[̟9�8��q��jA����lAK�y�-:f�%�lq�!�/mBO9ˊ�D4�J�H�gY�ʸ�I�9U4�Wm���?��bMw��
7Kc�42�j�6D"i��f���>��"G�9;�Q<`qKj�R�m̊Ͻ*�\V�*f$+"�2�;�M��Ǎ2$/E� .K�h�����	��~�!�_WT���*�Pd���ư�-�\���P6�4��{�b�̠͞�dLO.yY���9_�4(K,�!�iߕ�W��Nt���X�Xz���G�j������т]��0��C����\��H�/uK0}��ԥz�y;6��F��$�ux��Lt��tJ��ߖV�� G�]q}:\t*T���z��R�����d�C�t�W�rCBĈ��@�!9��lG�j_Fr�����Պ����qnl������u��O�>�l'�����>&Y�^�P�.$N̋2?~-nHU�g��EL�9D%!��%���N��Bg3L���yW�ݕ��	�����3��0�j�܅
s�����Z)�Id���=��cWT���Z�9��E���KNz�
^�#D�j��txɟ�;�{' �E���W�!��
7b��w~���gn�/�v�-̆���o����=+�P'��i�)����ұ� Ǒ��^�����͹�[N����v_��f��&ݰ8.e*����k�wy
s���]���J�Dh�vvh)#��G����q���h9�Ct�`�{ͽޱ-��碊8>�L����x
�ŗw�vTj	�Zg�w��ikG�a�K+<�F���w����^��C#˝��8�A��R�_s`�L� ��w*�V����C�v�T��C����twY�Y�#Ի�$Q�Wj2y�+��M/��<;�Wz<w{د\q4`<z��j�.v�I�{"���2o�Yr�� d_J�t$v.{��~]z���m|�&���W��)�v����7^�x����q�4Ar7�
�e���\^ȥ�[��$A0�7,�����d��ms��QAP�L�i����M�u?sU�l�	 �f���X�}�)�C+�Z�c�+���G�EpÈ	(	�.K��Rj��ʞ�R�2g� �y�j'`��������1�7��-J���%���9l���d�fjO��j���c���#�M�Ah�����(�E�ҿ1&lY�~<��o�94m2��&���c0�B�� �4�(���lV�F��ht`GxK�\�5J����q�O�9aW �͋����y�����K�w��R��c�O,1M�L��/�ʨ:��x�E����!u�j�'x�,h���	ڞ�Rg�hF�IȾ�1NF�B����t^J�����(]�$`n��K�7_���AȊ�m���t��j���������r4-�R�ם�(wi�o��tve�u-�Pr�,m��ݥ��<[�_�uW����2����,Ύ�"��d@lR���Ӷ�ʛ�k�Q�����rLܥ~K.<Z&�� [ٮ`W+�N��V�&��k��#D	����Fb?a���ݼ��=��#�nDܻ}��Τ�1Xj����R�O0�N�z;�?xyw�*��䷅�ܱ� Eg��Oc	���u.vx<�'y�H����[ѤӉ��+IwC)ܦ����3R7ϫ��F=[O�=/l�kK��Xu]�jNv��>gHY#:hQg��<�q$RPU`���R�Z�T+F�S�tMQ��w�7���9[�x�Ie�R�2���ϒA��H����B���D"h0�9-$[c�Z��{���M��`��r�IA��>ol�:D.��I�4=t,�Ѷ�_R1��?$G�����Br��CG�ا}���^8�ɻF)O��Tk�Sў3��tXn�@�i�����w��l����ꤩ{&�KM�?o~��I�V����$�:�`!���
��D����/F�����8g�\���1WM��ʚg�d������|������zȀ"������9K�59�{2�T�I{*q�Mh3ex��;�1��-�ǡ"b3&sO
f�MBa�vYe�\�%aO�׮����p�u�v�����Z�5���Vl�yϯ��[�wd��Aku��u%�Un}�������RR��xj�s�Z!HE�i�B��ٖ�
�t^��w��{��W�݅��܄�n�)qj�fΪ��-�|�r�TJ�Ǽ�ꄹV؂2���)��	H�C���TP�t~��n��>x@�cGmq�h�U�JDm5B��s�t��Y�TC��w>Y��r�z���Y|FH��3)�����/�:�>�/L�>H�(�x����@Y���5�ZԤ����<Y�=H%����	$D��PF��`0��F�w����մ�uh�g�$��?^��)�8��G��'L�������@c1��}u�үR�{��|#�e�V��D��K-��5ܴ�na|4�7�,\N�$���R�(맢��PQ�A�WKp�Zd��AX������~u~4����@��J=˅2�4�I���u:�k�����o�m��V����T���&�돡>#ӛ)Q���cr����7�J#;q��T��M��g5$�w��?��>�B�~(m1?._���q݃HV{�q�2g��j6r���nxA�ق(�R��ˀ�q�+32��*�1$ְ�C�gM~�����
	ׄ���@[���7��g������u�ˉ���z�t�BmG<6�V���'��w5+�_71ӉN'Z��'K�lD�X\�O�s˶�Ђ�\H�m!��3>ֶk�i;�����-u��n�J�`r�D�2�U7�t�s���nzc�4�$!o� L�y�jHS�ʏ����%�+٬x����}̈́��O��/�����u{�v?i�\< 5L�>M2 ���qp�4�*���.C~��'�T�L��EPdN.�u�h�36���L��:�:tJ��0.��w�m��W(���,�r�b���"x�N��=K*zq1\�aQ��{���D}p�I��������~�����2�t�F����Hɪa�7|k��̞���t�� փ�h��ɹ_ ]�t'-m�7�s�Ʀ���}�Ȑ�S4�zs?;F�#�֟B����F�;b�����ι2{x��_K�*:j�G?�֏s���n����:B��]�)s��KE7,(y���F6N�`K�#��Ԏ��� ۶Ӟ02�asm�+�F;|��$�=�"��2Ω\�K���Ƶ!^��Tc��4X��<��KzDZ�����0�����e��2�D<��2�)�ZEL���Wn�f����-��c���Iv"ќӂ�8�F�ܬ-��uۓ�k�QA��EW7OzЬ�˾L�@��a� ��"C_SF�[��t��h���I�ַ�f���?S�U'���I#'$Gt�v����ڍ���歛3{�3�Ժ�/�쉯[^�>hx�;Dé��GO�e"�~X���F��%x��xe�y����{���� ��D��O��D��6$�7[�\��[��.�^�`Y���J�&�o8+�K�F{G���(滯*y�M�g�v2���}��m�2f=guU�N!��
�͋�s|��#ǐ��Ѐ�@�S���E�s+[߶,v���$��^s�O_4��^/Z��P�����Km�[��g\�Iƪ�w�`��T����K�L�yf�L>��\<Ŋ���u��5z��������L��4���M�&��Λ��DFCJ5a�L�l�m>��y�����f���̰���[�(0�$�AUA6���v�83Ŀ�&�QZ[�Ru�<t�:�N\lh����\ V�0՞�:�@�.֑��3�~�f�TS#}��<�t���̝7��xD?�O��y��"�Zw�?����/�nwB�".&cd��qT&�Jl�
�d������R�'�V�+j���dZ�c���2���4�ޜ2�E������׼%w]�go�c���s�RC}�i���j�F4���K�� �o)ֵ���A��	�d��P�#g����9j�v�C%�$�<MJ�����Ǵ��Too�I�K�@��6�u�̾�H\ xR�ȩ;$Q��P#���0�����z疐���d}����	���X�'b���5'2G�'W��( �Uf��uJ���t�u,M)_�2��ǕA�D&�}�|���<���N�7�U��l�j�=�\�;W�����]f���Q�pc-rk�ۂ����	H�!#1�W[��Irg���9|C;����7=U!�w��UG�$���Uǌl��I�ù����3_H�B��*0ɫ���e�a%�݆�+��uY����l��Z6�g��\�r\-����M}��n�TyAx���)u��|���8�z�(���vl�0�q�J�1�7]���
a�U�+-jh�X�.��dQe1q&�I�b:��`�K1..�*FG. V-�o�c-���)��y�+��}^9M�x��_�;��׆ȁ�+��o99A�˯����j�)��a���D����(�T?���e���`�?��ř���dX�L`�BKL��!��T�*]�8b5n�ݸ��^��W[�
{��U��h��4.���� ������_0���V��̌�^e6�?�B̳��I���7�Қ�]�>&���)h���-<	q�n�R1�;1F��0T��Q�5[6�=שIL\�2۟L����
.4i�kLU���Ev]cD�6=+��x���X�L¸��ֹ�x��y:z/�#Ȫ�~��T���J��c#���FL�]��6�Y�	ao�����z�un5�Nj����&9"+T���#]D���x��'�~�5�����&��nш�eߋ�-'�X�Y�#��)���Y�3KA6����B�]j!f� <j�<WШj+1_)���g>3p��ʨ�ܵ�3�����T�Js��.�c��͢D&�E	Ak�!Q�;�,˃�rQ�o#r��6����VU��O׳ٴ��5x{ta��~�v'��P�z8PK�n�V�������6��:�f��+��KȜUyD� E��������u;OU�{ǀS�Š��sU�?bZ�f |��t�k�yZ02�a3�&����풳���Ͽ��hC�7|@�X@!䇅�F�:���b�'C:�*kV�Ӝ��0�ęf 9е�(E�g����A��o�ְ\��F�zC����< 9o�`o��^l��}!���P1f���!\��_�,&�����\s�W��QP*�?�y���@��Ш� �������}BE��J�C��D���!/I��ކ���*�t�o�N��Q!�"��w=U������C3�c���`��@��Zpj�6��W�5)��(�6�;��aLWSw"Z ��O~̯�z�
� ��y���P~�;����#��b�v$ݜ1U�a�jm�a[����mh_ra���"�?/5�텛�0g��s3� �z��:�S���r́���	�_+lV�J�2�ϟHM��M}����f���J�U�ϴ�ZNz�C$ ��$�UՈ��q�k�K��j�U�2��]o��ʸ)����ހ��Se?j�������B� �;9c_����X���Ps��L���n�����i�����K$k��]��CZ!$֜�o�5�Tڢ�v���d��&� g=2�2!W�9��2�"�5�{�X���տRLH7y���T�8�����ƹ�O�0qt�l�.{<��|�6�"Þa�nqg��	���3�C�E�T�׷z�sw�������o�l ����e!��_e�3�)��u	�n�ӈB�3�ƴ���WiF�Օ{.���k3\f����L�]6���u����~y-��v*����F���yY���� �~�4MXS���{��izg�?o����A�<=e;Į�N�5Ċ��e�b�e�U��L�{��a{�d�4R(�B�?��0�����`���ky��o�!�d�j�sL?G2.3 #�$|�l?vpc(Ut���
�	�A%ۈ�8� ���,f>��-r�y�~d}x�����$v��K��f�;���#�����C��Jw���R��Ǫ@߉��Lf/��
�g�Rȹ(^��������~R=�ڄ�?�p2�oW��Q(
�D�Q�1��}�4$�ĩ�><��+��Y���U��[bUל�7VV|�����;�?��b����Y]=*�H�y7�z�'�*Ǧ>��ݎ'E�2�z��a�ЏE>�������m��r�y9O��j�q�Wh���5�v/�]��	#��$h��δ��b�=9�pxz�u[���"�`��p}��It����,���%~�1�X;�t_iNj9�p}'�����E+�ka�B�l��4�1p�6؄�*y��7���d+騦���p���R���ae��J����Ck�4I��+�G�4�v��A�Ӎ�����=2����6�����^|��#"e�6g��k�"S�w;O?���b��4�L��O���^�k�H���r��^��Sc�P�~%�0�-Z_���W�I��汵pC��i`��>o���ȷWV�U*Q�Y�YQ=i;U�ޤ!	�2��:�-=���@�w�zPb��&UY������z�n���\�Ox�*l%[X���eƏX_��%��B�9���Q�;+J���&n��5,��ugۂ{���2�\a���P�&�2u��d�"I�~�����
|��{C�Wv�H!�Sf�Q7(�I�u��!�~$�z���w��}t�$&Ϗ2\��0Wz�t�-���{>aeA��mT��q�&Ӽ�zBk}�'5!��׼�K�٭W����nw1�������p:s��v�:��u��y��NhJ٢��a����6Dks�/�9�8��Zq�ڃ%޸u�K|�W{x7���k|	�m#�7ܡ��yO;�����ߺ���'���f�훉^r��#;R�0�|�ew4�tH0�����@d����ǷH��a�s�K�+�SlX*�_P~0r��R�	�N�\dbU3����0kA��dF����4�c�?tA���S{��$��<�+�(K0ұ�y��8Zg.?���A�Gv�$�AN�Y�@�g$���i?�	�DpA�	�ʹp��|�E��3f�ڒ�^E������^O�Ai�l`���8��>�� �(v��9 �=��������>CTo՝�� 
�Mys�ĉ_�gAoIK� ^G��g,���N����:I�#�}G;� %��R3J�_���*�[Oy؀��od�����1 �Yv9��	�.T�3�%c1�M�K�������8�ke�ݔx��Tk�l�R`�3���[�
m�W��j�e �>Cm��8���fg������(ZI�qR�����OZ��{sт+.bַ̯1di� �p�V��E�D�{4�W��ݏ�w7��G��h�M�(�Dx\�I�*w��L�8럌� y�-�&�� �_b@A�q7��m�BzkW���R��{}�Ŷ<s����*#>zQʀ�'� ~N'��_A��8�_�ڙO��U�m��!�eO��]��i�'�C�/8��g;j|_�[5�.���4/��2֬�?b_Nyl�㈋fY�FR���=a[��x�ĨБ*x�����o����^���O5[�[�V�	���YHCR�"�F��堼a�����kv���|G�M��"��i1v�H�¬`�Pfi=��%0'8!$�����������f���Wj�Qr}��(+�B��XC{v�2ûu�.����.'��9�����\)~�d���djƏ�o�O{?��K�
کWb+,�=�O_'���۸��~�*��?��>a@FP`�N98x5�_�ׁ�p�#��x�L����@
��v�~�140�r�?��/�� ��$�����<lq�mc������񂅏7*`v�?I:$���(+�B-5.O����,S 8�J��8�H���(	v�"��%�,���-y��K�I��1xy?�%�l��YI�"Z��:��I��E��u"W7U���Q(�>iqvX��G�w�����ۥNK��2�JB7 Z�F(D���'x�kID��S��l��ݧ����;Xo!LnmD%�c,/�!��'mX�Go�m�UőE���&��6��Rho�7y��8� ��T=���+	A7.?Q��Q�:� �`k�����[�x���Ni/��=r2�i��/p��w���u�]�S˻6M*���a^�����wa,��T�]����9z�6���S�;��(���Gp�S�����U��܆6��H�L�(/��"&py,����f�v�H��Σ�譄��[T ��,.7�Ïq hb������|,ђ`��u�/����[K��qΙ���@���-G�> }�a���^�� �a�ǥ8�ɬd;Nw�8��}hT�M��Hv_�Ы��P��a����ퟟ���\.Im����v��@m��ja����z�k���
+�V]�(�<G�'��Z��C���㰜V��:��*���y݈6t�V��V., 4����'�c�'v!��F놎1	!Qy��"�Bk& ��r��MJ8}qM���`l�sS�9��<��g���r��y�����8�GB0�UK0��U�ҡ�6�͡C�`p#l_�ѩy�H��O�߁��E։;w�u`��b�k���*����H�'<�ː*_�����a�*��ր�q8�*m{XE- ���c�g)]�U}��m���_��CJ�A��Yj1<w��+d���1��EO;Z���5�M������b�8��=�
�*R��0���G=��j߆�m�T���^0�
Qo��2U��]�̥(�0�+�1l�K�LwpZ�)�_�J�J��2��R�\�M�>��45�e^�P�U�!��WxE��Q�s�)���*��E�J+Vp�S��"r�(�6߲P1D)���4�HE���Xƅ���$>��O���6UC\ڿ2�j�քn0�*_Jw���!�r�{�;�����2;��Dy�tP�=�r� � ����?by�D�y�H`,$mPH_h�A�HYT���5(�4��:�L�̱��OL�Ȯ����#�sW�to��Xpovؠ��-C3d����q��v��Ɵת��@(��;Mb���[�����:��$V��B@�����U�*�
[���������u 9,�;��6pK��l�������k"�c�U��[kt	�Ӭ�g�)�ۮ�y업��F��+�Ľ*�%51�3%oL�4:Q���yQ�� q�V!V�NTl����:<��F�~�0��2��S�cz
��m�}!!y�w6���ޒ�����v�yu4 ��		]�������{X,�כ`��6*7z�_J?�����i�}H��6/7���Ud��3�n��� ?�?uZ��lA׭���ZPq��Q %��[W�N ��&/j5<�c��w��9����]wl�*�ÞL�z�-����I���&aLW��.kl�m\���0^���?��Mp�9��Mi��rl�*F��Y�}�K�]%�=�?�9�ñ��߇F.GU�wGB��{�'�	`���Y?�A�I֬�=e�4���Jꨲ���B(L��Rdr\��.���0n����}9cpP[n�˚8�X�>�1r��R������u<�y;Լ[)��|B9�l�^��R:P��x�� �ʢ�-���N�R���2�<��Ɠ�s�Z�U�3/
e�J�5�ZZ�*���;{� ��F!�JhX�p�V�|�6���nX:�l���'�
zе�E`�!i��Z�)�fO U���-�KEX%!I�o�ˤ0�N�,�����Ic�d'�j���Y��O�0�W��Z%@�C�L"ۡȋ]�V�	&<���%)���+&�r�鉜��	��D0[֮�|D�`��m��}��,<%�x�?�\_1nz�9���X��]ʗs�t�5�(<J�M���KJS��,�w1*���|	ꁫ�j�\"�������D�?���SƯ�B����WN� �r�����G"mb��P�ƣ��d�k��Z`�Q�8��ʕ=DϟC�6���MR�(�c׃���#%%�Ht��Ms�-�G�q�p/w�,��l2����~Y%`c,�7�J�K%�0�H��k�_d�l#�Ӳ\^?�PF�K M���f��>����f���9V{��9������ l6F��$6f�V�Z�/x0F<��#qp>a��M*�CZf~�9��}h��<,�Qp�6�(��1w�3yg�W����X�j�'�-�k��m����jPѤ�糖���jD��(dNQ���W�������2�v3�C>�C�$�Q�2��P�b����1�40v��j�}�7�֭ǃ�=>҄.�^W��&�ۋ�~���z��(|+�=@��}��{a7��F,��f��G]�g���B_"7[���;N
�IALmr�ʬ;!��1���P�*i妅���@f�����>�f]@g9�[v�&M"l���s�(�KT�!KM8�Lx� � ��c^��ӵz$�R�v�D+Ks�j[����&��i�	�Ԡ\����sm�߰|:3dk!�xl���u $�3P��}�.�E���u_��x���2�Z��F&��Ϲ�]�3�'�(|M��#�Wzo��񘘮o�������!;��2�.ə�AK.R��z�]��ˀ�ю�z�F�I��#���m��J��g�ہE���3��\�9&�c�>ݿ_L����M������v�jd<U h^@x[Կ��&���?�5NZ��v���wk�/�`�WXxFꡏ�"_8h���T����kR�nOni�0����y�� �򤺑D�����}&E�zC�R��Q�3Ob�crɰ��Urɵ��̈́���MR�P"�b���h��HFu,I��x����I�����`��.������&��1��-g�A��`2��?��g��<j3���ʯ���u���X<;%��M�#6�i���uw�%jo�4L���W��~�)Y����Xc#K&9�RT��� b)�Ȣg���_�K� �����g	$S�h*�d�ud&�:U ����"�����,M �]Юv�A��=���.Q��_F t8z��!��-#� ��Z�G������J���r�	�����=�b��,P�&�kV�Ҧ)�?�1u'�9�Bγ�I8$ >EF�R$*�����T�R_�@^�68 KD �]A6�$��?C�I��k�SZ�/�au�����A����O���O���e�RC�S����]�;�����U! U �3��J�%~:Т�&9$�&P�1�	��!����w>I����j^��﬚pr��̂7�H���� �C5S�C�+V��xF�$��i��0#�IW���z��L���jۧ�����U�(v�O���_Ү:�5�+�7lj��{�\���kz�k�ȹ"#d͵�g��ώ~4�����=�8Ō?EN��?ݙʤ(.��#t���5_.h�r�cx��Bx����A����(Z�&��q�ޓ �K��~,�z)�Y<�sy3Z��Vl�Q	l^*�q&��&�K�RA�W��|�����e���]�M}�H�g�)Z��y���w�b�?� ���^�Uv�w�剣!N����˾��¶������M����%<r���!������o�<9��d^\~�OsÆ�����M~mBL��BARw�,Q�H��2���<!��m	sӔtbL���p���9ى�܋tf���Vl�, U�K��,���H��8JI�+{�)ZJ�#����H��뱷b=Q�]����Yn����!ZD:��UC���͝�-��H+���A8!#�%w�v|��X�w��w������ь;����WR믨�ѽX`Nk�ԡ�n�Bi)��+b[����b�<����`1���G7�.ir8��C�;�!	�y�-�M��H����֢�����Me`ޭ��8^����c���G�+Ċ���?�ɇ�~D���L���CdZVxc��@�Jg�U'?�.PYl���h}'�Y9E�bK6 r8�x�3��,��f�A����O �J������i�a��`$8=$���3�ʹz�l�\=���>�������.�Z���* �}�9�����p^��2���E6̲9���"�A{-���/tCM`]�%���W�mm�,��s#.���]����
e��a��vgtqٯi�%N�wiqz�=��W�.�w�,��T�k�w�d������"�I^A'��o�UK�ӹ���{����٤�/���e̳�?JT=�\+	��+�0����x7�bኼ���\��S��d ����;�.]�yn�y�o]��t	Bp� �B��,ZO�b�x !C��/W��D���aʎ�H�ސ���ؼ�`�
��|ZsZ:�O���j�bֈL�JZ�ڶRG�aL_v��!�$�lo� �"+Jl�Q{TJ��FڪW�죇���	w���<	he��I�v4#~�ID��r�Q$l�Z��;��e����L�����W=\���^��r��[e��|� [jR���ұ�GA��v5��y�SE#K�[Fd�9��*�4�Xɶ�����y�+�I^%�rߊ��3Xt��������o�~����k._d��IF7л�5I$��]F3-��ɉ�`���s"OL	}O�'0��#@_\X�.��S��b!�p�'wEd����4�P�"xC�嗹�x�@�����	�G���+O��NKPr�҃���@0�.|�"�-{�!F"~.����q�&3=.���6�����Ə�u�� �GA�o!.�Rv-J��Y`1�O[c���c��&�%up�s.�5[t+`[{@w��y�8d� �96y�����hi�Z����۸�U�bp���?G�Ė�fq�8G�0,�n��M��߻?)��T+ ��x~:��#n�������Bq�0{��5"�*l�մ�M��:%V(����q�]������:ٺ.�4t6OQ��S-�R򥲶�:p��-�8^�����J=����{r6�}G�����W�����+R�KZ���|�FAE�wZ�ОB�6;��y�A��� ��@t�qc������%	��uK���n\F{s}sb�1r���k �it��Y�zʈ�u���(I�(�nd���.�9S������Kj�(�3�z�JG*��l��)�lFml�!7�xg3/���ܒ���KOy��]@��	�>2́2J0PI8�z�2֢��ߏ�*��sB���Ea�	���A"�T����T�Ԭ�@1lIB�@'ǢL��g�����q#?�����D�i��/ը�wCcV;�Ag<�,�Ю�&&s�= Q#���?����Ѧ�8�>Wt�Y�M�Lȯ�%��~d��I-���"H �qBx�m�Ϫ�?d�玱�L$:б���#����$���Z�"�7��yN>���?�1n��!�%�H�:�]#�JkR�X1R+��j��QC�;�S�Tx� �o(8��Q�1�K5���5��0Os���p��!�!+��$�P�:�4��_����B�jGy�|g�
Ƒ�QCe"8�ע��Z�*+ i���cRJ�P�4��5����*Х)a�����5�Xs�6�&0v�v~F�*�D����o���B����AH�~w����[���F2���b2��;�C-CH�CV���vh�	���Oїl�ds��g���̵
<sK� �;#�eƍ|_�G��u\��bI�?�����hjH�(X�e��Gqmt�#�*�J�v89��QD I���]�L����HQ��y�h6�)ů�5�ɸ=�3R�X�qHW�u ^�ϧ��3��#0�:���TU/����_�ԏ�8����0Y6_��(��Y�ɏ�{��:�F^�۟���⬄�9�[n�z=�Җ��a�?�����A"�/����M��r��ӷ?%�Jp�Zh���:v(#�;
>?r$j��M�"($�f���8�n��cJ�\{:	z=��j�HxbyX�m��Q�N����$s���"�9 u���zО.���I(�rV�;��+V�;�^�hq���ߖ�u�C*�1����
�f#N_��pl�⊬yU%3�5� (�pN~�/�>Q!ű�ւm_�%��'���	���e!R6�#�1d{���Fa�*�MyN��'VL�U蛠 ��?.,ָ�&�������T;?U�ՕF��J��'a�nmy�v�@��8i��u��EN���VaI�D�M��T4��~ n%Z��Re>&�5�q�DB�2�w�v*Qf�&�}����۬8^Թ��v���Cߪ�}b�U0�3�Uk�1�eK�!��ˀ�m����$�O۾��ʔ��f�$+M�X�[�c��0C��AՊs^����mQy��x��U��eVz2���uݬ������j�t���lH�օ�S��<������<��qjT�j����?��k���x�sW�Í�Yq"	tn�K�{��e��3�p ��� ������S,���7�lLB��j-��]ѳ2�$h���X8��=Irr�> ����z-x@߀mw�H�W@%�%����v�w}��z i���V��W�������!�~W7:�azkl��ћ!�e��`�!H����5�2�H�-�ȓL� ��7M}u!��)�)N�V����v#<ID���0�*�fS���#�%�?���=67��)L�F�:���ۯ���D�7f�ͦl�I���T1B_Gq��{m������ո�z�>X��0��d��XZ$p��B5��aJ0�W멩9��"��6�	!vQ\I���8��,!	Ef[-}�����{��k
!8w�Q��JP�����"���.�ݎ,[L�p]9�o�m�}jsGau}F4���v�<�B��~�~�Y<�q�	�{�X��fM&	��������S!��Y�uP/F�2`�b�w���.'e���C��R&���5���,�z���R��l��,S:.���ȷ1�^�~�<�M��Q3��_Juj{LdTޝ~���K�ߠ��ON|��k�r??��{%�&�����h�e��L�ҀMts!k)Q�d-���F��!�V�N����fA�9�ZL�c�6����p�h��+��G�zߩ���EX6`7-��5&�b�Yi�o�|e5��*�{,�ep#ՙV��	��1t��B���~P�{!k���_�t�y�����h=2�����㌲�3@���Վzi���q}�DFk�]%Ya�C�U�ZȣX���g��M
�H�����ƞGk���#�l�O���=cҦ�+��q}y���Aş���|E>�d�l���ƞ��h\d��z��P��s�A���a���<������b>�8I!�� ?
��0o��l4u���.�!KBQ��`Y�����P��r�-�۵qw�E�]��wJ�y:f`�A ��M��l+V�qy����n(yK��~�i��tL���E��e흧0%��Y��,=�x���#H4e�M=���t����ۍZ8��h＠e��������9�,���l�'��!K ���x�̴k��DBt�O��3�&r5�ۡ��yu��y2uL}��t����&E	��]g|��D�����v눼_1��A0�܁�d"�wkG�ϫ���a-'�s^���z#��lsH�������9�����B/~��pq��@�>�URt�����LZ:ҟ�]/�\�J@��Ej��8q�T��{zl���ڢ="v��Z���3��S9n�ӽ��,d��N�hY��`��^vZ�T�B(�8���4Y�W\�좪���m��A�n˂���c�g�҉/@�m
�)gB�_����b<���Śrr�E`��]),�%l(�E�Mn�2�]��A����\�]?4��3���@��T".~剦)���]�A{��Y��yW������XB��[s�zr�)�% #�H���
%2c0"d����X'6@�際rck�#c쪰.�-)��ߺk`&,q#Q�8�]�}i/p���<���h�ܺ%��I����|;J�p�~#Ҳ����ԙ�����QO-&o�;q��D��&;��V����VcF
�)�9�d�뛄��!f.�7�
_�P�<����{p6�P�!����j��7H�+6*����*J��!k�1���|�3T��y>v�{��niھµ=36#b�����,���Un���1�Z`jA�	����(�ƚ�z���9pO/��Ӡ��0�o�n���͎�6�l�j����ղH���7����.�*%�_����ANx��O�!r(N����Q�Cڲ-�aF@FR�g/���
�S�;�|�� s� � 1������3��ԕ���SD���\'G�]GԌIOy^FR���Ű�4Y��YzV����)�ľ��%݇��7�YE'r&����$��Q��S�����O(�J׫�����G
���1᭺���E�U�� �#��<`�E��4��\���k_�x�B_&h�A#��a�Na�9��S�P�@��dD3c1���e�a7�d(�8rx��R�udڍ��*J|�|��%��@�f��KC}g��P��Hm>Qn�ƴh�R�������6��:]?�I8�`�VW��HK���M_1|��C��~:<�Q�&t|UuE�XP�/�����Ҳ^~�'O�+k��R?�0FS�����\9"�!7{� ?l�+��PE&��=�,�	�E������E���.@��3	��?TL�(�3E�gj��o/H�(�a�/�i��z���3#B��Z7�S��B�W�!�s����"�fY.�gI��>D��p�݇�k�����F9�tw��c�#G19�k�*��>d+sN�x�GC��ԇ��X�qɞ!&�Z���� �0�V����h�ZlW�����R_���@�`<�5�e&2;<E����zZ���LS��Z/N��1G�&$k���>���%}7gf���XI:�1MЈ`L��S/@p��
P,��
�@�����@Q�稤衉�V��;h��rcr���[d<��/��ⓦ?0�7���ߠ���l��O)������V����U4ٳ�f���0�5�{��������(�FFt����b�T�G\W��yj�
��M���T����I�_���1j��8}ߞ�z��sƆ�a������{nֱM�������o�L�hվx���>�/�(�A�IS$�I`����a��E��	�������C4�XS�C��j��wk] \�]�"�0�ɑ��F7��(�c��-�Cm�T���jTgha���G*�M͟�%"�в�cM��_mIw�H�R�g-mr��@��my$.��ڂ��S��� `D��,B��"���ܑr�d���=,�S�¶Е{d��}���ު��!� �Q%�[wz��=�>����u�~���Z�P���T���~K	?��$�s����U����0 �bY������$9FPx��.!��n+�1*Ƅ<c�eN�H�hH�)��04ə��o��ct����{o֊�ax�L����$�f%��0�M�����iZ�Ҿ�]3��1Ie/���l��~5����;S3�=Rc36�*�v�7�(<�Xʼ8�Mb��#�$N��)�-�B�9

z�c"�$�W�,�6�a<�&c_��K�h ��C��;���nX|B>������#�O��"�J )���/.�rv�2uT4��oc��H���٢ǀ��8��r�,�y���[4i	�rx��GԾR����w�B�[�5W�	%�x����dzE�>E��;\�)ܽw�Z$�G	ҵ�W�Ī������A���d�v:�g��/�p��_���W ��z���v�@��'��#�����^�!��z�'�"̂��ky�ذ���aLU]�Tk9"� �V<e�5z��K(0 �?Bt8!����<�:f��;;��Ճcļ@��/�O�G��ҴSˎJ#{<D�5�籪�ċ%O��Lw��+;���p��T?���Uky(4@�r��v��x!�;��,�t���#���1�HI��U�s��c����&�ĵx5�T�	T�Vu¢)��յ��K\�j5E0>0A��u"��U����T#g�L�+['Y��/�&}�6a���#gu�K�o|����_�>�t�1�׺�/�m��եF�m�N�3*m���\P��Af�儜�>�KMgX�1RJR����7�&Wd���C}VK�X��&�/`	���X0_^��s���{��9g3�V���h"^�'^q�l���v~}U��R����j�}���#-����Oy(p��j���{��V���
/n�N�JK`�~*	N%���m��_)����E��N]N�u�%9B�*�f������h��Z���H-�sSY��s?eP����/>�YwB��|�8��B��;@��Xy��:4��:�I(O�:i��?\�4�hȕ^�-���:��y��nZ�h��R�h��Fl�5"�Ɏ�̝S����NVBϬ<^\B�^�J1�N�@���V�����W���;�����ᣂS�J@}�S�|U���Av��	J3�x�JC^�"b�������ʑ"���Pr�T'��Q�@=�v�S�KJ�2� �=�:�X����Ϧ�P�� �J�^�]R![��^�"CN�2qmA%��)%s2䊠Nł`-�	��#���ZXl�XJ�Ӓ
�6�=��^8�r���q&Ou�8Ѐ�Ui��׉�ь����]��Ʀ�iK�M��%c�t^�i{j���8�z1��d*vې��k0�m���}��q����ݐOiH�rA#(��I�<w�Ɋ��7}NX�S�x���E�����/Q0
�$��Hg��]ɱ6�T�_�f�����͐b���
��pH(Cn��+ �@�hH���^�s�H�7��G��'�� �c�r�8y)��ם�#I�G(�|=G%S����{jE� tG��N���:#w��c�w�>*+���P���P?fy�C���K�j}�~__A��Jǝq�cTMTس>v�b����r3)�lH7Ęo#T@�{1���h�%�Lj�m�-���O����^�B��ij�KIv��\�Rפ�ܵ{=��l�?����jhp���b�bP���a,����4YV�?����Q��ŀԚ��'-�W��Ic/-��	��6k|�mi]kF6c8��~c>���`0׌��.�cpr�!��t@EѼ���`�(����t�~1�˺�ɗ.x��+��׌&��KS��Y�������g��s	^@hov�E�*��
��Sr�p ͽ��Ҵ��ļU=W��Sjǧ /�����R5���a^���A���_��]d�<�]��}!�4��q����ўm>����e\���v�)�wy�]4E��'���NC���}����W�}��4zx�M!EB��y�Cw G�G��rx�jZ�ʧ�9sי̺��N�.���=�Q�������#�	�F��h���v���@f|CN`xK��#�u:�#���=�8�-��cU�#"�-f�"�'*"^�bBS�?c��-q%:}�[���:����:$�O������o��Cۿ�p������D�ysCqK6�~�"�g�]\@�[��@�Z.���	J2fW.˦t�DlO��x��E������d�R�f�l��<q���ә=�:�w�Ldk<,X.<>����r'���?e
	4uy��ɮo��6��f�����M�	ק���`=�m=w�wxR���\�ńc�@�����F�<������gK+�����bN�!P�"���oun˃��P��SJ|?�<.�ϦNG�k�e������?y�*HhR�5�Y�G&�^�TT�aP��My'3�M����6�4[H�iYg�E[,���y�5uUχ�P х�Z4S����O��13����C�H�,�'s�j����d�GJ����+l<��b*7��������;�$	/E���d�� �=ZuU��X�b�0������Y�g>,����w�ܔ3P]:�2 ��aApFlW�I�%J��L^�雕���}/������kg�7ˆ��	��&!�d��];���0K��?�"
.Ba�~�����ڈ�bېFMT%nX��Bgca=�<�h�N�0��t��JJ���$��������+�=I�\ô��c3zEK2�@xa�]f)G�8���^��^Ke E��/JRTĘ�g���\���A=��מ#�V�&�Nދp�^J�����¦��T���U�!�5���� ��Uk<�k<�W'5��^� �����l�ⴳ�-qߓ��G�4��z�[l�eB�cK��&~R���A�}��$m��`_0�8;��1nC�S�`��ؼR�V��/��r�!kHe��v��� id>��h*p����w�5��:����jc,V��-Y%&���OO7Jg��h�Y��a��@ގF�l�l?��j�.��K<���էB�֬9��$O 4���Y�BY |ew:ޢ0�}n�%�2�!wyk�,˔@������=b��Q�T)D�@QL ��2��xѾ�5��N)��pU�
np��)�m���.0naK)�8�9�:�G֎�hv�-���#�"�͹nI����L�0EX�tapi�)ެ�_�j+R���Toe-}�8��#��MD�gy?5Z�! ���h�3R[\�V��CΙ����F$�aғU�)ec������sJ�.�o�<;X�#Ӷ����У������CbX�x8�Rf������j2
\t���������^x�u��_|���~�5%���f�L�Z'�����޲�����H���|R�4')��$���Sb�G8(;Xk4wB� U��6��t��#���=�f5(�S��%T�U����
����7V��'ĭ���V�3v�k� S�j�.͵���pb;�.+$]��O���'�=���䊥Q�k��
�:i3���{���G�|����+���ٲ�͎/<2A���8Y��{��1��6��J ��z-I�w� O�U�	7��D�/�2L�e C�!�[��Tq��Q�y&�`	f_j�,[��~F�vW/�����Q�b�k�C�u@T�:z�B�TK�)�q�=sÎ�����s@�RlIX)-�-��q��V�i��3����ɟt/���lI��rLw���v�O4%仈?���$��mG����	����pm�zX<����}�).P�+c�m��av���J@L������T���^�Ek���b%�8X�ӵ�7T�(�uHv]$�����C�#~w�ԕri`ˆN��O���2��T��hjD�����A�Z.�����}�M��A�H�INEx-��B�û�~��ڕ�c����a*�"��'�L��S^^������D�肯F�����_	����5pV֧u�*�:�EZH8O���C,[Ԏ�����|I,cR���I��ⱷ��n^�Z^�
�������4hv��8`Ir>�� '�B&,B�'�W(�Bỉ	��6�VwvCy���Q����c���W����NZP�I�r��C�3rv8������lc����=��iIv$2�����qh���,U^�`"SM��c���kL3z:X���k��p�o����+-�f?���蕉���qg�HeA��lP��ΰ$��-�5͛�l�UK,�Te:�X�(o�<��2a�Q�2: c�ѿ�5I��j��f����p��ۡ�+�E�����S��v��:HA�]g�E���u��D������w?"�ު�� �[��hZ��t��9�`�؟gH;�`����@S�D�o�ȱŒ���cҿ��\�
4������^&9s�;�]����ۓ\�v���G4�f�nޗ���f$�CO���{���F�l�ʭՃD�>R�2R���kXfެRf�/WI�XaZm�V�Y�@����,��A�+c�����%��PT�$,��&�D�?�|��s`�W�/�n��'�	�3��Eѽ�I2E]��
��.'u��Q*]�IE?�ZuRѹI"��x��N��9;��Wn�D4�P��P�!�9��嶤�4���0n;���9O<�s��� l	h���}��Opew��*�V�g]tT���DA���q5�P��F����C�"G��Դ����ap�x��J̒)��B,�[��}�[��-ez�;������M��Y�N���?��T�0��ogxQ�)�P�J����ė��@L?��q�6�<��b�$�{w�ԯ6D��T$:�:��8R��Pۿ�do�sd�?Nt6���E�{���������rƇ�x&��o�����t�d/a}f�?w=1����A��I�ڋ�_>�>�f�� Xť�)[�_�]ߦ��uM3[Coá
!�E�f���T~]C?�2S�$�v�4�iP<@�xuƺ8am�]��(M�e��ضs���p`����U�emG�zR��ө@��F$6�_����N>�'ҙ?��� �C�)S{:��ͼ���#�|�H������>7�r���[3&�s���K�����]��z"Q�F�o�-��_��M�,z���.x!�7"I���y��Vd�b��W��u�g�IZV�.���l� �z&&�h�<����z����ebb����y,�e6̃ӭ�+�u2ͬي&�����R�?�=����:��:��� ��]���%�7��[C�{ZHB:��U��%A�$eg����>\%�/�iH�Z��g$�l#N/$p�u�A��	q��R{j(Q��o�#Ǧe�R�}�p�ej4@Wڰ�M�
�WW5�SU��Js�R������_ձE�Q�w�%Z�\1[:���5��_��ܓ��O���l|�O`��=焱���d���A-^/ή0�v��ɇ8N���ۯ�|7��eO������G��x9<�R�.1 �=ϊ%��c�nY�02�e ���:K�B|��ev�!�j�����cZT�$˂c��c{4�rf8X��)���'Ÿw��2�U��Я���_N#�d��?Ukn�B7Z1 �h�����y��z��1'.�u�����Ο���r?��$�q_	).rj���H8�Ϛp�F�K:�+��z[%�>Ǧ��`�JL�S ��Y<j���?u?�Zx˂	�:����(D��ݓ,�eOm�� ��iN%v��h㽆�yh%^ ">"%�V�7�'��*�2gTl�[�����E�p����~xl�v� þy��Cܱ�O\Q��Ey�w�M%U��w�4��zIdd��
� ��p[~N�7�'�m�E�E2����o�%� �O>�߰<�m�٥1J-ƅ���,���Z��XT�9�:t'�̳ز�;�_;%�w���F;FB�8�,\yxT�2`��I�4*rܣ��"�����ɬ�L�T<g�{��^	���ٰd�����x�ᡯ1��ʧBјkOt�&�PŪ��0*iZ�LZ�A�XM�]��Ŏ H���j��ɪd�Iv�.ne4C�{�QT�<��,��ݬ��gL�� »������ %��Ӊ���;�H�	�B��u����>{�B��02�4=��b@G�����H G�7("���'�1PL�%`��2��;�R�� )WC^'�����(��7w�U1ߧX8��L�]Wc���Du	poKqu�C�.k������܀8`�œF@I�g�?���귱؎pF��m٤�OK	�0��{�M� <sub��bYC��$ǹ纸n���]�Cc!"�J�vT/���3�i�vq"�6%3s^��P�uL�V��p+�_$6"�Lm�By�|_MJ�bD?5�����D�<ٛ_@��S��vRk+�0�
�TV��C�&"��u�@� r�m�� �S/6z���$l�L�}
���֛�f0�ԕ ������Cx����\s�%Ȩ��o=ۧ��s�m=<R	�Nڏ'��
Sԕ���z����C��%�s7!�)у%|��}���oYC��^��i�:ލ�'���F}O��H-�Ka�Q	'�~Yvr�3Xm�cp�b44�t�9���/Ф�a���y�pG�q~GE���*:T�;���jT��shH7-�w��E��޵^�.p�)�F������|�/�H�իt�+���B�&�굙��-@��M�(�d�P���]�� �ݿ�2l���֪D㇩����\0����J!(ĥ<�eBP@_gt9t-�0o�p�ڴ�{����Kp�:��(�f1� ���\u�X�5��n|�aJv��M#�ܝ�2N9_�ڡ�D;��0;D�o��Y�-�ͨ?��E�BATh�V�w�t�N��?-�?^�'Ν�Ќѝ��cT��%wPU�1��mV6��>�Z9�r�<����֡ ,V@�t&y�=^��n����q��.yQ���@
v@�]�`�
�ׇ}��wT��K/��l�&� 3�-ax;�N/dS�m�2\�Xg�_~���n����R}�TT|��иbW��N�%����r����Z�6��ѹA{t�0�?�D�B*�_\��v��r�����Ga�7V����u�r�۱M%��ȋh�Z�8Ĵ7� \�e�Z��)4����&*`=�MDO���wi�Bw~���W��r'Cө�E�]D�{�����c]�Ò�i���2�.��
,�L
��7����%�h:1�7����1����!�_�!�qY��g'��^+k��܋�g�\n�>�i'��^��֏�-�^��܅.��]s0���خ_�˫����Y��)R#�6��4�U�E�i�EF��R���@u,2�r(��8b��	��� ۊV��>t������:��!���B�����ܮ%� �m�@�l/�H�f��A\4�H�j���&��ԣ�-��g\Ĭ�i�op
���^%��5�Zy����g2���Zt�`��A6��NIU�P\n�ڷÀ��'�$����}������E�=|B�\��l�2W�0��U���>���Y��Hwg��B�V9RRR��H͐W���EĘ<_ ��X�{S�M�,��G.�xx6͠1�l7e����IQ��e�)9FF�zƀ������I'(�r[���".I3 B��ˣ�E�n.i
7��}rq����1���o
z��3[k�C�L }���F����Pn���y-����n�m߭�p�A@�uD�兂�h�(���N_��.-����f TEb{��F��3����²4�Lgs�e���;\�\��9\I]�ZV)} +��ė27_�  y`P	�*~`��(�7�%w��#ҏ6�?a�����?=R�TX��|�f��ō��*��K���E����4��L��'gl�1�	~����r\Ԋ�<�m���=�*���6A<��������U�{�8S �=��0�01���@�`8�cg�<Z���)�sm���1���6�+L. �#���2�/� . C �PP�fPd�`����!�+������|�|�ʽ͢���*qz�)iS-�g\��I�����a��>��<q/�{��ˣk�m�ܸ��zaF�SP����"����!�̚�]��d�svݿf��K�T/�_�7���o־'�e��u5���g_�Ͱ6 _����Z	G�����1ԑ,V����J��ŖEٙ��*^'c����x�]ZG��?��5.��ұ����{����j��.�	�s�z�6ˁ��[�1L$܇/��U����8{HB��v\�Jy{őJ�*Yk�����'̿�wQ2��c��̹�3��\����U�sF�$���*����F�u]�SR���vs	���s�.��/0:wwpq]c1����|S�0�GB���I����Z����J4�-�H�� e���� �f�ښ��L���C�Z.�j��DT1UiF����m��o�oF
H�K��Vs<�ҝ��s<�/z�
Q�����,��2������I6d�^��"c��T�����G1U����T�ilԽR����3��J;�v�~}2������ẜr���aA��яT�A%��Ǡ�͞^ľ:����Y٥�A�qi��:1�ADr�1]�s��GR3�o�N��ѽ�uVP8�U���~p��bk7T�M����@��2�.iHl\�o8���m�M��_����:�����J���G>�����p�IK�m`f����<�1o3�&N�"���NrO/U��?��=4���g��D�֨:	�ԅ��6��:���Bp�ߍB�'�g�����܏���Bi�<�A4�� "�����2�f�~�G�E�6��$+%.��ny<���k�����}?b�Ok��S�N1�U��a�Ճ�q٦da�h`y���\P�#�/Ѧ��k�P�ܑ�������񲌏��W&�0�(����a?�����k����WQ��tnӓo��}�{��m�!�	��ouUae��,B�K(F b�P��s>$��[i`��{�iҕK9_�i�P�f�]�ƪ�°'�F*��/��~�a0��/_�8�����c5�V��mb�A ������;'ۭ�����L��9�8��%�h��n���~�=}�{���&p�$=|��'_��l��ퟦ"n��G���
/g}� U.
��p�������]��bOp��;
?���ԫ_V�p���4�d[��TP����2����ܵ�,��%�*`Ks�7��S����_�5E���`��s�=SPTY�	�k�_�x����Ak���/=�m\s�Q̆A���!=tҸ#cN`�G��7�tUI.��>�|ڱ�q��\�������9f�v[��a����,��<�� �d�i>4��|�v��,��?�i�$0�����mo��:�iaӒ����Û��8��Zz,:�}	�n�>�?���L�[�,[��S�j41��^��鹔�����w��_;���4�4+^�R�:�އ@)8���= l�:�l=���}�����"�|����䅘�2�*h�Bm;�ȼ�{�Sv,������Ӆ&*����@i��ڲT��@�au�KW������wgGN�D=�Pq���;��j�ҿoC�d�qy��{�A�D2�=\x�-U�t�OB�?�GI��L���᫟R�F��ef3��eU�)֋�cz�/�$`f$��q����������Q󬝓���zI�腲d�mt�7b=����J�;��T��]�DT ��e��5Q�/����VCZg�C�/���[U3@,�$�4�F\Q�PL*�d+*wT���u�@��hҡͧ���ݜ8�BW�g�.��1ߌ��b4׀'��
��$�&�ŵ`!�GeJ
E�c���.4���f)��,�\ �:h*ԓ�7��21:�VǗV��l�7#�G|���o�<�E
s�7�tg�T�x��I�����?$ k���r��k ���J)^�x���~%S�������&uQP<�C0��"a�)����L�s�C��zN�Dh��Uo� ���=�!���]KKa���e���'>�>q�ѧ�'\*��H�k�g`�/��D\w\����bw_]+��n�����y����+�O1X�Cע������8�h��<@����>�䱥]�ߴ��h��yD!�4�&�$���6MB"�����9��x����D�~�o5(�m=K�ϻ_sk��ˁ������[�3�l����6�G���{��?�)x�础� ��_A�\B��kȱg��Rx4R�����v����ni�]���� ��ȧe�[j�	GƤn�@��z"�A�MP�f"�([���ez���и�y:�\�FC)<x��s|��F��)qZ�D!�3�]�pj�>^ l��R6�B�/V���������[q����wI�,3�]�y���P|�-������F�>��8ۡ]�^
��W�zXnj��.G�'?fn�*6�?Չ.�N�
��g�/�O���s��ԍk��/>5���8������9��Rwd$���,*K�P����._���o�}��á�iL�͋����u���Z���b���3��KsI���b	[�lWW3w�������?���a�|'P����N�33�9[d`wZ��ܖ��e�k�|���no��w��gD>-�����&f�n莣��P�ϊ�̎�O��P����.ڙ��wtm�֟|=㰃ܫ����p��3���3�Yf]Al�N�Q��F�]���6������ zv5|͊ELy_�؛��7Ua�)$
�|}8|w�C��یlV�$�~d���DL[�-���}S5F&YY^7�9�/d�O������1$�&��E���#h�J�خ�i\���!�L� H!>��� �!{�����t�O�� �b�уL���T����p����VA�n��'���M��,8����a�ܞ��N=
���D�͕+D�PT�LɊ>e��/��~�;
��ҡ+P���Z�G-Y�n�13&D��*[jh�R�� ��t���{�*y��r�x�K�n)�~�K�u��
V*�^j�e��[�d�G�S�����XQ����5x�� ��a��m���߃n�U��o����9G����X�؃��IT����R�.m�*��Kw���T޸�Ep�;;J3-XwoAN9F"y�22l�c�t�'�U��3i��M�fk�0���~��ǮdxR�}ǠJ&c+�����=�&�f�]�E\b�f�[n9v�U���-$GZ$�11�许��L�����c|(2���k�D�
����5�i����C�����n��K��tհJt��)\LΣ���ەX�	��4��<�U�3��zNw���ı������F��	����er:%j���}����c�0�!w�?�����bc�V����
�t�"�l���l�-,�3X�z�J���/������j����)jS�<�[�q��I"�
*x�7�@V��|�I�B����B���� �0ݷ�d��L�풙`���8�)�7Ӕ�\R���0P*f�u \��),���d��:�@��b�T"������POC	cĘCò�� ���,2���0��3�s�������2>�h�D���|�͙q����BA��w�w?�q��Tg>˃ί�����8��$u��eI�>��q�����̛��d%-����^�B��r�X݊^e1v�eS��c�������0�R�:ç��B'��l�z�2c'�F��e��C��F�(|���d�Ə�?SW��&�؋�ÖIO[}~�{Ov���oq�����[��VwgOv\;]~����?�Ӛs�P�T�_�A9.,�:��}��٠r��ݷ��ŌN��`����� �F�tv�1w�145��n,{���Ŕf�R����?K� Q����`^�����5p��
��rk�ȗF!LO��O�����/$�\^yW��f�G�SaL��D !���z�Q��r)$mܖ=�?���_Y��GiO~���;�����cN-��
N��8�S��5����!*xc���.	e4�2�؄��ךb�$F��c%����iG�SKr2�P�����o��,��ݡ�YV�"�#F�B���Z��*|L~`�<�"�bp�ts��c�f�G���BBM��/X�с�u Qz�/�����}gY�xV���;��r�wh%\B�a��*������O��<on��?�S��`kv����^B�VB�0���
_�mN���k����"�sv�<	O��ە���d����u@�3!D)>T���I��rV��8��-�7`���=���6���?�$���ѵ8��P�[�J�K��n���x,�!�?Ʌ��a��3+�e�N���cГ�)�ƌ<az��{���^���}���%�A��
f�,���ӆ����2�QgA���x�!ls�zT  H�4}�t.�Wz߉(;;S�ǃ�>�d�����_$`����*����Q�~�K�~�Y�nrqp�8L�dd���8y��y�8�{ .2]� ��͉NV9_t���[��K^�Avy�l��y�$� s�v���!�Nt� ��Ab���)�c>[t�~���1f�7T`� 2ܓ�PŖOl�X�E~]}�)�*�z^I@0"���-�op��a�x	1��9o3�7_?��Lt�+����"��E��*�?D	
��7��F5{�i���,�M~(�B��@�G�? �s}ҋ����;�gTU��k?���]���~\�Y�,�On�EX�T��B�ɓ1����@l�p�=�(ɫ `�4�w�&S4�6PV�~K�q�.�i8������X�5c��0P��Z�X`§�S��x�$7�.w5�2ѩ����.F3��|K q���/���'��Ԝv?,ܴ�0p�쳇q~[��҂�Ա��Ð>��lN�)םo
N�'+�,�}=����y�䔡4�@C�"H��˝]I�.�F��{����5�4�q�� ̖D�|������:�����BҘՑ)@��3���	����x�t�[!���|d�cӣ���
2/����Q�`�H�=ev��W�n��]�[�H0�nj%�t:0YjnC�^=/]\���Vl1�rP�nL��}��TD�(I�*��,��$x�E���Σ�G�=�<3���\^p[d��
ܵa��3�Ө��`F���P���<�л�����NQ˵FOE=AG{��n����*�Z�=��k{����ٲ"��C�֬[�Xb �q�y�b0`���T��?��
Oo�|i�Ծ��BF)Ζ����{�|~H� ۘ0�����̴t�u�{mڴ)�QcdG��	����������qQ蠴sJ*Dux8o~+0�0a��Ew���C�Q���Ҭ�(�v9�sNw�O�;��y���V�rmd�/Q��
v���,�@�"�0���1����~Z��<��0n�_פ��d:�
���q��3��BDj����@�.�F6^`%��}!)�>"&oJ��:�J��X�T��a�.�F�ݼ�����s�8T��S$70�Y4��Zc%(U���%<hͰ���"����&��dx�_�QeE�1h�KIz���(��5���k\~*�3{���qea�oW�%zO����:��"?ݪ����.,y��F�.7���ǩHh�h��U���٭��F�/<7K�DE*�(Aҙ��v�lI�B ����P�r��o�w����g��C�Yk�Mx�]L�+jT�&ea��@WT��@�EE�9=^]i�ݖ�}�/��3�>S\!�_��CR��AA^��/8v?�������L��'��␊����ٷ���j��?:�u���v�ſ{���7XS���{���;w�?a�8zo<��l-�V��Ru��2�hXS�c������Rݭ�_ ����2�xt��HGa��`b��?q���ILԩ'坸�}��x��s#`D�g�?Q4���Z���PsE�.P�	p�о�rq\J����~��#sui����\����>��	��a��l����d�7쬄ҥWw�Ðm�2�u���g:��g�2�(=v�>e9]�����G�EZ��<_��YFFMmTh���q�"\�����*Z��9�ϙ�V����i"�����"�}��8 �gi�F���Q�x������U�!]W&pz�n�vV�������n���!��/>��Ơر��k�?�Zo{{����ۙ#��˂�y��oyæV�ٱ��I��S?Y���������EI�#����I�;�������Ǣ�ܥ �Qe�ϖ�����:,�N�����H����Dħг["z��H	��תd��q9���̏�F#N�	�p�����IM/\"K̵���?%�~Д�E���$���f.����w>n�bp�K�:�(Q�{(��/���1�!1-�9�W�"c���L���O1?@V�(t�Aq\���K�:O2#6��6�bp�����f�BP�F�����;���1��������`�>"ב�i��E��dc�&I�/@�/�!�6%�=�ϼ���L��pO�&�����NM����w��ҫ1���2o;�Enc��Y���Ը�!��o�g�')�ɦ�%$�]�뫔rGrsZ���$�o��8)�OK�S���*�Y�#��v	n'}�JF�n~�5A�\-Rb��sU��y	�� �������Y����zrŞ�5�����Ҟ?ԧxt�� �������9R����%�?��<�,#Ip~,́� �!��p+:A3$����.7%�<��Y�%��ʱ!�t�L��PmS}?F*�/����g!J��7��)d��M��T9.�T�$i&BC'^��4���<i�#x��$��$,㍶B�����㍼�R�� ��_٠���ݾ�uĉ�uSFF�~'�E�h��;w;.�,�ˡZ^4��f��87�L�Hok?*�K����4�Q�H��kQ��Zof��E����ț�h���_�w^�Sm�[�O����ͺ�=�@(�u7�';�(%_�ha�u�M�},�6 ��"�KrgL�|�݇�v�S�)��o�H���7�[�f�{�Y����_*� 6m{�H N��FR��)[g��W�)$@�M}g�i�aeXż���C�E�[�q��|�;��lk��/�o|��n�D�N��ğ[��5E��\�j���a"tFF$h�U���HJ�Y�b^��fw�sY��_ ���u��y��՟����kF=֨"&v���V��;hYin�V����hP�Zyu�d"zb�s����O��̱Չ������b�\aĐg޸��s��(��L��2��a|�1U<���5��&�t��G�,Y�А>�4����yO�~6�0�Ck���&S;r�T��F��q�[�.�]NڠeE�.�b-m�]�P��ꇲ����6���8�Uq���s�SV�G6߫`3�U܏s�=��Ǣq�?�]R&}T����I-R ����i���p�פ3�4T�Yr�������I5D_��QXB��0��@A�gǺ�������99R#�s��l#)�Y~�Cj޺�BR�+�BR�`����R �r�������Ã~ Wo�8� Ã��łrI�v'Dgx�B�A�"�S,��y-�؉�k]��>��vR��pn�LL�yw���R��#F�	��J>Y�Bό����`�/VER�.?��kl=��Z>8۵¶s�n��R]�)$�x@&���`��\q�9��k �wj��uɊi4�Vh{xؖ�\��ˤD9��G�� [n���)��4��*���8�����p#�|)�W��m���#rd��HeK(���%�th} 
s��ؘ'yW�x7}���,���2�9 c-.us�������q�"��'a<���8�hv��Ȇ�C�
OI�bZ˶2DF�* f�^5|)�>Ե�j���D]$�Q_
_�?�خ��c�-���+u��߀�B����Ґݮ��؁ڎ�����n�w	��qF��+-$��\�+�JsE�I|�h(����;0�hCz�rE2s#K���sS�]7m��t��b�u��	m��(4~���+w�2Mf�.y��4kh��U4�[�`J�ǣ�5H�T(�-���៓�X��Ь�2Z��}iL��Cw�h^{;���I-��eh*}������v����GK��&�<�Q]�w'`���k�>�d�#ɇ�p{���DO��I�r��,-jyșo�z�(�E�]1cp+t��W�17���rM1CL�5G�r%��_RG�5��;*����R�λū�@���� � Q�L����>�@��6��3#�V%D�U���_�F��
��;�WR�A�̜�Jz,��ث����bO�8�I'V���k��ɡcЪM���ǔ��uL %��n�Ɯ$A�k���ߢ��$���G��>��v��WA�!A��j/�agi�шR�l�+���5�]g��^�u"<Ho��v��2;ffJ�D_^������}���6A�BQ^��1J�1`�a��a�8u>�5
H`�6c!Ti,�$+{�)~�h������fA*�P��G��b*Ě��u��`s�q/@�5H`�t��#VVϾ̚���id��w�0U�[|T<ZC��)Z����>�M[-�vP��0C�/r���
8;�ƛ=f83lg
��ۙO�[ѡ�B
2�:�,
%8㵔�B@LN4>�p�_���6�Fl�b��}+��'G���0X��k�d��a
��:�u�mc���K��Ȃ�G�mv�����~��ΗwmyX�dy�G>L1h��M<�?�7����̕��(��̞��z���� ��Ă[�B{�7�t0�	&��������Č.Ֆ],�[�XJ%�R�S����\�S�����c,Z� m�Qo�\%��T�:&K�F��"X!>'T`I?=Ɯ�`����l7'mE~)i"m,.S�+�h����^�p���.#�+�1U��5���Ai'�I����/��m©��:���/h�I�P��L��;,g��� ��=-yu�2��,���ꪌð�g��i��Q�_}A��$x0EOG��ۈG�K��jqf�[���#:#Is�01�0aHB�C��¶C�p\�UY�Mr.�f�;�+������{it�ΑR������|ʳ���	c�8�ť�s�G��(�JB2���Պ��5~I�v��P:(���U}�R�/K�,/��ߵ�{�W�!�hl�J��X5�溽�f�G�
���ܗh	�7&-��$__:��ݗ>�3�1b/��.�m���E����p�N�]�=y�hGt^�F*�N��߷�	U�d���2�?�Y�����s���L��I�K�/g�w-�egf*"?���+�[J����G��?j|���Ð��������2f��ڌ�������&�E �;�^g����F�V��v`�r}]�IP�3�RAͩ#�K!V�g�@�/Ρ�5��j��{���>�+�b�YYzX6��������^#��<�Dd)�d��v+�t�ͅ������*�.��k�����2��i��`�����)�ۆZI���"�_��8���oɎ�FR�+�n���c�n��Dx�aٔ���æ>;�{�����LK�O]m�ȅY���u1���f(�Pc��b0NX ��� �M���s�8�����xpt��i�i�$���9|Ì-2*z ����UٓH�͗Zx!�s������#�U{��8�,�ʺۈ�Rq�!�Q�N�z��P�G� nz��8�4���X��:�\��~�k�S��O ;���v0J�0�ͅι�O��1��ǥ��h�;���Ȳ7'�ݓ�!ü�K�;-�S�2>M�)F�?\��տ��C�y����p����l���[��΁55�����A�2�(q����W�9�C��h�B�[�z@��i����&�����{����WԽ浛�:]�mF~d�MpKÿ��֣b�2>�
r�!��*߱�!�߸�U����ʶ�˸@��hU�:�c�O��u�i�1b�;�PQ�A4��{|x��*��|*T�^��'J̬��J'��L q"���ʼ?)Ny[���IN��ρ}I���.�dJe+%����C�$Û_�8ɠ���$��\;ƞu�RP@?,��7
����`Kt��|�� 6c���ԔvmSڼ��C�Ph~V�؎���I��h�ڌr�cyp�D����#U��o�<96o��$�.|�`T ���QSc22��$l�P�>ܞF����v�`'	����n5����b�(���w�}?��5T#N>Iu�����ɓ�$��8�R�&�dMkr�z��Ti�w����>��~q����f��7��%}�ĝl�6\��
��g���z�6b�I��<[���T�E�t�
��X�Ç�(d/QJ���H�SSEU^a,�̮m&;+'���*7�jN���:��@�eanRԠ4��s�q����$!�4⨨���N�j"�y��UՄ8�F�ɳ��{0�~r�&�3KlG���f�՚B&<�	��Z7V܂Dϵ���0Mx;ft|���]o�P���<L�I3�.?��u�{]���t��&s� �*>��E���oDw������������B�6�+V�T"��z�Ua����W4r}kߊC�R�>N��*b"�PkO���������|7V�t�i,�2�Zm]�f+��	�TW���S��v3�t讂�W���@��Q���|?3��]��o�Y���!؎��9ڼ��m�N�	����o��.��R�3�WT6ϹmQA==3J[2j ~&{-�e���[�@Z��&�B/�X34���|�M���&	q�A�K���v
����Q=&nS{���$Y52�(l�p`
�I�>$DӔ?�,�O�_	]� �i��k6Lp���|Ɏ�
	*�B-M��V��� g��@�b2v=�zw�����!�8hhH(][�:�4��K��S����Ԕ�%�>���cj��F��\So�|����,:�)�J�N|Z�ט���n-Ԑ�`8��*tApq��j���dt�)��ǀ��I�J��$"*��	Å������=r�<;�,�s�@�#8`�!?9a6��qR���L��h�.��uu�m*��k;�;�_�֏\qd�3��j�������~U��c�]{�� ���+m�3�JV '�[�ϴ8@9�������j�L�>��m_v��JY�1c�nH��o�'V�b���!�㙷���
�_y:ً��,�q���MB�e>ވfO$؟y���%48p"LH�(.��|>�G��r~ձ��>������z���<e���Y�T{ڒE�dfDW~!d�S��O�C3���>�Hz���LW�ڰ�?K	�ZsK2�4)�)�I�~��Ä�{�{=׼�~���z
���<�U�0��^5�}��v<S�W����L�~�ב�E��'��V ���AۜXW�meA"��LZ<��?�x]�=:_QQ �l����eI�n�7*z ���E�i5��߮ٚ�4� ;h��W0�+�%H'��n9��F"Ц�\48]�,HD�#������Ւ�'8�a]�C�/V��A���,4,$)�:L�B$��^7z�/��JA�V8p�O�5��G6^d��@�/�4l+�5�:4�p�����'S�s����F��`�ܟT�#5g��2�T�.{�jB���L_/�6�t��4�F�oZ�kI������r����.E��>2���Ԃ-�z��ù�'�B���a�I)�#�K/�R���n����s�4G^W�#q���n��8fh
E��A
>��b�=�Ӑ�X�L�8���CЮS$N͐h6�&W�ĥ��­�I�B�d���M1������&�2���,`᧝�E�y���L�{�A�Y��۠IFo&����,�9>��{�^hj���q���oHF� ����緹G�h���[�r�<���!cQ�Ħ��J.�3GIx�6:Q���%�w�p���`��8�
f�p��)�U������0�O������X���Ң؀/0�pEd���)��}#	�����x�T�F�}���Xr��������R}O�D����*�Y�nK�''Rz{���8���z>ΣoS�r�;]~���u}Ɵk�&�B^˴h��}��%u����H�}X��HQ��e�]�����%�B�r��sY?��&���d &�.,!��GD@4��7��G9�}`I���th7�R;Z�͛첓�
����O[/c�F�+ٗ��T ��\�)��xB�>'��X	���8����<��'sDf����(�IuY�Ds��w������G�eK����5�Z!�����_xDO�]�jcpE43������~�E��姳�9�����7���eE%�ٍ+��6�Ei�k�v��N�%��#O w��5�,�/W�U��]H;8�}�U´:T�F�p����}�m�����ԷF20�Ɉ$��P��u��8 ���m���PT�E�bܔJ�3���ǸqgzCI�_D+�3���,����ac����β,2��-�`���(�SN�S�#� �5��a�
a�z=˰�%nv)�]���n,P�/��$!���J�y�u�XF]��t�U^�\6iyk�X�B4�/+=�����Bl0j�~8� �����.aSx�,ܬ&�|7����p��
��w\:�ޕ��}_��e�"����߂�[.�M���o�uj��Qb��a�jb^�W��X�lG,y���^��C=���|�w̃��������4O»!c�|U�;Z5������T���0��	&ɴ����`OF�nk�P1�VS%���ލu�mk�Cڡ_	N������B�EE��S���Gm@T�楓@� �����k\w+��d�T5U
����-��^4I�%"��;���f�h�K�xĢ�:ֳ}��*���b2���'(p�gK�Q�.V�(�*&����"�8���W�䯎�o���JH�tvi�!�A��>�á�gV�-;�H#٨�!���/5D����������='���5��m#�R\K<GD�)d������Z�ɮǥ4!�8(����u�L)�h�� �|���� �OJ(iMlc��X;���~�P�̯�m	�����3r�zI�o��7��ѡF��4.k�޽�����PxjTEܸ_��Y��N���D����j����˒���M��V���-ӿLBGrV/�}�	�
�V)S�N\ʽ�70T�H#�B�$Y*c��me7�� ���%�D�nK̽X`����X�'	�������f/7��4�Ə���4�c�����!,��V8ݙ$N*�N|�-{U�sq~�jh�V2�`ܚ �e�/�pq�l��P�3,�8�LʰKέg��c������Nk��W9�G/�
�GNh%ӊw�����Ө4<���+X9��cf����]:�T�X�0�yp~��~r�j����]`�5��K����n-x���*����1��<��<DA��#��P�,��|��ǉ���<���9Zr���� �g60�^4��dl���p���%KE+��J�M������h�K&1��G��L�0'��}ʤ$�E� ����pO�V��|���M?gd��v�w�,Bu��$���1g?M��pp�N��&�C�z��/��:�z��ߌ�8G���2��]��l�P>��܎�%�=�[�����D��nټ�Ke{��S�K�p�'�F?&�7��Z�+�Jg�����߆,�14Q�Gj�
$%���(*Ⓗ7� ���N<���,⼪;A�O7��\�y?Cބ�w�T�Ф,�ԝ���
S����?{ɥ\�j��@%�f���?lǵ	@��{NL-:<\�3�Yr �����رX�����M�]��^��⼂v�­k�)v�_��?歔����sA���Jƕ�E��~(Ŀ��r��s𿰙����,
�P ���zr7�Z�W�K9/@  �P�Fѿ4,�Ӣ�I�W�b�I�*�ynOdɛh���i�$��n�?��4���`@�[^����!�`xDyȫ�U����r�.ٻXJM�bW;�%MJ����:�=;�6ݖ�5i��53�8�"˵�G������*�ʕt��/m%��8Pof�=��-K��O��2��3l��2"o��񼣓�(/=���ċ�'Sb�"2QK���4���56J�\G�2��Dt��|�Җ��r!'������xv��-d�̜���A��/rTZ.�D��Λ�{l�2�����]3q��?l�5�.o��d��q����{m^�{���~�w�ʄ�R^��|�c���yY�5�`,�+�/>P�Ay�7��m���}ؼ�\�2=�.����	տ�;a�G��v��k�e/�&+���$�j	��?ƙ�Ȉo:�&.�t��JA�i:�{���p��s>�F#ߏ{��o=�_E,��<�S+Vuz ���`��{x �*�b�ڧ�X�[�S1�i�/ �?�ʅ0�bI��R7�/�xzL]&zQ�M���G�w	���9j���6���" ξ\�'���q=�2����K�Qpm�2;Ah��j
�IDHut�)��C���^=߼���AY��{j_R<��u�|T=�ئ��F�t��A��`�D��?��z��1�uV,+����B��b�әb`T���A��c�S�2�׋����<<Eԓ�磔���0E	n����T�)�a7P��f���Bx�'�ܹ�����Jd�S�區�N��VU遖_���P�rV�����0t�`�z�o�d
�t�XØKqi����Am�{�:x�F���'̾$+o{iry��4R&��e����F1+Ps
�:Vz8��II��%�A%��2�����#��F���2o����=���RT���E��Ci������?����=��.A
g�B�1���]��S����=f8T�5���D���A���l{#RKcd1o�w���%X���j�M��O�ݛv�f�,V�|�CL��uB!�fԜ�a����D�]�R7d��^�|iƫg����U�ք�t[3��R豆�Qܷ�;���ƁP�/$.|�$H~�쵽�5�
"��z��Ki��Lg-đ�}2,�w��-h���mD�6�c�c��Y2�#_V��|�ɶ���(]ДZΏ【����߲l�e�y,D�)%=��3�����4�3���K8�w�%� *�?�����K��K��`�uV=L���2K���{����xU
�+5v�զ�4'T]Sd^���������/B<������g8���۵�f�yS�¢��wo�[v#�5��U=�tzO��	4�S�É	��}�6��v�~�C�>N^�P�?	�$mB'
�:���|_�*�����8�&��s�G�(�K#,\Ԑ�?�6�ѣ�Ԛ`�n���Y(:�8�����f6b<[��\p:���o
򚻵N+j�Bo���}H�}W�����rԬV)���q�3n�o,P���<���xIF�!��r���ۋ��x��)����I<Q2O�ae��8��e�@ͣ�1z��:-��f�Q
a�t�ú���]���G�6�Ly�TG��������ӈ\��l�l~��.i'R2$�=����\�x��ď3�"K�a}���qg������ʦu����2g�&���J���P���C5�:�Je{�kEi� #�986J\>8��Jh�
� ��=�8���D\��#o�w��hpk��
6�]�bď�Y\��:ͤ0�Z=e��I�M�H�+�����'��`��s���*%�-�%fX���F����Q�\A�ǚ`ZX,��8H��hͳ�_�HcI�
q�#񎆏�X�� j�*���J�r����;~0\sďkj������Tp��b�qF~�t��'��Гv^i��z��MӶe4��@�4~����혇=�����A�2<����J��_�&�T�\U�W��#�*����H�~��/����P���x�i)rY���&i��1�M��#B,�H��+�e�/A�2^��p2b0cH��O�E���W�a��ba�16�w�L�vP���y�rK���ds��<�u��p�[7�l�����a��0�ǟ6��&%.O�:��i�t�r���x��|CU�ޱ�:�S��5fov��$��q3��{�H��S�݋��N���L�⅚�.��3G���=�7;is:�s��d=�|oN���-_��匆�l��hx�^2��{OS��/T����ksK(��B/�J�P�ݭVhO;rcF~�٩���F�y�Ŕ��Qm��_���g��@��#`3��[$W��IE����;��=sɇf��ߥ�nF�^����ɀؐ���;J��`q"_P����<{������(QUrL2�k-x���;���҆����4�:B6I�LBg�E3�0�Ư�bpZ�!+��}����e���G��r��7�dO��Vu�5DjQ���D�`�������I�D��+=ٿ�� $X�_�!"R�cnNB�q��� ��`8��D�;:�o�{��U7G#o���bUI���BZ-Q�r�.C�o
:��)(`�@�tɌ��� ��w\`��oYb� ّ�i,�t��ql�$�u����Ӓ�c/�ެ]��9�X�����_�P��T�.�w���3pM_�!��ǻ����P3�ƚP��	�'sx��;"v����I�-F�p�)�`Ǒ�M����#֢Ns��|ԡ�1�ܹz�KE:.�F}w�Ǳ&u��y�Z��:5�#��������e!�jp<l��ʖ�*�gP�<q�e9`[e��h\-����8�"��?����$��'�k����W����z6�?�%&A�:�s�����ʛ����9xǹ�Z|���>��\�%<���%��3ڥ����(."�IGU^b�";Ox�j��0d����~����=�BY�a9;幤?L�d�#��u���(�~n��2�4��/�����Սϰ�I�f46�����i�{gS�Re�s�,��Y((�O�L!��56�l4�X@W�\V�f�7��B�q����\,�M#`�7N�U���渿�r����@8�ƞ�
E]��+D���Ă�³�:V�����.Bถ�oH#u��!��RZKq��Ow��j�%=mr0���X��.��+}8CF�Z-X���Ԝ(�q��x
n,���XN˪QG�F�lL�̮���8T[g>���=ု�И*Jj���Ui0'��F+�nh���LOM[�%�s��a����H�7>Z!,�R���ß�_̅0_D�2+?��g{��Y���xm��N�0�+ؔ
yB�d%#\��������A11$n�	?C�!j0�	�ާ#�w1|Y���}蟣�
������?���Ak�=d7��?}��~�PtA~�"��>e*0�\ N�� ��lT+[��V*��bve�i״v�k��CU!v���+��� <�c{kK��q}X�)�'ۆ9X�#^�)̬�z�P���\�P�IC<�C:��_Z�OK��IX#�)���q��%Gb��wF,
KMM~�随_��AI�9�h~k�'���IMM��QiO��=���F�[�q}���7��qeG�4���|�s�ܰx;��ҳz_8���t��l)�-7Rnŗ'���a����N��荱v{c���"��M|���&`�N�{m?l��jQ�����aa�(��.�$j�Y�A�1(�||G����)%G��9�?�������5� �p�R n?�n���SNFz�+]����.��蹚������;�ɰt��G��M֍�M#^�C�d�����+���#?>�vg���" li��t[��.���e
Af���_��d��Z�8�.��P�}��z�;�R�},���g|��-l�}Ҏ���$�"�S�+�'c4�/+�WtԜ7��~5�F�Y���Z�%hf��&�ħ^�����씒h`;
�y�!�l%@�Ǉ� ƴ��Sna�4�J.1ЌM�.�g���,�@n���U��o��Uoh�2����z���HQi�{�-ez�L\5HM�ɸ�N��ƾz=ݍ݉�M��w�8ς(��m;�cx�X`�vmR�s��g�٭2�Z�%�:����bƄm�i�th!����Y*�)�"9?�*���h&��bP�1���2�z������$q:���s�<�2z�
���b�� ڃ�Z6��Q)�e�ߑ�Σ�a��� o���b�"D����I\��]���iJ����19���&�r�ڮۼ2��

������rof��@C)t'��$]��ȓ�@��CJ��b�W+_e�)7�/�ٲn�-Մl�?���d{`:A؝�;��j��ˠ}�`N��y)��HSf��� gw-B�kaId�+�Du�,'���+W�����B�>J�&���G4Dq����@�ׁ&�P�-M�E�2��*��&���֔\ll�l/E�n0>�il'q�"ΏxAx�~;�4RR�jgP܏F+��~��hf�z�o��|�n%x�p⑘n�3u�}�ULs�`ןW��Q)܌��&��v/��Qa��%�<rxX��=<[���+�}C�f��ƨ�H���ڇрu���������d�����N��@j�? t���]�sv�nk���#����Ѹ!?n����������n�k��.��1%��JcY��u��J~�܇�gd	xJD�L�~v���+��*�R�j�6]�xԄ8>@�.@@Ў��Y�����t�6�]��ܹzO��>q�9�Ld����.GR�jnDgF����zp>|��:{F�`��ݗ�t��	C��#F"
x�C�eX��s�*<����z���*�D�r��<%.�G�(H�B���	Vz��� l�=~�_��9T�6u"B,e?q��k�� q�̕o��|a�͸����K̐i����׾H��.��p>�+F��󏞝�B��0���������ʖ��U_t��J�\,�����x���a,G&���$�{&^S�˃��2|�eNx����T��L�{��YT���K�3�?�P?)�iˮa5��<Z�il�-g��>�&?*�M�+%+g�xm*@���З���)�\��;FDz%WuDRT� ���?�� Ec�������h�
��n:�,0�{J�`^���B�#��<n@�X5]�Kw/(8�L޽��}
��X:wn}t�M����a��"�*5�U&��n�g��s/�ub~�)s���$�j4m�Ԧ}�Rז�L�Z�l��(��C�J+ZQG�H5�qѹ�0����`�<>��JzQi�1�N�@D�����_D�?��-�n����y� 3�/P���C�R����u=��O��K]��Z��|^��Jmo=(����	�;tW���la�Gx���36D�%{��I���:��z�졥y���t�3/Q�(�.u=!�d�!�H�,{���|5Z�
c-Za�����o�%��b�;rn�)�si��^V�QS�Q_y�d�K���P��V���|s��-�*�����tG��8Z�B����0�7#憴���N��bL,8�tO|��f$*���3AS��;��O���LB�/��]H��:��c����R�ƫ��IW��ʝ|���n;��1�Ϻ��&6V���J=��:N�K���wzd���-:aI&~YKh�bg<��|�-C�h�����T'��P��7Q/��߀�����(�ՊU���xR��ĕ4�Z�z���YnpM^�b��j�<x��Z�꬝�hg���w'ԵW����	��֍���V�I(�6��Ĵ[�v�Q��k��'����}�L
^�r����ϋ �"?���~`�>��qR�ch�r�E=�i���.�U���� ��fR� �����7�$C+d�O'N��/g.�����[d��P�m���4=�4�_t�8�������,j{��[���������Q�~'ҁn`l%C�c��%>TS%��P,�Y?����c"4����Ӣ4���_��us�⋒d�a� s�K8iN�h:'$S��Qz�l� Pv��Z�!L��j�2��`����<���i��A�a�A����&� ѿ�(�g�'�+[�,$y�!�*�[}�c�pt�q#R9����$|/Q6~��[�ȶ'���3�]���Psr����O}cJ:c��h$��>�����|m�8ŅՇ�B��*�y��3�<��`��t���IG&E���}9��Q=MaC�x�M��#�OȋHL���{4)�e�=x4t4Wv�'v(<|��b�h�,Oݓ�Ĕ����Y/��O
��/���y����n���l�mk�K�A;�7��P��t*��0�Xk�������^�\��c�> h�����6.%�I�( T6o�p+�T���vD� Y�]c
ɪ�v��*%A�&�,�Y�
��]*8�不���-p�lɌ#߲>����b���������YD)��rZo�WhP������]�|frD�#�f�HO�hk5�VP+�d�����D��:�oG�+�iXBl;�k���J���r0D\�V�����h��kF��:;�cU�������/���V���t��Ǖ����S�Z͐�A�g�#�~:,u��cɐS9��<�#1���1z���k����Y��[7��Ԭ���,�X���zef=�ݩ���e�f,�eXD�Dg%�����t�\���g`. p�J�I�.��6g=d/�BFY�����9$,?��`T�M6XAs1���K? �0��(3�,|�)���!�1�Z7�
�+�[�~�9WR�t�u5$��&�{ә�ĕ�d.Q$tّ�ق�p���������Y��&1>�4��u��c�Ai�|��JVE���Z�M<GF`#s��xX�O�K�ʿ�Fŉ4˶U�JsA�Λ�`��h��K�u�I�̛~z
�<�Hb����Y�� S�H�v���KP-׉:u�=��� ֡![ҙ�	,���C�i���A!���82�Hb�;�$Љ�S�b,���犉��r4�]f/^v�hs���X�P%N���
�n/hFP�*?��](���-�n�S`�n�5��<��Ο�"���M�e'w�mP���Lo
�G�F����0�+����B�T���	V�p~��9d�8q=���0�I���̂!�tnB���8��_�i����b��%h�x7�O��H7�]��R`v�*6Ꭾ�k?�j��ƀz�s�t��5�=l_q����V�-t�$��i�mW�E΍�E�7����`��9�D/��=����G�/;C�o��v���m����ނu�w�:ev�������taS�␲���I�� w�G���+�vC�M�K��:ڊ1nmС�J%j���4�I$���@��3��Dy��R�h8�dt�0���z%��ҝ�4��E�e��,�a;, ���n��Z��[���2�\f-�A	����d���t8�z9jX�o��+K���6 ��B(�lt�z.�� y�F:l����w'-PN{2c�*���<3��0{}��a�7]7��w�� �N�#�~sZ5���P��6$0�������Z}�K��n�+��XJ@oZ���@0�,�3�x��sP��b�;VKf���1������Q�'�0jXZ�^��E;����v�FH�~��7�p3�o-=�ޯ_��@evۍ�dº�koYA�]v	��"�&���30�+S�,j`>,>Ee~�r�M����܆A�
�P�+,���F�G«\��ސ}��D@A�<�J�{W�l>�s�~�-���=�K�,�^hn�n$���Q���-S�@��67��9���ix#Xf�q�!�Jҏ3H8��7�p�g���r[}�|6�O�pAx8�Y���-ݔ�a]?��J�s�z����0��[9rI��>5'�PHrt��5GF=��J�=�Y��� r�����ܡ�J"��L��!���8�=K_���'¦8�G�6�g�@/F�xg����n���8���HJ����|��%��x��W��\ЧF��i
go����k�*CDbS�U=�x�-�D:����ڞy~�!U���M#D��9��z��6<��7��,�\ �}3i��?�����߫~/q�\?�~ɾΗ�b:�!�XK�n��9e�|����\��`��EIv�{��s�"��U��7���ƈ�����Y�.��B[�k5�ܔˀ�^�^����@La��M�]���:Ybϸ +�ƶ�I?*����W~D6��
T&uͪYRj�Z#�i��4����8�f ���J����~>�F���V-o�@���n���"ZU������P�|�q����O�娆,�C�D8�/M�`1��/8�[r"����8�P�\.��ܚ��;h�Q
3�f��*D^����*��Ô��g�Fv΁idUU�?Un/�z�[u^� $d�7�B�����MU�A2H�~�ܙ����'�<�Xl��(Q?���t1�Ul�&2�L��_�[��L}v�jp�>�,��{��y�U+��Hx<ŵ0����u��Fڒ?�({��.m�Sمo$<?�#?\�n<iP39������	x�7:K	x+�fg���w
������C�.0��
��'�g����.G�o���&��96�6	��D(��u|A`�ΐ F,[�(T9�q�x��I�d(�%n�oׇ�gx";�Bj�6�7�(���zeô�ɷ����{vr.Abg�$+���z�Cd��U%�αSKsϖ�b�"l��[զCLK�༿�V4L�E�Bq1�#�iIߙ*[MY�3r�m(�9����"V~9����������Qc�|b'J5��Б@!�%q_�J�%ڝ���� ���O#a��t�����>�4����_ͣ�b��(�ƥ��b�U����>�P�z�t��ȇا�{��< po��#$E'�L����z�J���&gv������Z�ZO:�A��a���(~�R ����>�7�bY�1"^���0}�n_�@ ��= 6�pԦa^�8�r)(v?#�_B�፠~�ĺKv��85��=���!�K��١Ҵ��lrL��+�4�8o,�:����`��謁��L�'��3����J/oY6�%8��`�B����v%=���p�M=6�-fǘ���q82!5�;}	�rG��"c�aqqC|��x��U ���MҖ���m�ďQ"D��_�b�/_f�l��(�<��4��!����u`�&��i�&a�ޛN�G����h�;p�X�,�[��*;?�E���l}}	�v���UP���h(��Vc�R���U��RI���/��NK�)d�����&�x�`��R ��X%�H�n��{��H�������(�2�(	@B�I�����$��2"袁o+�}-����V/��$T���ے��D��6�{�jÅ��C/<wo�s���ݽ�n���aVY�����EV�lb����2�(�y�G�!Ǥ�nx�P��JH��g���*���v����4%f}�	>�<Z=�t-�\�3Z{sNQ���CD���9=cU�I��3��w-�ҽH�B��D�6�鑱�Y�� ��6��F���=,�+I�I��_5x"�d�,6޸�ͳ@B��{6�Y��s����a�����|��'�³e6�w$[]u����'uL��w([��n}�����sK�SW���pF;-˲�7\�ؤ�x�6�Zu�+��<�P��q��3�M3}IL�g쯫���	���gbbCw�Y�P�ԉ.�{_c�;5����|�*���s8<�h_��fE�xd��@�/7�`޲01��$U�5��%U�7�!_��0Գ��/����|)U�~���/_�f%�}l��e�6����5�����p[����]�	�V%���s_�z�:��J�n���G��dv`��~��>Z�cs�U<����d��D4�;K�ۙ��*JS�S�8e6�=O���E��v��זZU�4��翛|1�/B�O��0����!�Qʭ��Q$R�4���w�.�C�h���M�˄���a�K��.|�UR
@�A2�L���}��JƘ�Lg�L�i_˅�]�*�i���q��K-OWw��U����z����ܤI�a%��Co�pE�O��Vb�'z��}{� 9�̩��{n��x�+\wݍM]����(�-��`U��5�/b�M"CC\>�s�� �&B�DF	x���jc�PX�]w���̗�XD9I��p�Vb0���4�S*-�����Ó�pr|1h������j;*���"�����}�����vq��q�Vn������Bi6��҈����TH��[lE��h?i.�I�.>��[�ʻ"�SllV3�n��(���`ҡkC���Q�1g��U�M~�-^�k���ٝ��橞��4����KoY�@����s� 	��dD�ǻ��Q�+��7�(ϔ�� ��$Q�4���s�W;�$Y��UA�C^q�581���ΤsF��:4=�k�4k�n{���ε �͜���h7���Xn:�KP[�O�R���>kG�\�һ�\���8 덚~r�8����_�=zMw�R4���u�0}@��s���q�k�1�}�,�̃��1��FV*7FmmR������A���պ��q�s���)>�?A�B�@�,'�l\�sB��/���pMk����������%e��:��Ui�Q���G^z���S��h��y3��Ճ,tG��M6fn� oq��j�7���)m�a��x*��R	o=}f��g�X?bT6���r,�;�D�^����!���3�/©�8�E�ێ\fX��+��%P������ �>��d��� ��O-���I򯨉��b�z�s�#�q�)c��9v���BDK'���Y��-�tc��o��<;���*�ܠ��K�.�����x�e������6�z�Y{O���콴�\W�WZX��L$kq�V��M�}��/�p�|��	�h��΢S�c��i����P��ŷ��K�[��&ZE_a1X�m���xH�բ_��6R!�FY4���D#�3�gj�� ��hj��0�䉯��Tb5O��ġ2
�����`��'Vv�[�i/v�/W�a�c�2���J�dHB��W;fY5�YJF�}n�V��]i�|H�+{��ǃi>�3�5�P�V�6��9�V��~�e��%,�ў���;'��IV�..4��(y&��ܣ�N�����HhmK�!�[�С.�=6&L�|�2(L���Dr�w�Eߠ~�?�f�G�d$t��T	#�e7\�������-8�g�-lc�4�!y��(�I�y/�_��w��[F�m�ƣma�`c�kj������Ȑ�\����(�U�J�s� �'��:�F��%�z�f���ŎV-zF�~�W�Ġt�g�+ �o�ԾQ�6`��H(��7g�������аV���L�si1�.ɍ&�� Cp��r��Y�ϒ �lB%�C�d��h(�F����窞"��Ố����w9*�@�Ez���A��[��r�?�E��]f���W�>xX남�*�$� ������l�c�|��	^�q�˟�C��ny�[��	��U��,x7z�G�{ڴ]�R�=K���(�.Da4�U ��@+�X¸i6vw
�p�����VVg]Kl-��(<*�D�D�Mf���?9��୩�sHʏ��@59$��:��c��\OYm�����X5�Ҷ���W�s-C?/Q*�j��"i6�ˏ
N�3d-c���u����$���d���w��螐�l�a�� o�߱$ʕ�6y"�_}�^����G�qDT��wd�Ȁ�#�0�y��״��0�!}+;�>�Խ��� �L�[��>����L��̤N�K� �d 6�)30F�
��l�J���C,��il��#�d�B)vU�D���C��G:=۰�ȶ�Re���ѭᝅt`����R�/T��O����<� /U��;���B�}���v0�^�z��u���䶚�m΀wrM�?H�A�l��oe����y���o�1���%U��k�Cq����^��r����~)�������Z��a���q�ld!��l�IW'�b����b��#n�	6f"#���U�#77�0i�b&���I�dYx*���D����
k�@+Z��Ҵ+�g��n܂)�,�cs�N���wf�2�v�fd�u숯���W��ff�9�N����x�Z��	��m%H�U�O��Rߔ	�L!-gԙ9���a7�8Y��흔o�X��:�+;�eϚ�q�rt6^ۉ��?VΝ̈́�N�\&���$g�N+����1r:��%��S�s�'��2� Q�?��+F�P�c��чA�x�d��E�DE�%+AL�=���7gM��?)!�7�!�>^���q緋ʧy�ǌ7܍T�h"=�v/�XK8�}�(���Q��$E�dݓ���X !���6�z$Wf�P��|��������U�a��#��
�N`G�����D�h[�iQ���V;K�I��^�q��#OMųq��ʅ�+�������<=��!_$K�kO��+nQ�|��w�6[]�A�駌;vcHZ�[��_�0.d��K=���ō/r�0���-ž*c�?��̷Za�U��0��(S5`"(�hsBc�������� qP������c�s�u�pf��-c�x�{G[��,�� ȥ׸�+�@Aow��X	��pى72��q'�
ԣ�Gn6?8�$��Z�T�	�Σ�C��Ǔ��R���f�Zސu4��3Z�t��hx}���;!{��j��"l�JT���yI{f5���aMQ��v\�,L]�D�i?9nu+����Rl�i4�ȑ�n���~T5��"�����s}D̀p�n� s���f�t��4$o�%"󩡵��t:�N�F�}PlJ\Ld�q�4�"�G�k�#+��P��ꧾY�e���35*rNG����W)���|T(��cz��zo�#��F�}��M"��S����O@�w��\�D)�d	E/�{w��F�]˙	7��H*��<y�}�!���m0c�x(j��"�%�D>�a@ɣ|��VŮ5����u�\�%�u)�Nݨ���5��m>�#G��`�1C6]�A��x@�X�S2#j�3�-/4:�mvj^�{��ba���X��lڔ`������.֘e^?Ag�k����Z�W�o8=E�4/�����!���(�Y�GN;!�yL�h���Y�i��Z�����D*��}�Y�f�1��n�Q�̃XHA�O��!ρ�:�1{R�d�E���m<���9ф�[vޘ�cuõÛe�;kB+%��v.�W4W5����&O�<��,r<MZnÈ�A%)V�Ъ��>��S��^ ��
�jKA����n�q�u]Rw.1W�Dg&�Fެfy9������ �G*�d�ˑ��a�1�BׇR�B�V�6�e�����+BXc����S�!q�q�D�`������Πy02������+>Qf������"��$w�n�.O��R���N�[�ti�
S�� .�]��x�&�Q�=�OgQ?��+1D�&8A�����=�0E�3(�t�X`���{��5�vU�<�TW2�wM�kY*�f��@�H@f�
.y�'V��$�R�*�#8]��rb��Rf�k�mRJ�������պ V�5;G.�8;-������2a�yCO��(>�� ���zWפh�Mjk<]$}:�f�N����{z^h���������@"���Q�����hΛ֧��0<�n�ʾv���}(a	�q����J�͖�1�����⬙v�k�_�QU�j�ZP�Y~��y��~Q*�f��J�;^&�ۀJp�C�T��|�į8�9#�N����)���@s`�U� �l<�b��R��?�?����=�ײ��h�4\5�M�ں7*ȓ�d�WJu=�h�S~�A�����|���W�qЈ�����A絔Z�z@Y�l��V���'Qah��ƖB6�(�R��2�݂�c#�D@�����<91�O�$�~���G&��o ��z����v�m��QP�.XK����A�"#��'���΅ 퇜��;�>e�D�t:�Uy<�*�L�&���f!���	T$x3b��!�hÄL�"Np&D��-��.�	���$�p��3��4_U˅�Ǩ�!^ň��:yt<k�9y4�?��vk3�ly��J\k�����`�����-Pi�k$zFg�+n�sr�o
���BԠdP�Xɯ�}ɍLx"��䁷�bqE����@�2��=��[/�MNZ3L7ر��7Fz�C�>���q�^�H;�#d�Kz[��头��zt"CS�N���.{l��1s{Ȼ
��)1W�̯�v���>T5;�=�KS+�k��$i0�H8Ȕ��3z.����11��-����_�i��EZ��,��1���keߊ40FP��cAt�F�#R�3��"�9۽��[9}5*d���sfP=�-	d�����v�����W��7#E5̘���M�V�U�bx��c�*�2���'c�o�c��L��BG��S���O��%=]�P��ύG��zu�xфӴ6,�"������wXc˙��ᡤ���(�xgLN:< N���aJiRM
_���� \�ON/�1�@̗����al�q���5�AmBz6�Y����k�3(�3Ϣ���64M=^����4�w�:Y�M��y=#���ndz�=��?GMg_T�!+��h&��Ήww��![�$�)HC�J7:L\��ƚ�2�@S2j�%[�d��_����t	�vc�b|�8v�3-���?׌֔�{��R��	�:���*�r�+v-�z�..�%�H�^	�7�)�U~>�e�U&N�ww�Bz��ٰ	q"~0�����~־�3�����ڬ\أ.	�*l�Q��3�ZP��9L^%�g�Ծ�mqHy_5`Bk�TA���h�M���)"�W�7�p���<���(Y�'��ܡ۹9N(�:��$0!�n���/���#�ñn��j
�����5�D-��T�ռ�ۼ��f^H�*x�N�YZ�/�t���U�7��ld�i��"���wx�Ď��'A�	&N�7��r?���T�#���X�1n���[K�zeTZpY��
��rp���4i2�iL���u/bVh�@�x@V�M^�k������'/�5p��q#�l吳{S�Љ�b�[\F>�j[��&�cCZs��ҥWm��:0X�-G�E�$?>��XJ(E˳8��L� ����b��oI�� ������ĺx�!("��d���^m/)�Ӌ� ��i<�{�9_)����Oeb�����;qtX�4����~!���(\�����	ܽ	N[��i"�E�j�E����]q���Z\?��ӊ���/�}QToôL�3N�O�}"Y;?�>8?�qL#2��8��<�6-�;�{6|IwTi�7�9�` �2���Ŭfq�R���a�����Ҭ�#�#����a��L�M���<<n��UJ�Nh�<ûF���Y6��"�C����I�)4`y��h�ӂ��[ڐhr�c���j���/�| ������Y��6p&c� 3�1Do<�6y���?��k9P����YBJ:c��X�󤞘wb��yw�X��	����9�lQê�L�[ ]:M�K)�8n8�;Z��%{n�zLᇨ�VH�L�j�U~C<��>�rv�GA�,L5��捗B�R\]ans�	pA<k�jv��:K���P��d�
Y�H��N<|�_N �����~��a�ԥ�ib������c�i�����CѾD�",��]]����l��.a;g_$����ێZ4�f���~��}9�;�Q���ԮD�^U�.o�G�a��![�$� �ӥ-52Ӫ�R��y�:�P��QBN�>��XbqRX�U�cJ& 1\������qر���0?�,!~���N�:ae�-m��#��D�U��L�ζ\Qhu/~|g"?Ĳ7�����|�g�<��ؕ��]^�: ����h	+�v�:�:�DF�&
��A%�o�uKEA-�� �0�&����	�b�������L����R��
�M	�Xe�̗_K���F�R�XCj�'s����9�c���Cp?&7��Iq��}��Ev!ž�5H��*㨽�U���>��FB��y{o���y���jd��Y��9��6��յ�X�ݗ�wpZl	����@�D�k9���h�(w�=jF�Θ4i�5�R���@�-�����7JPofT}A��ba�$���g���E�R�SnR*Ɵ� ��37n�WE���LK6S>��EZ^�M2	�&�钼�ϧ���ϫ�T��E���ćb�n� �Ry_7�G�!���j��d�*͏إ�j֤+��:g���]!Z�"���b�[L7-:j�$�����L78v�Ql����&�,����2K�C�g^&�,?���S��>�w>s��a�b��GB�|7U�������Vt�C+v�Q�1a���>�F��ZaΗ`+��t6�.r~*�Z:K����C4�Ӕ�Y�Z�LE����ٲJ�e�PG�%4��tGt�����l��	�笄�6�����.[��[R�*���<DNl�kLh�����%(����w�do@X�`�D��nS��"���:�9h�)6<�ә���cg��}�}Zq��)?��N�@��(ʹe�(�g7��b�	���������]�tAZe~4�Q(�H�Χ��I���^��T�] `��I�WS�3�hQ2Q1e�����bXy�.l!>��kB����K@���E�0\a�:����f�}�Ti�AZsEɾ��U�D:Cd��Z����� �8�vGbc}��{��������E�h���$�y�a�H��~� _e�2�X�K�WxO�2�y�KPM�\�J|h/���}��E~A�м��#�P�P���z#�;���tX�H���l��l;��A�0R~6�^�ѵi�p������>;|�~~��ۣD	�ک���B�$�"pY�'+����~-p��1zբm53��hlR_��@5P�Օ�?S���A�D�NY��qgܛ��r�dQB��k=޵���܁~���N�}t�~,�^ ����!P��������	z�����P���w�*F�['������)Ƕ�v������8\@ٸn�n7�ݾa�Eu�H���$����f���-�1uK5��;�(�<��=6�x9n�a�RPzR@���$�Q4#��m�;�GFh���m��X�0��Ua>d�Cݘ��G�$0�y��I9�@XK�a`�K@V����aWoC�LY�L*��p�W��u\��%9,�,�͆�ަf�F�+���tzN�mw�ܒ1C�#���c����1��݀JQ�Y0��.�p�)n8�PR�R�p�n����M0E����:�8��[����/���i�&?IS�bL�wR[9�\��y��e2k���p��O3u�[��\���	����C���:0��G[����^L�5���z�{�e�����[��&���r�:�w����G�zsuQE��y ��H@c؊�bce~=��xvtm�%JU���p4)UԷ��ى�-'N?�Op8�Y��<��.��8{�0���C.�P�-��D�B
EL�1�<�TbDdN�J������ܞ���Ѝ����	YX��gl˨JT���ol;���N��C���T@����_�Z���_���M��u�f��������~��߯�k�ѩx�Q�{��r҅�cJչ�[[�-'>�7C��+ggcq��1l5 �\�z�j,{g��;�r����F�q:��zkG��)8R��?����(~ �Vu�[�����T.z�)��G�=z�����^�'�*zI�.LaW@�T
�v �	Nm$$�@�?�*�	�tզ��f��H#�_8}��ql_��G�N��Uw^���k�1��\`�>}�o&�	(T��d�LaP��l�;]�b��Z�s(���^� ���O�QEhh�#��t}=U0[��}b�6oF֜z�c�$��>Y�]MT�g�X��9����N�q ��!fV�� k�0�tH� ���\�d�ؙ[��������j�i#��)2o��=`}+���m�wG賛Q����q�a"�7����7��'��Y�3�5H�����z�ea J)�jH�-����'��/������h�P_S����R�c��b��U���&�;��Ab��*G�]̣y��BhU(�F7B�-�sZQupq��nƛ�7c��Ci��W�eߗ����BJ����H���1��#N�nqx滋��b]!����[&!1z�̹l��^�� k�i�C!��j��;�g�@��A�h�;�RP����>O���_e�<�Cc9��E߇�|�d��%m���>��c[��
�AW�'?�!��0��ҌFz�>����4y;ޚbSᧉ���aޏcSL���m���qa�I;�J��6��-	���M��E�p۰��@V�,�v��t%2�&��ze����˦��
2�(�&��<�.L�<��Bǔ����q>��� .��J8��>�Kl�Tj9"(���ac����R��T^l�Ldd1�׬?�Z���A���(P�\����
��hĶ�&�1�C����L����͌W�\FY��䔹�ky���m����z��|T�Ud�0�M��P�l�_ �_R�
�����<#�{�Wpc�B�B��I`��].�#K��=�[mX�-۾�y���(X�h�Ʌ N<=����<���I/�G�4k�����m�3��,`�M����5m"�OW�{�F�y�w���/0ba� B0���w�������;��#i�BW�`��0��i�`�Q8�^�}9(��0�Ͽ�����A�μ1�\N�+���Ԕ����f��V;-*U|�wIk�&.z���">�(�S浅��(�����F̽�^Q��/�+$����o�s�q|���d�/��<����پ��W>���1���n����#���xcǿn�0������6��S�3P�/̐k�W��yH�g1�=�ĺ��3�+�>�X����ک��e�p�x+��$r�s�2��BLZ�Pu��]uC�U����t��bL�hGRsf9��X���Wi�����Tz����,��'�Z(��a���,擊�'[�g�{#��r��Ћ'�ȃEΓ�j?Y�h3��(��R\<�J؊c�b�g��:�AA+����	���c$mvá���L4��7�p������X��2`�Z>�Z�Jd�>�r:!�bR�����]�h�=��(m��ؒB��y�neC����S�:w8�P�I�AYn�cS�=%X-Qc��lt��F��pXu�����9 � ĒOr/��U@��t��B�8fxD�[ǜiZ����j�~�5�8�౯����ڇj3�xmux��G9ٽ�Cی�2��A�S�w��e��|�n��z�Q��͚F
�i0t+E�鿢����o��% �������C��c�>U�[��B�����A�ȇ�؂
�X�D�/o����񫭂C��R��Y��؄��GYkɛR]p��_Z�-���s��,/��N��!�,t��e;�^O��y�-�=We�fG/���ĩ}̃��'��u?�DF�p�F9<%dҋM@�w�.}>o��N� o>���J�b��șf9�~A���U��^�[�%ј���0	��k��A�%J2:hK̈N� �.ι��YUA��4�.Su�.P�t��RY~�G�<�޼9b>C���(N�\�E�~�ȿ����}�w���ޅ��4�ԫ���`�uu�[�iP�vx����)���'q 7m�m�a�� ��Tk���r!B?H�(R�y���m������=�+�k?��>��4X�0,�y��4��Y��zN�fc[a�>�U9tx���� �kh�$�4k�/lo�S~��w��s�za���f��	�T���j$-�X�P�_j�H߂"\%N/�u�G>Ae��_���a�u��f�R��'�齵,��:�����F �����ܘyX��fa]�����A��X,�%�����6�����0	�[=v�L�G�W J�!����w���J=c  ��ۍz�ڻ7��sgPbH�QXs�Ȫ�.�k5"i5��4%s���@�]�ë���r�+�n������7R�a�O(��>2P{KT��_�I�+�,|+�+1	�P�+y�s��e�}�~�k�a醃���,�'�l���-��\����V�4�o�Lk>�a+�ܫي����q4.B5,}���cc��;�ߛV8ac�w��>ë�@n��xh����D#+0�>6*��y3�׆}Ա��S�J"m�u�B�$h9 ��6ئ�����^V�{>�t�B���?*��S3S���`�kX��S0�|j^7�_9���$xWo�[l��2o�K�A�!��f�R���*/S8 ��q�!����a�S۬�U'}�z���yx�z���krgm}�"���}����1��(�y����,a�R��"��> 6�OOv��%���M#���-�N6���E>�����t�O0!�#L6R�!JJ,\A�d9��8���m��ۿ��`+�p'� �?Sw�K�ʐ�a��{z;B�Th���ˑ*�����X�Ӎ�u���)G)[|��H?P��}��$�Ht�leN�Zэ����mX�]ɴ�1L/���(j\5�S<U���a�t���]��Ѫ��	|�X��Fd�՗�G����=m\����+�������N t�"���F�P���y�P(sj,�]C���$��a��:��c<�1�[���6���s-�����):p�75���:��e�*7)�6�"!n��Ť�(��2U�����y���oJRP��4ClE�i�
oM����f�%`o(�Z� e:o��×�$���y��7s��]�=;���4�z��	��J��~^r�}�����9L�8�n-��ɏD|�P@R����W(�(һ���zÒ�I|�R���*-Scj��͠�?��۷b�`���E/�]�$璀�:����o��I�w߆��M��/��u�3�H8q�����]�(��f�Td���&J4r}~ �F�QWb=nq</�'�*f��$T�Ç!,�u|�^���'���zD`���� j���B� �eόQ_2�4@g�/2�k՚�Rȃ|O5V�E~����,Gwl�����>cP���_s��4���v�����yqh�l%�@��CG�r�h����J��� ��Ʋ��%@:+)T?"�^]������
�ρ��m�n�"�����/�2�b���r�~-E���Wa����|�c��Ϡ���Q"��jize�<��d�mc-3��}W��ո�����<-]�;�0F�8a�D������7�i�����YBV}�w�I���_��e=�Y?l�U���x�'�����E �eΚ帣b��˧Un�AO�6�j��	��������-a�o��p�t.4���%Z_�*鈣��-��Y�e�����7q�����U��]*�1[�K)w�؉<���\��
.��ų���PI�><p���-�Aߜ�A7�YDb�_��a���Z=�`�k�e�Q8�!߶!A�_�a��{�p`Evߎ�T�R���CpL����P˙^�Ă��@�:w�rqx����{]��j�5��BL�X�������kcH���ԽcE�R9�IB�F��p*��q�|���t%����$ά"Y1��x�w���)	�i�W#X�UC����XN�4�`��dbjv�T>���냧5()I9d(�P�E
M��+�g�u�m�R�� �ݮ�Q���v�^ϛ���y9���O@�㫭�Yz#�?ɲ��o["�i��fl!��N���Ɂ���&��`-4
N�9�#6&ΰY5@B2�jj�h��G���h�~@���|��]���Z�¤�RǿO�Wi��ל+��{-@�f�+�^��|o�p��+�9�Oǁ���V���Gi���p��l箬�3ܦ��]6΋Tв�j��%���Z�b�����k�<!��u�'�ƚ�I��U��>����FyXU����^,�*?,ޟ��1\\��vT��q��F�Σ^f3��������]� 5���<��T�b9������Z�s-��-�";^|
��+T?-�*t«���e�b���������M��|�Et/�:�S��R7d��VVb�A�<�t�c��@X�����g�v�&<^r�|�w��M��F#H^(|��l���[+@9nq�ݯ��]�C�an�����V�h��F����=c������v �S�m�U�1�,@�z\6�69;���u�����n��޷�Y�=����w�x�y� ��-%N}�Î�a��������>ҋ���O��-��EY��m���+�t0��p�;R��� �r��L^eEo�Ck�s�oUe�X�v	�ʽ�$�z̢(� 'UX���p.�|�D�a&l�%`�(�L�,�
�}��	���K?u���밥 @��C��.�i=������W�}��ӟ��FkuQ�Rõc�v�a����-O߻,���wC��.M�?2zĀ1���Z�z��{K���{�҂@��u�R	�9�VY�;`8�!|��}I�`u�s�l�m4�tє�ٝ�(92�C	��*�7"�y���>|`sω!�y��'�t����u�_
m"�F6\,� 0�!1}hS)o\��.�#8�k��M%a&�^��a��F�hN�#�#n�Hhba�i��%?�rﰟ����6\����b�S��Q����%�8��Y�l���P��jkU�cY����Ho.d't�T��iI.��]���h?$�w`cpO����<l����螧�>1)06�:̱༎#���-[�� fJ�M9��
�M�߬8��?��|����t�1�O��g�s�o�G�Y�8+��Ic���/`	��)�G|�J�ꢏ���w�h��NEMw��љQ��1&��ʏA�x��t~6��^h���]0�|�E�@0��瑈�Ợ�c��-����J�S=:�� �s�[���g�q�JWI�s�҇c�i^����R$���舮˚�C�3-�&@���-dNkr:fU>��-+�~>�a��ҩE�L�� �-�Nd��`�;DF]d���T��L�����'D�&�2sO�b<�=i�al���J����ٿg�)�zDǱ�5��xs�!��̈́��u{L�?̥�$� ,{�¡�1 X�\=�x��L�Q�Oٺ�Z���d�����p^F��ҊD���Mc���@5�_��B�kz��2I˄��atўtH&�����S�L�yҝ�z8�b��U-�(y����Ϫl���#>K
�h���>��%�\�TC�(0���D+{�Ẇ.����DpCύ���^M�^<}}�ٻu{�@d櫀
�U��p�g��=p��˽:@��8[�t�>��̵k=�mO�_0��F�I���K�9��N��,C�%�9�������ѨT<[�]�,�~7�ɏ �%^�,�TP nɗ��3�W	z�Ҳ�U��E�8�jB�-�S+z5��n�\�����c��c���SU\�F�݂���d���W���g�k�")Ѩ�h��0eM/�#���6A���骾&�M�g>����'�fu�alҭ��@�&ǞR�.�O�$�q@�A�gtj$�J���~�Ċ"��1�-��>�?w�X����O}��d������g6��`��^|��b';"��&���x�	��-���C'l�4Z�9��
�����G �P/+��c����FS����q��E��I���ڜ��`�:�O\���b��`�S�8��/�aq�iu"�⟃˕�猴l�E�9��,��|i��ܮ/RS��B�6�2@�p�r� ��⣍���!���=���E�?焃�.
�$�9U��Oxy���>��--��D�-S��)��:F��*[q8A���_>�3{����~��㤿�Z43PS��0��`2����[�(vA��q,҅ZE.b֑.�9��	�����Cȅ�F�o`�T���c�_:^Р���堎�䝒�P���U��&�^��P��2�Z�de!\|��y�v����M��Ow�w�D�nO�n�&d?n�g���ݴ����Za���*�i�:I�믾�����Q]!h��v ���!��vsI\��h�������%T�T;}Zh�֢�sͱ���i�����[�K�;�7��Z�ru%���#ě���������1��6�g�V�9��_�fɼ����sW�9+���X]�V���cp�~�)���5�.�qzu��R�
jfo�|���M��5��$d��Z�1d�`��8i�D��5ߧ�0l؟>�u��UC_i��Ov���V�H6['Y76��͋YK(oHhLJ��yٝ�4]Ӂ,�h, ���n�6�x�j�Q����F�i�gB�tf+RY
Q>��ϣ�RQ��"��t�ݐ91:�Y��d��N���o���nؓT�"Nbh�����z|�)p(��SHzB�X��V���bHsiІ�����!E�Zb�W��:nXŀ���ؘs���v��|�q���X�t}Nz�F�b��W�c�����&�l�Lg�>���6��>m'� 4:�6�s�&~=y�W��nd�%�4�C-y�o�_Lp�qߒ9�����q,�J��r=�7C{�Ka%������E2�*m�_e�l��^����k=�%b}�a�[���K�N�ɜ���@�6���j����tz8[|]'�)ԃ�cv���,j��%etO�盚���f�������6O�+�P������v�_W�M9g+p�a+�҈��FA��nʓ��Ǟ��ν%�Gɓ��w��B�e��J�Ȳٽ,��n.�6Ӭ�\������eQ�)�c_DB{��R��t��o��q_ӈC�������h6.�t���	�Jo��y���u�����/["��R��}��m�H�� ���^�@�w�ʅ�����
z�)%�w�`��и4|i��X���I������r�b�P�h,X�?>�"��������5�N� ,��5�^K*���x��i�������K�
�ӵ�"ٿף��3����6��r(>�[y�86��"%��[8�Eb=0O��"�AO���B_?&l�%l-�<7�ů��TN���?D"${��Q��N ��=���O��"�?�7c1y;�G綮����so(�E��(�ѹ ���Ǧ�O�������>�wA/GҮ�JFCڐ�|{XP9ѡ��_3�}���j��UF�ܸ4�@V��2Q$�QЌ�d�{��b��P�G�ψ����� �,i$�Ի��S�5�&kM|�é���bf�>�=f�Y���>��jߢ�6��r��c7I a��"��N�w�f�cS96Y��S>�K��+3����x�&3Q�GC�hd�8?�ܶ�eƼm��dz�W�šs��i� o��*��;~���d��z��m�OOr)B��k6��+s<����J�{΂�o�~AtJ�?�l�^�$E�+v��̂m��hfh&lgV����;Ԇb4�Τ��%{O^�c�.1+��%���k���/�E�5��ps���S�40pŎ�1և�c ����hu��DXMcѭ�"�H�
1�|�Ş�^OM@�Yqw�d�����ۼ��fS �?]'��i4�%yQB���W���٧=l����|?4o�RX.uV��d�<��@&����K�!�(6=ټ��g�9�ʲߩ;�S��Z��x�2��ZC˗�yHBnL�k�v�)�2�G(qABى������{���sG��s�@pސ��	?(=��j�9��|1#�w�yA {y�h����'�_[�`����3�×���\��z�@ܜ���[S�`u����sW�z��!�ؐ�1�q
�Z`ø�'ߩQ��lS/}>�R�6&��A�h%��n�ݶ��'�J�d�&p���(8}�FX�����?��� ����o�6)�YЧRUi�@��?!҃�4f/4ѱ|"���V��LxY��ܷa3�ɕX�!:JE�i��p��f�"Г gD~�b3o���A���M��7A!��9ֳ�q��Q������x42�m��C��wIj�_�7/��2$�J�����!Aƚ��;^E��7G��|��DÕ�.T7G���J���
��Q+R�D��)�D�b��c[M�
�����~��+)��G���hZ�継��$��L7Uf2�^=��Gq��K���1��]?������2<3B�kaK�y/r&UX�L&7Y���su��&�-ڋ�e��}v�*V��rf��$1��6I��+�QH���$Z?ԝ
����y%�z���D��l� J�6U��K�dH��Q�#ѧ�S #T.;k.���;sC�K�[��K��L�i�X-�\�_x�$U_:�['x,�cf=�TVv^�Y��x@����oc99@�����1�{��C�j����U�d�<ٸ�J_jt��M���x��%H=Ӯ��2�;y'p>�e�u�̘��6�<`�
�'u�vq�@)���`@Lo+2j�S}���tp��X;����,�"�\3 ?a�c�V�e�b��Y4h5�r��e�N��D>��r�}����g������h>��ݏ�o�Ð:��ojk9{l��ʩ� \[@o��̭���V)�U�&^
�P�G�� ߆�!D�s�g=Ⱦб��v.�f��`�>ʔ�a/��16��`?�+�q�4k�}��b�*0�6��"���4�a	���Fԁ�w ��O�D�M$&g�-y5��/�þ��[Q��W�>�[c��r���֞'	o߂��(:$%�gy������K`PK��tM ���46z����z{$�r~g=]��lXүH(�!�3�)��L.�ڔX��ႁ� ���5���-W�}VH�Ħ��-�Q�U��z���NI��d����Vj�I�����J�w����#��A����vq*쑄 �tL�s�p�xܝ:����q��3x�
��WsJz�ñBN��E��=s��K��o��#�k"��g�&8�͗#B�_�?�{���8���u$��}5�c������K��Y�"dU��W^=�L6��Q�;e�x"NZpJ)�[v-��z2�r�8����<��Y���n�y��� �O���*�\�%�]��.����,0&�5�da��݆?��Ӈ��w�>�>H�7�j��e;�dh[4�Ŝ��p�r�|��E�u`������c^/|Qc&�q޵��+Kt��-�}	��0Hj�MJVNy;�B����Qiq�]�W�?��լ����F0��ϿGފ��*��w�Bao80�i���mzKf��Dmw���2C͸F�熹�.<�FrvM��~E�ў��?�g@J6���Q�FV}=��}�O ra_�v�����X(C��s�2�����߱[R��ur�3��NE}�MS�bR�깒�FLu�`y�TJ�m"���k�Z���!�qM-��	����I�$�e�w]��v*����-��"�����&�c[�[��ی��>���`6�c���o(�Է	& �����D��Ֆ�E���[�?%�Q��\L���9Ѹ��R5ҫrCT��z�#�Z�O�`����N=&�:`R�zg-2�?R�2�$���ꊲ:��Q���dtK2r�_w``Wށ��?�虹U��vY�6��U���k�sΕ-��`��yr;l`�S�)ѯ_X��BsZK@x�(�F����̎�_.讋L�\�(g.��:�]�C�o�������{Ү�k�G�U��b>HN^Q��:��:!I ӫ��������l<��,�L�6��t64�\���0�R?�ә���[B�R~�i�1���U}��r�����~���V���ls&�4	���R���W�	P�q�%�J�R]XFq��K��
��vF��C���Y������`,g��U7����%��M�5(:m���
�����f������/�Nim��^۪����T0d탱�0qQ9�R�q��x����ޛ��Ⱥ�g8��
�s6�lwƣ�V������ua����D0�g�#��d�ON��p	#�����0,>��!����wN�v,sy�NF���
A���	��W
�Tl$g(%.!�P�e�19����N��[3&������^^�����)z<��S�efV���΋_�-�O�%TQ��污� d��O0�s*�2n�%^
�9L,������}:�5@�a�M��6�a_E�/��}O����M%�;�9�h�.ڏL�����hl�ƭ����-�CNYqcY�I����ق���5�VE�ꉡK�G�7��vMf�+�dＥ9�$�M�O]������Y�h =�B�Ζ���c��a���߬C�Lì�;]H/l�"��,K��\�{!��X�}G+���c}XyJ�s���^��h^:�(��f!�?�[K
��=�ŉ�b��Q���蟰�����_����q��`��d3>尬pDt�@ǀŨG]�I�,�Q�/mwx��G���O!�����E�Hw�Gu��E�{r�#x����b]��v$71�T���_���d���Q�db���Z�(�ƕܺ�h~�{P�= ]� ���MQ������1���WkA�XZ�bTFcM��r���q�nX^�������pT��tܿ�ي��Ja��-̤�FmOW����iI׼|6xr���܍�,�PQ:5$}��l���m/;�X�>������t�=16�NF�x����T%�� 8q����n+Z�+�C����D%I�Cc\+�඙��B��Ҫ:'+��2�[�9�C�����6��pD�r]j�F#DH�����Җ�2��C���"�e�i�}ls��{yxw�c��Ԕ��/AO^ �ꅲ/�k~�Gc9����>%.j�i�<�Wo'�U�\8&��֕]�*�ե$n1�6%�����#��D�ɒ^����n�7���R�3:����^šQFu2�l^j~e0�������i;쟧�����9��{�ȭ.A�oȬp��;�):�΋(��V�k�׸��2���H�r�>)����`�sgp�b=	W��\�;��gI7�rm�8<L�Q4N�2^TХ	:�7���������N�����c�?!˴� V�,jK�9�3ޗ�,}�c�e����xTG��J�iR��]ٿa;M˥�lb��ggETJf�}�$Q^Js��Ko����}|
(���h3"88���5 -?�س�.{���,��B��y�ʲK0��lI%@�G��b�P��<�$��	��M���,��j�`������M�
�e��)�/�[M0�Z�6
[\��|�I�?�vk�J�)Ҙ�z��sg^`�1�@>t�q2 ��}�N��2�ޣB���8�Y�g� (ܻ��1x	��u�8M����H�O��{l�)[$︰O���;�4�Д̌ĦF��>�S�V,������A�G9h+�v2�_d�iz����9_!�4����f?r��;�cX\�J�4�(}4`W4��Q��}�!�-��|W�̸Fl��\z:Z�^���k���Z�XD�$�:.�m1k�QiG�T1tX;up.`C�N�kzQ��W��{5�e��6t����L�k����P�"x�h>K^$�!�)�B��^��E�@��;1�$��%F�?<�bd8�Q�u����<���=$�OAP5)������ˑ7�=��'�ĩ��C�8?7��c�=��4T	f�ut�k��8�*w�EVrڻ O�<M2b~2蚮tL�1L���Gg����/�䱤����4�s�.�|Ls��mC򿎱Qݲc^���M�F���cr���p��N�����u>*�# ?lu:�k�"F�ji�i���pU����_8H�0��=�lY9ќϛ�����CB�u�dؠ��f��z�>b_!M>:�H����//�s�L*���
��+Lz�h��e���)��[O(T���	��g��s�0�qK=�';�K9�r��ކ�Z��e��@k�o&��9b�-���׭`G��M����-�ǉX�U� W��L���z�ma���;:j��t3���ӑj�����~�ۏ���K��QAQ� U�L��^@f�����m�n!K����Dtg���r�j|�H��g\����� ��u�J��$��#�q)*r��QZkVl�yO���[��n�6�nc��/z��]��y��$���c���l�1Ũ�U`�hO�����%�����w����l;�7���(Х)���<K/y��i��t���<1�kE�XٸK#���R�0$ Վh&��n�C�*�-FZH�ՄAbO{�`ѝ��8�v���E[!�����%H!9�t�����m͵�Zy�뾠f4�1,,��i�o-��vh3����h��_2!�p��\���'�� `���g��\�!1��ǃC�W���x �Kc���H+;��)]��",n�$fjˊ�N�|DЏ���/KDp�����)�8?���?�^J�v��,��j�3���DQ�O:aI��8T��(yj~���7��W�}����n�9��u?���`��Vӽ���6Ʊ�F`mt��Z��ތ�T�qm����FϿ�]��'8����:��ys���j��p��?����2���Uɾ��^'M'C��H;D�W 'v�Ť��g8*9�9���(�џRXE���DR�郻�!߉�sY׷����g�A�iu⊩/�D/��o�L)��̋%o����!�i���ff��)zXb� ��j�����*�р�i��JW�����\�7��p7]=��t�7aG�<Z��b��Y�Âko>Q�Z�L�_˨,�k�د���)������)�K��W�p;�Њ����]�u�j��%�[Q�2C�#����ܕ�y�����.�g�H�j8B������nC��hL[��и�J�z��j��!�k���~��4r�����@���_\��Lմl�]$po��ء~[�ǓL�q#����fDG�+#�7���WT�2>�$)L��qs&k�ۑs*��/W��	��'z�q��ô�@��^C�x�#��4w����u�bWn�	Y,�a���>_38Qs+�q�}&���x�Bn~����g������j<�a���'�֨Ԫz�
Q�E/���ߵRy��l�s���@(̷`�yŪO0i��_�B���L�Y��
��R�t�\�,�}Ǚ(\���f!�OFҸ2ϲ/�=2�W��!xD���N�D��mJ��g'�ծ!�}!9BċzS�����H�K�^yB*���Vc=O��>x�U��"C�j� ���_ �aӸ��ИqB�_�ꆚ����蒼4�f?(n_U�����{X� J�8���=�5�5�tz��Vb=Lۘ��4��b�B=/E�U�bk�6�ة�E��rУ1y>��0���k��]��P]�'�?.4˘�EWo]�ra�^ߑ���!sFd���M�^���E�(`�=8�Ϧ��`�RTo�ߴ�(����P
��	!����"3��nY���7l�ks���?C��:zd���0�|�x�HDQ��#w��m���aԄ
r5D��@����jAu�z�a�U/�MGbW��A�=�iuQ{"Ô{:��9�s�ſYHCi�ǽk,�;2�}J#��gI'f�I>p�É��C���_�j]m��_
���?���"\�h�>��!��W���-��i�Q��R�wn��~��xy�C_�M.�G��p��_�y�h�6����#h�"����M��\ޥ/Z�?0"Mj�v���>�Gc:f�����E?�iIx�q|IP���)f����+U֣]���	S�D��\���z*~�1;����;��C_+�> ��3��c�:�=J�Աr'E���݈�X��NK��K�;\4��x��uR�#�^��w�.�c��(�KGX�Ѕ,�d�A�a^�U�vJ(��VT!L�T�@;��tp_���4x�	�`<@3����-��Z���u]�C�,И�d��A�9[7��cQ4tK-��:?2�K%�����w�vi�үޱ�i�K��/����ȑ���n1P�A�'[>#(�-vs�8?�A�9c·���rQҢ��-W\0Yg�1|}'������r2+��N ���"u ���K�_5��L��_����`�HUC[�,�4_3pw�Qi�Q&^m�Sj���6[�#�$��p]�㹛�o��n�	!����4��_�](F�E"G��1�m��cR!���-�]�"��\o�ͳ�0�ֵ�|�:�m;��C*o�Q����N��y4	���Vzk�R�Vt[X*��;=�������8B>����qJv��Y�ʤ�hQ��:�Q�^�M���q�B_$�5Z:��(M���+(�x��9�"�j��Q��!�V�%V�.�|�Bac1�S��%h��x�� J0:��1-�V�&��FX���?Rg�jʝ{����7v��R�+�d�"
ԚEcF�"JY}p��%ѝ���4P�m1�Qx���7�O���˄!֛�MK�n� �d�Ťp�� q�ь2 ���f�	
3f�f�O@��2͒�Ю5���<���Lq@ް��l��J����ڗSs�T�`�5bLsU���A�/b%cgc�X

�1�+��.�Q�S_�B�|^m((�It�s�[yHr]� �W��T+;�Q����y��	�w����R��5#���)n�L��J��wmGN�����tgZ*d���5`�
h[[{�y�5/��AdU̳Bi�L�$6����xo>�`2�P
�^z���$���7�c��r�W�m�X'���L�	[�纅c*�iSW���瓪	ǘ����3d�-)�ѯ��q?�����&T` ��#��Ȍ��v^���5��~�V=�Ds�6��=����Z��\��G�q1�Je�8�=Tz$G� {w/��<ׅ�Hp��|9��# �8�����9�u�$F�wG9�`4��vL`��~5��^�����#���%d�Hj�K��H)ο0����3���!�������~�HF�'��5�~I�I��a|��",^D�e-�F-���x^�[�^X=���W��?�M7 (�AY#$]�12�h�L�	�������@�更���b^�s� *�l.����ͅ,�u:b�ۦ<�� ���j����^� a���o��+P+�J�/��K+e.2��y��9d4ja2~Xg�Z��|W-s�^��sI���"2\�]#���X�X�Fch�%��Z�x�?4g���Q�܇�*L����s�=ۓJ�%��R˾	��A �1�[��UIh���w�ջ�U��ф� 6��ܕ�2�+�F&I���`t��KT���^��<��6R�[j��fI\����.jd�SD��"XYK�F�o'��>q�����樇T�6��NM}������������HIo�>�]�&E�o�����P㷭=5�,���!̀�yo�W�QvPKą\j���n���x�� x?�6�9��n���i�\�/¸Im�iV-YSH���%ҵ!�B���(itbi�M���L��P�/�Ir��)���f�t�F��)7�v�xT%�W�,rS�.�m���ڃ�˲���X�:�rx$ہ���g��I�5��~���k�gº��s��3����9��i�O.�(Y���A�=dc��8��
P5��ǽ�_����9�~��o�#p�=K����c���E."J����;����pS�[b���e^t:U��n%S��6� ]w2�5=�	�-b��@.ŀ���Z#���w6�m�l?����Q^�F�G P�%_�6��m�O����c��H ;TZ�Z�Շ}���3��]Āz��( y/��+Q|���ʃ�gT*#���,�U/�R����)��3�b��_dec�I4�5e퐊m+s'�;�����
��lyL�9ѽ�O�8��'���`^���ʢ���$�Z�ܒ�z��s���/�vǐ�L738shf]h������[��B���֢�0؍��^����BK��/T���9��mq%�z`��W�b���u)OE��3�K*-̓���K�܅8qc�wU�:� ���� �0I�DD@a�e��z�*���F����p�*kS���ax����΋�,��B��`�$F^�\>��p8?/��Q<^ɡ:]n�AE��Q�U[s/�F�QV�+.�.�,X6���L��
W4�'�4Vtj".򱛱ѳ�b�|UDSn��pkj-�y�S���J��K��h�c��	��q<���	ٜW��Ѯ2�ͷ��W$;T�A�,���ǀ8uW�F�s?�%�9 �A�3����)咷�&t�C)�D�;��@@C)�L�=7Wh��V������*1m
GPS;fQ��CE���a�?2+��@�S3S�k�<��f#1�骲-��sLe�����_�Y�V�Ȝ�
.@�Mi���ڋW95���XN���u�����/g��3��X]�(
��n��Lx��U1�}[ƪ���o�5�"˩>^�z����s4@���ʨ����ܵ�<x�09,��ÿ�Sd~�x�7mWJ��nkMc�C�!F�ɡWG<QT�(�Z�7��7p�RF���W���_�+�*:��	�?�S�sɤ��5kit��}�� #Z�LP��R�s[;Z�i��y�p2I�L��g�#����=�Ǯ5"�j�4��-��A#�ۺZ�/�fס�O?���V�����d� d�h��Uo)4Y�Cn?���p|Y@��Eq'(��u�3ͷ�;��mX��G��P�����H��gZ<�=r�m;.�Gz?^*�W�Η�}Jӌ�Mu�i�v�"��#_B�PRwE���s��r�q�"��M"����h����+�8V�dbb ��˥2�k�e���OكD�	�N���`\�|�N�e�5��U��÷A��$�
;��`:��k���{1��K�2����t��]�/fZ""DZ;R�p�<��ҵwI��j����|��-�;k<iׁ-����A�%�ċ^�}�:���/��A]v��A�u�G�ibk��!�mg���Y~6�A���+}a*E�$�����BC����ib�^��>�lȆ�����y�b*���\�{y�h��b���T���A0d���G�����0���t��d�Ox�*��H��\kw���O���π�Ą�S��C�|�&�k\��* y���L�FisC�|/��"1;��F^�>+)��ڷ�Iz�:SNٽ���S�0���P��N�s�Db:� ��=3O[�{��m[�@���}�g�C#.�ICDteF�L�o'��c��P�M�/�C�o2�o��&�xͰZ��(D{f���pҗ�]U�|Uۿ����_@��sK��h�'�]x���>�+��}U���¾9ڤ
����m�=�y���<���أ|cJ��
��/[� ��Yo3�Sĝ.����C7�0���$�b����ˈ�}�D���=0��p-���ҿ?^�\��șj8{��*8��=�6����o��<ؙxb��`�n�	\�\�>^�b a���WyrI�;���������X-1�|*a�}h
��$&�����n�cG��ɑc����^F �����
[nQ���l�?T�`䈚L����Յ�O�h��'e�Mل�.(,�6�.#��6��Ë�N$g��K����^y�sv|�1���0��ƈ�9xs�٣����1C��:��RK^wk������
X=_�p�JV�ia}��-�����H��<^>���Y�N�d�!Ls�G�ڏ���%��<��Mz���hs-.>:�!Y��AMl XoaA���"zyH�M�7$�.����2��D��li��D�_��HۼT����	�=�TL�Ѿ���K���tϸ�V�d2
hey�x[�3�*���Q�����j���^��g �8w�+����>��?2Q/����(���wݙ�89o��!� �,8� �i[�mcB_mQdT~����On��$�6��w⠤"C���f��H��e�)���N� F�@���e�[�1�f�#�iͷ���8!�?����Wf|�f���j67\|w��to*��^q�[��i���al����4�'W�!�����+47`��H���_���)Zlo.Z�_�!�lv߳g+��
Y�GA����F&Ctz-���R`*sT&���%g-�����- �	FC��L�ԗ,'n�[r��0R(?gL���*���	��vE��Q�ЂÍΰ���Q��ߧ� ]򟎹V$�d���'�{��J۔���.�t�E֑E�����2]���s
y�i��.��ҟP��C��b�92P�;Qx������1z�+��
Y�z,��-��?o�l��_t迊svM�UB�o����C�	���̒�����ڂ�-���}����bt�͊���0s�����<���q���a�����_�[9��&z��3�ȡ/��a�=zLV@�A)Y\��a?�ĝCk�i���¼J���q�2!�oz��N�P�).��k˗e�\��|� M�_D���`�c�P���s|�r��j��v�_�S��d��3��T��1�"�h�M��2w� ubݑ�S,�����C��c$o�@I�$�M,���H�s�%��?0�Q��xc����*L�1�^�o�a��w��>� ���u����
�o�X��j��F��^�G^qR�,�f���RQO�ӽJ����y��K��%8�0�̈́TYX���9uQI�4�!�~��Q�`Z���b+�И;k�kh8�{�b��2l�N�!�[��ޅ��k^W��?6DU�W����5j�p���m|1xd��=A����br��o��(�c��B��S�ҡ1_����&�P��
Z�K��$��6[z�e�uq�R�GA�����Ү܏�/~#�i�v��e�>;���H_k�BI��C����jz�]!
`F�;`����g~��i|������m�����:��#A��}G�Յy<5���� C�do7�T#j�ʎLp�����C�,j�UR�^I�ħ��x�܏6�%��Cz}�6�f&��s�31.ma@����XlK
E؎�����m>$��;T��<F�y��1m�	g�o��و��To.�}�`/�+��/j�|
mh㺖�С�I�!�eHiHN��9�8��vV�}���3�n�6�\���uS�&�������6�0�sL���N�1ܤ�X�������-}�|�׀�-}����*+� e�S�:Yu�d�9�h��bZ7V&,�<�/�p#�7-��_�kv����'ҕf��b�����b$�WSy�Vq��P�n7G��UoH{D����{�hT�`_�C�1Z�oU���x�rT�'ہcP� J $�,J��k�Q��	b�b��=���bn����G1 '�"QL�H9ͭ<o*�n^�«!�I~�r�*{S�X�h�p�;���m��� s��G�T��#�u�8�D<��ƿ��0�<���t�rp/,�PL�4�ZyV�˗�WG1Jؾ�H��HKS-��(�h��`>򜇗����L��B�����x��aJ�ǽ0�����Pb%q(*�(n_@,�a(�Dx#������h�4;i��E�Z�"֌�w�V
O�^>��`=��,dA�;Q�59�x��/�WP->��H�pJ�F���>QI�e�(r&Y!*��S�p�r�(���_������j������x���7l5�EW��.���������vԿ�����hޝ��_I'f�(�k����E���.+��OxM��%b9J{����%�g}'���$k{���u� ���(� oZ]f���%G���\�ܘ��iOt̲����2�s'�՟@t�L!t�g��թ�[��v����>����3�on4>������� �K�T�CL�^B�s}S�H�������D��F�09�%��~�O���3�w]dz�Qfhuq�2��ʲ�joҝY�G�ǎ2�*���6}���BK]K�[�����u����qX����V5���S6"��z����~���C�E��{R�	����D�Ʈ�,�����_�kH@��ٚa��HX�f\Eb�:|�=CsG���q�+q�@|Qȅ�O���q?�S|�X�Q�?@$ ���{=����/�R��'qP4��泂�z��/J��n/՟���~���J-�o-4J	��J��_��}���&dM�y�`�! NԔ4Fr��S�����vU�n{d�?��G�)�5&S\���ʾ�+��𷲅���X`Mr�)a��+�h|8x)�芨_�ʷ@uZk<�~�8���&h=�7���NY��;~���еWN�b���4@<5�:�Pu<�f φ�/Yu�O����#*nx���0��{�d�x��9���Hא���R#{i�
�'��eKɯ�!G��!Y��T�F[
�:�z�GL�`F��`�$��j�y�����hY��bI��uM���6�I2;u�=�S��C>>�|0!��"���!��gǋ�؋���hYO�.�%:�:;3��+N��W,����UP�������P������i�{ƕ�s.��r>Yf�0ʋn�HC[�&�B;i���tRb�M��NzI�4q��_w	Yx<>������š�y��ϲ�ILǧ��*�������[s���NEg*���+c��(��d'l�(D�)�\}�c��3�f�52�>����E��J ȱ��jS}"bn&  ���S8u��(�G���6ܟ$]Wo����R0��_���hߌ���`U��ϰ  _Q��/�3�.�o�K�Tvi]�/?$��/`���>�`ut�oHa��d�h8&�?���;J�X��;렵RK
r��m�c�{*h�~}��O	�e�x)xpCSi�r�>�<-0�P�}��$�'�=yR�W�mv\u��e���f0�=٢�Q9g�1��52w�>�[��N���tx�[�@ �H�O8�;M3Z��("�6�����V�5|Q�2�F�
��I��7�g���!WDrvxA�0b�ޭA�#e �&�.K�r����j��y�<T�E��|�ֱ5s��=ym����OyZ�2����黀��ߌ�ؐ�8/�!� .5�iJ��u�2��c��缯�]\+�;2���������zm�5�t�J+�)�6�e�$��-�&j���oOM%l���D�K�'�s�|0�<����h����2��a�eϡK�һ�uI���
���(+�Ug����������������o��{=sL_1-X��J�!~Yehs����R�7�����b��l�ra��s��������R^0���I4��+i��s
�td�̦2��=�iv[��5�4U�P�i�򽯐�,�?���wV�s���e��@5�ǛK���4ڧ$7%�~�����&+	��;��/���&��a� ζ�h��	G㑆f��s��J�֋�j�xx�ؕD:D�a�+iDX`���!�&�:P�m���j��"\S��,a�㱗5�h���d����ꟷ�UuxSX�q�!Ճj*
7�*���~�����g��re����q3_��Pڵ��uE'�>�Խ{�ҝW�O{t������7���a��C�պ�v�Dyߛ��r�Ͻ�	3_1h?4_�j����:��������&�m���Z.�.� ���0xX1��?�9ۜ�$�+�\QI�'��c|�io��X��#}�R>�/7�.���$,�.�e��OL1tTS11�N��Ζj}9ت�b����U�dq*�)��U���ݲ���g��v�P��m1G�"��E�#�Wȉ�:bS���̿R[�屲�;���uWE-f3��e�d����i�>}��ITT�X�w	"���E��΃�~~�ZY'�Hl�����y�R>��u�֞�֋g��pI��?Q �S��<�RIޝv�P-�h��_�A�����D��n�߃����#���
)KfhM��V��>8 �R���(�A'7و��[�)�����6�L\����	����P)c��+��� �l[��8��ޔ�ϫ�hW1c���T�m�$��M�2rϱX��r�K��w�,��*�d��6J�{`���h�
s��|6	{ ��k�nŨ���H�� �Yt��/�� �y�������W���X�el���D��'O��[b&ٶ�I�����3��p�1�S�P�c�	�N���r��1²!́��V.�?p�s*i����e������6nSM�\瀠�,�9�<��K�����H�u�A��Ym(>`�.��-��L(�K]���ލW�5Np��-e���-���5�,Q��.�l����SX��RQQ����I\��X���(;�U,l#��m�P���?c�`"u`�r�H��*�~G A�Hܦ�鲺*���?�Q�)a�� �h#��] �"g��ُ�&��CE5�Ԑl�M��ҝhC��n�6}+�]ǋ����8����~ah����-P����Y�i��Q0ϞA*rz=V�WWY�k�5c��W���/l��X�or���s���\z�,5�m��0&��N������S٪(��-�/7r�2c6��Ǜ@k ��ڴ���Q\?���j?�����x����|/�޲ޕ|���_75 �T���{�	�ْ~���<;Ն�o�Sd��l�Uy~�:�f�S��Fu(�!�"�E��B������QE�l����� _\�u�����X��Y�C�p��Q�\���F=�I=OS	Lw�S�*�� 6��&e�`��H=�q�9�"�ݱ)o������8;�Zd�������!�jP��K��[�*bn��d{�c#^������D�Ԇ
`���*��o��n!C���OV D,�����ܖ,[����,C�ewx�sbi��' ��+<���{�z�of̡H}�ş�BJ�苑=2c����q1Yj}��iy���	�s�2�'���V�\2*H��^�V�vT'�)�}alKP���Kf��|��^�$K�8M�=��l����P.�M�5���N^���W�SE���T�T���!�Y�E��������tKW��!���.u�QR��&�4�x��aƌ�Z���FeeS�����q=�A���8����2�6�О �ޜ�/A�[�OJI%�+h���Ӱ��M�W�fHurE���d���V���?�,��� ������<O��Ë}��'�<+�qE|�A�s��K�xs><w�15�׀���T�u�l�2n#cޡ��PVZY�O��s����`W�;x'�?��Y8-��������	1ګ�o�ĸdT$ٻ�  
42�ߚ�$�[��-6{��H�C'��,5*�~y+ �$��Q��N��4�rN)bTaF&&�������7[yѰ���^��w"�&����=VdШm�S�������g&פkt��.��L��]�V3���,knm1V��J)�(��t,�������;�)����N�d���KnU�#��E�a�>&I�seg��3�Qu �o�D�%"5�),�Mz�٭��%�r���ʄ�h`�#�_�oX�����A'��&2��p��הQ�;�(�Q�B,�����B1��~/����_�[~pjP�-�?�㘜�4�dwG�.cl`�nU+�� �������v��"��4�0y u�L�I�c1�Ӏ�P�yeһ��=�� r�LT=�Օ�􆒠�X�O0�b�>C�����+i��V�j�}?��\�!ҙw�S�Rwk����QO��Q�����Y���Jr�Y׮�,^�C#�d���\����"HM���b�vw=|zkA�
�=mj��w�]vۖ�z�iq�66�����w�`���� \#u8~$�ޣ'�4�_�z`�{�n��S.���qb��-��ȧń�C����s��tJ���-'���΁H�|���� 7�QiO�p��y\�J�;-��*ン��^�qwv �X.�'����H�g�;���9���jO�����@�I�?P6�EZ�עM��M�0�Z��YiQ��d��0%�c��У̰�%�yn���L���.Vb7/��A�<����J��l��d�l&*��VX�~�xz��TR��|��ȵ������F�D,�/@���F�t(
d�_L\�5����VE.�n���]_)\�"vh�/�羽h���\�}���2�GHQ�n*
��?��T��"�u��a�@��1���w�b���|��QT!��b�U�'.č�N1��	�k�Ż�/}ɱ�t���&�����޶ў��+��W#����(��v���^Z�(`��|�Z3N~L��z����4oP���G�Zc�^�f5�#=�V 5^�*sS�6����k���2UAp=&�Hc~@��E�C��6�F��4����i��K�-q����]�����F�EZ�]����*U�D�@]�ED��D��8�Y��������]�L�DE�fKga�E�0�M	 �Hʮ��=�4�}��͋�t��:P�m]^��ȯ.;D���^u��~����Q[�HX�����|a���
�x ���3UѦ{呒��)�(�1l�VV�M��8G��}��?�o܂�ц� ��uz�\l �UN4�d�wx�G��w�e��܀a�P��^G]�R��O���g�4�zC���_�bF�����_�q(pR�\7�9�o�h���%������4�K�2`�z�iN��}p;�]	��a��WX{<޸CtUO�"@��Lc~��+mϛ�8����DFii�L�$�xR��z+�<�����Q���g�����_;/�z�V�%Ϣ���ͣ󼙰�!|k�A;p�W_�$_<t=�s���n���%�c�x쯳'�'x�� ,R-���0/#�&ߌ�Np_��!�Z�Y�R�p��u�e�W�%7�3W���������S�Z��k�Lsf���%�F�x}�a:���lu{�vB�������rx6��5�>.��\^��.tO��6aV�S��x��Y��Y/�E���/^D¾��j����g��P���O�D�'�����"Z�ߠ��؈F�O $�yO��(%6Ys���^������@����~/���������!�Y�]��Ho�ÙM����M��F+���cى*(7v�υ����J��+�|i��Or*���U)�(7�G�&�~�=��8|�+Qz�8�f���I�n�}60q����~	MYB��+����sp$��4C`9��x��?ǂi<̦���y��܅ЉV>T�鎀�Vz�ڋ���mx���	�=�<n��$N*�:#J�B��	Q�ǩG�l끙��G��7�f=��q!?���rݨ�2iw�׽�m�����K"$ժ�����Maܹ����l�1N�R���T�N�N,��#n�4�Y�j�>(�HBb#>�!

={6�4�5���iy��M�ky˙�+��O6��wE�_7(�:*�Y�)^ql���w��&du���*B��F�Z8�8T����},��"҇�hX�2�ԶRs#���u)Z^�uǧ�)��R�=DޱL�LϪ�.s\r��s-�=�>!\*r��g0	>۬�OѤH�0�2��
V:�&KV��&%�!$�ķpS���;B2xHlJ�K�ºdK��n8VMX�'�s�+����C�J��r�Y�̘����*?wl��-\��E7�;U�	�^-��)0���|�V�0��t1�!�純[:u��C��%7щ_[��jj�murJ���(ZwZ$U��U�2�{�yn7��m$������jjQ� #�J���(2/4�xA�zhn����J~���z�h�	f��P>։ʄN���ѪbDۣf �&#@t= �Hh9"��������~C���@g
�_�#tC\��ȣ�5q#�<爈�����#%V�ı&����0��`�.�f�B}ԟ�����%T������� D�� tx��߫mh����6ꨋyi�8��P?z��K�R
�w���p_�P�1�h�@�z`��\�1��p���)6ĸU�8����]�(����r��-�/ ��<Xt��nL�<�'�*K�pCk�������Psz��v�IP���] {:�|;���e�>������Sܪ�`���!`��A���z��jy��pmo���������4�r����w*Nj�̧��v���$��.9��x��Z���g�+N���jh
�̢�����,w,o�-E��4Zf�)�J�Z},�^��)�֖��4�_7I��ź0�~X���N��*�0Jg�
�����j���I}�m*-�ݗS枊��e�b@(�t��	�<��`C�� 6b��(%A��;,_���f3w�id�L�H�	�`M����[��;u%6�(�'"��6�Z��5��F�lX�]j8���qK�a��q4<���W�j-[{�
^]��kR>�k{����|�g�\������Bc;<%�L�cx {�I]r�-t<i��@��\z�Lfg8-	�z�t�7�j�n�{��B4���n��:�T$y�0��7S����|��Ğo�D㟨H����PA����3�Pd�&#Z~��A�c4���y�,�:Zm�#�u$ʄ��%+u1��P�6חi���k��v�Z甴�H� !��*,��r9���1�qvD�n�Þn5���~�N�\఩��P��R���2�J���w���?�]�7��$X6��d:L�
6�u`Ά���h'�����g������'�x�y)M��F���f����B�ģɍ��b2�u�U��4D��O��㰚Ci�Y(���Jo��g�|a�ջ5�J�Mӏ�~�R���P5)N��I�����J�A͹��J���f��E��h+Nu�6�3{;���h�����m5W���'2{�i/��e���u�ݞn�����bk�)2wr������r�;;���m��,y3��-�������3������Rg��?N�< C@
{I*�Y��u��-92Yy��%s�|����M@�e'��0�}��D��W�(��Nӻ1;J/C�'�M�]uU���`�n�`��Eh�:�����o���_Ӏ��s��q�0�k��FtR}?$��N�f&C��%�4v�r�gQ�T�k��X6U��!���:���"ݝ��ο�U�L�hҝ�ŋ��M��2L���t�q'��p�P��K�v���ȿ^$ ����sB�e*~ۓ������m�m�Y���%�#f�I��?�cz�����)ݾj�_���_�!�o�N��$ɤߓ<>JIalt6F��9�!М�#|�Jd��Y:ː���a���}�� ي޷��Mv��Kz{a$��4q���=�W�����SpN�d�2S% ��Oqɷ2�t5�QO��GU�������=HU_��`�{Jc:C��iӡq�(�����d���L��c����A������|9�O�q_5I����^=��|��$�f'\8ìDt��kdhW9�"7`.h�=����ά�`jN{���R��Q��?7�EI�|Ӷ�I8`�ֆ!o-�I�����_f� ;k��>�O{g�:�=<Ɩ��V�	�Q�I��GϩPI��A� ���'m�����R����$|!Z{�ͧ+���� ޞFÌ���n�ƴ���|��/F��I��~�:9.�*g��$ P)_����bP���M�sf���=B�I��dA�Ɇ9�=㤨��X����9�x-��m͵>y��_�a矒\V�k�������ȴߌ�uv�/+tx���,��8д�=;/�R�GL��I:��R�4�A�� �A����U���&t�Ʒ
G�6��B3��mx�tD�A~�N4��ݶska�qaӾ��Έ���t8rTt���h�l<�L
*�Tc?���-
�1�����ʥ�n��@6�R�����+�������O*)�ԧ=���|֮��= ����XC�|(J�6�!$��0�SL���YE�.��|�靡+>}�U�q��oo��H�*�s����a�����.'h����W���*����s�࿗P��pJS�	Ի"
^t��p��D�C<X��3II�#^�^PH�ܛɋ��r��p�~��zW�B9+t����������!�Y�|T���F�B�w��U&	O̠�m�\����"���&��	k�$v=�A7������L>��S��Ja�	�`o�g/�2|(�^���0������<B\���!l�W!�7��H������ֵyՏ �MKX�T͓���H�Oٶ?�a�t;�zK#Pq�v�#>�d�G��SH]��(��n2p��\x1�����0Y��,��wC� &;E�fƅ{�$�������0�wh��GE�݃rʺC�Lsm��r��a@��rֻU�H|�կ[�P˖�_� _D�N�)1��z]��[Ui����� ���h#�o{,�z���7}�-�ηj~�]Ju��o6��cRt���# E>z��Iu,��q]�����)}��lY'���c��|mb�瞌��B�ߤfs�z�6E's'��ZTo,j#��3-͚z�F���y�R5��E$YX�:��W�Y�n��[ZR�g��h�0�7�DR#�\<Nq�~n����@z?��^e����-�`Wktͨ��D(F�%FL��d]�xB���ڔ@P: 7�������C��0��u�����.��OH8��	�`n0�K4�$'�E�\^5]��[�"��Q!DU�e��Ds/��l3��0+5��B�����fm��Mxl�#���) �H��z	�pg|��	�;�J~��̷�Y���gt��ޞ8p�Ja]������zpZ1�b#�z>��7f�A]�P1@��c?��;Թ������Z��{/�Q��nQ$"���=���+d|��ww��V<��Xo�j��s+m:��{���J��W� Bh�_���E�'�G7 ������r����#�=������F�(���fs3��9�kB����J��;��"5_O�m�\F4�q�́��i�m��0����[ۏ��D�&9�`����t!>�2U1aP'xf\9�tQ���K�{�6b�,�8a���'0#,�8-բ�xi�zC���s �t�Z�R�̙�b�M���)i�?t���f �[��tB�x�|�*��\�<&
�:멪�)h \����S�m	di��H��&�翝��9{E&�y"��!�'�����+4�9�z�N��Z��t���S� �@4���.لl0B����.(A��P�b	%sy��9EeVZI��+�-�� �=.?�=�jPO���	c�J1��?E�~#c�����S��9YY&������lN��Oq�z�o�X�Ɛ����m����h'�����l�H��q~+�G�9�n�r�[��̂�}h�[<`+�t��T��r�I��.L��!9*^ �����˷��l}����|l�[�t0�p*A�2�i�o�aV�ҀD��һ�*�B�o��Kl�v� ������Y��ʉ�ʚ ������NG����Mhi�1�t�S~I�iE�ԗ����Y�={����z�k<{�����,Dj��d�w-�1Q7Eq�勷9ӵ\j�^p{��P3�+(��:�/�A��eF��rWN��jࠦY����˫.�r�Xz"�
$[W���X�ڍ���`�A�����lc<ݛ+�9��uq�|&�B4�2r�D��ͥ��S�G��^�d{tT�C�2��{	VD�@��}.��� ��Q�������:�m�g�H������p(i8y�BB�h>�r��<����-��>�>���gwRL�����{bf�>rfN�|䩪�ݮ<��2�}B'o���9�v�@.Ϣ��p|�*X�c����8IN�-���u�������-����ZJ�97�)�Ӥ�,�������=Q$ح0�����M
���gQ�~y�����a.O��Ho����s�/!�9�:f�_�G+��=gě�5� 7�[h�1"A1���3W��='��=�߅,���I�!G�d^:��K�'��פ��Z���[Ӝ�D�"z�M�qD��H��^�>��֩�Qu��~lj�i�C�#��YB����S���^~��d���L
�X�ي:�X��LM-n:�(��ݘ�]K��ai��e����g���+r�B:�Z�Cׄ7^5���GN�z�㹦��#���)��T�a'�5L2�H��@N�Xl��>�$����M��H�5�f����Qu��D�
�iu���
f!��v�\��������+C*PJ�}�3t�a�]`F&l�����^�OfC#�W��Bn�J�o
�j���,C���0P�'6o�_�� ��$�&*���q4�� Wc`uX���LЉ��u�Z���T�Ǝ-�AC�ÛW���b��I�`��[�%�c�Y���� �������)\���^�So[Cߑ&%�96[,��gtx}ӷ[��F�(�`���
��J�|Ra��jN�=����I��W�B5�3��+g��k"��A	���H��xn������2��{�P9�bH�K9�ҁ�P(�,�8щ�#9��4;\?�#��i8κ/f�C�RF�c������%*��0쿽������ꦩ/"2|��˪�T�N.ƙH���/����^��i�A]�5TJt\�5�>�w-p�_��o{������3H���&��!�(��sew�N��E��bc�A3Jq�0L��4���u_���` ��Y�Rp~�䝥`�b���?Q(�D�+�8�SQ��u�Hl��}�rPDg)Kb���	�oDX������$��'J��/ne�^���A������;�͏^M�F~��V!ʨ��R�ʩۨ��)��D҉dHT`c���N9���|�غ���I�5�D��f��/�)d�0�wM��^f����7B�;�A4j�����R��h*ͯ2���1��/����	�����6��mf=��~\������x���0�?j����,q��~ڔ�A��#����.��sh��G#��Ј�<˟������@��r�q����lأ�0.q�@�2��h���������z��%G�T	|y�I�ҳ޼�|ZGtP,0���DU�C��X�\Pkf�&N�1؂�U����z�[8�b�K ��~X�4��.�Q�y�>ߜVTS�:��I���/�8Њ�=�H@Vqf&�m����z�Ý[#�$��˚�F��Ȼ������5L]R"4E�%�T��Y�My���Q8L[&u���x:uu�*�2k��#��<.A }g^xpja�39-�d�K@�O�Ǜc+X �Z*#��(��L�_Ջ��@�����Ї���B�NgԐH�l��� 6��n�F�:�*.o��=�M��ë%�Z����	�~J&|S�X덉�?}�ibv��'yv�J*h��TYA�[��~�@���q�2+3�tp��6�
�uXx����;8��4�x^���O���GfR{K����pV�^^�/��^~�m�΄���AS�����_�k�|���H7a�\�LPfd�wi$w*�)��)���/0|k����tG��X����q?���|Oo����X�J3ގFlJhV�6�s�}�ݷ��h�Ç �8<� bjs0���z�I��3>Rܫ|�cᩱ}�U?`K(B��	��H�D�cXF7
�-�s�X;V�RS�S�x�
И.̟AB0_Y侮�l��������r=�Z�'�rE,�|�,�
)i��c�'!�aq>$D,�=\��¬J�9���J�з���
�1�'V� k�D�q*��mh��R
����1�kE�s=GJ:K̞����~FI�4�va��1�P#�6T������4 �W^X6҅޶�獫8��G��B>��ۑ���\��9^F�p����ќ��JRB��F�>�PȬ^c��8��|�i
�>���z?Ö2���t�3�YX<��C�#�S��j+�>qH7k�Mi�a�ݖ�c��.��;,�G_6O�v2T�	X�T�����J�����I�DC={iU�lu=��-&Sӵg���W�U$�S'O�H���ZLH�H��0��1�}7���k%��F ���&�r�Z�ܚt�8$E���;��B���T�_Q�-��,����8b�� џO̬�8쀹�.�tt����iP$���b����m��P~�O-T�`B��M�Mow�[��Ai���x��k���9s��_=�8� ��˯5˴���,�NUR��n�"Ի�yM��#~.����i�lh�J3N"h�gU��ͱ�Sq.�3O`�n`��ehA#�b��m�A:��ф����W#�@����΃��X))���/=�n��B��h��^�m,z��)�Q�*p��/����	�$$e�[I�%�5�0l�*I)�i��ݙ�����e���Ӫ���>#��_SY�o��W���d�&{J�_*����!��^1����3��\|���-��_f����l�U�(�qI����ST* ��,�fX�TI|w0���}r�?�%,���Ѱ[~f����(h�Q �^|������\����P���W��5�U�]�&��8����7��z���
�ʕo,�/�Ar*_p$�0�-o4�_�{wޘ��)'� �d:���/xI<��v�-g12�ތ�2��7spY@'�\CL���s��Գ�usݶ��K>F�H[J�\���������m�����c�j਑�#⇊$J��P����7q��=7�Г����gJ/�Ե!*Xk>i���c�}�z ��{Kr?���&��R�x��fQ��m�|��+э�vv	Cp�z��]5��_Q��)4-�|�����U~�ǡ�j�ͫ[�U�H��#y�;�I����U�����8�����?�=� 8��D���-)Z�c�2��.��P��ܺ@���7�dT��Sgf�QKzy��ffoh��VE�N��垘�66���j��e�r$�5q����C�ܧ�5g�	&��n���_�=,\
|��-�ǷSA0c��Kv�8[������X`	<:����7^��5�������qT�0v���[^���%*�� /K��I�u��<�Jb-1���4��aa5so�A�k[�5眉ҟ�;F�ϛ����W��M|h�ʈ�\]D��c��(��8H���n�)*��H�
��1�$��*���ThX_4�aU�A�ϗ �lWC���,��s�Y���U�?p	#�ѫ?0�D���(�Mٌ�smܹ?C���rlO��=�m�K���S��3ch�ޜ�����[w�;�\�����9G�h��m���5�y�[MYu�1Rԭ)_�V�c���ie���y�۷��Ĭ !9`>�m�N�߼�E�|:�F�^K ��i��F�´kT���9c{�31��DEv��6�����Tu�:�YC����ǈ��b㘽����֐̤n��lVy�&��O���+1�E/���h�����$�+/;�s��.-BF�J>ߪvA"�ȿC��	���Õ<YP_w�-P������R�^���j�#�o/1)>G�^U��M�p_o��ZZ[�n�0�a�g���}�r��u�$x๭��LO�{��H�m������j0��U8�"Hݦɩa{OB'jҺ�*G���Y+,�{h���`�
��k�"�` czN�
�d����1�e�맇��M���ӠAߕw�K�܇���]��⠼�C�=�jܥ̩7��}����R+���'����[�B2��ң@C����W}-�浥�]�a��?�3��,�𹇚�tT����󇩽G?�PO,7���^����a�q�^L)��tH���p�g�5�Ws��2�����c�t.R���CoZ�ĕ�߷��&ߋ�J�ƥ?d��WZx2��ot��R�$~3���T�Z��CF�kr���OA���:! ɨ�)mB�
Y�
x�O� �������MF����a7���Z�S�uNM �g�������A��n�Dj��=�fw$�.�k&p��GӁL��(x�.$9�y��:��A����y&��b� ���%�����{*�I1�������r_��<�:��@#�Q�W��*�p��A�<(��o�d����sM�C�s o���� N��u���A���Zb�Q.۱v�eм�o��(w&�����@�+m,��@�L~�]�&)��$��l C�Z>/�\�!���$,t}��9��?�����@	�u��|�U��>�-���9�3�E�w<�!�|�O ��e��Q�#�����=M���0�Js5�`P�}����.�*�&�x��%����)���#Ah�������B����q��g��/�ɰ�Y��Vӻ����m~�he�Cԉtm�U��\��o�Z��Q1�%��0�Z���F��r�j�Lr���s;2p���#���?�a�("AlV��h�^MWK7]��)�r�k�TRx�<ٞen�_+k�8J^�׭�l�؉Y"6-��@�D�}���h�x{$ϗnd�4�նOvro�lL���^&d-:��|����
q��6��G��yU�c���Ƈ�N����n��1�:�D#�JS��Wi,9w�
y��F�����O4�O����+����e��&w�06mL�}4���a��b�vi�F
���ՏBnH��4޳���VА%��RE�ty�H���)�f�HYK�y���%Q;��C
�7?�������K͊���u��OM0��W�I�\P��+�f@3���O�����.|��V�%���o	XR�u\\�� &UC�(@&v]O���O�9g�BHBъwW�����m�h;ψ�g�֞�����u7!�{yh��Q�3L��;�!{E��K1�rө%< �>I�&��2٧�^�����=Lߧ~#=���XG��A��Yqj5g�E�ݪ]gl����n�'��!ԛ˻E�ֈ�7r��|܃]�,l �a�oXy&�_w�ߝW�E��?M��a��<�_>�Kp5�����X�6�'� �Ì9�0���Z�t�p���X�!w�5���=~8^?��!�8&!lct7Y�T��J��B;I� �'SʫAL�&Y��)�]�0ē����YS�� Sl%�a�@��VF�vI�9|��;!	�ы)�7	h��0!{�0����1N#z�}��C[8I�y���4�l�G���Es��߻��0�?���Jݷ%�𐭕$ ]�W�&B�G1��	BB6�ǻ h��t�g�j�f�Hչ���Tx���, ��c���UK���]�x�:���{N�C����E9/*��	{��� �U����Ob��qS��B��]��@C5+�i������'W�	�0���XjN�w
i�-�X���gÖӘ8cTi��}G�#�@�~��z�xGg+�_��!�����;��D��/:��F�!��8�"o'J`���&U�'y�$w�J������Z �����d}�����-�MS���5+ՙ��ʏ���u#׉�M[��U�j�VU�s�A/���F�$*��'7�:���A&��Uӗ-k���9�~��\�>��5���^�f=�ֹd�O�\ .F`��q��_��oG�UC��u�G��Il�g̟WwYQM���3E����.ʕ�/�ޟL*@�M꼝��H�+����pB�',��JLP�I󜷤#&��VRq�&����+�����voc�e���DR��9�T	j�ԋ,??��an�j,Jӹ�B�П��X
�-�f��2�0��Psn�9zn���~4�آ�>�;�#�n}�&�0����oH4�-�n��T�!C�`ԭY��W�A� ����tQf�S��$�Ŋ6�g�scݿN/m��G���}�����p�￑*l�.���?�t"Q�:�L"䤮0yCO���ɦ:c��G�� �:p�nC9�K1F'~
���y��K1�!�[�?T��� ���5���?Gp���U�9�)�B�M�;�]�m�uCFg#W��m����_�⽸�i���ڌ1Q�=,�E}���	��AK2<U;�5��V�f�9�fp��l���M���M�Bl��F�Nȉ!�XY�Д{��o�#H�!Z�wi�#�7��v<M��yD,����"k���la��,�)�NCX>0�'�Jl�~ԓ��l8@:6}����]EQ{m+�ϭG��z[�X���V�����AS�' �����0My���7�L��8�S ��L�7�0"���6y����n%=^<�*�\d$a�	YN��Q�J�}m`WFZ?��®jW�@�{�Ո>T�T�����uy�_����]�����;�{�'!�{�����(0�9�p����9E��.cS�G����]}�	&�⺘v�p/�"D�M<:h�>��?OfH���.�t0�F�����F��9B/��]0�ܺI�J"�V�GtC`�7�JWM�u�M��m!��-*� J�1�I>�ǈλ�0�F�Vw�2<ǡP�ʳYK���Y'L}��L���t�+r5}B#� C����z(+�}f���-���N���H��5&I�4�*����>��{:
��	�H�/F�~��5#�s������!��HB�,IMRQ+teA���<P�7N&��J�3e%)���������L���v���/2��E|�2��kZ�w`�6��ogl�uohR�\�f�=��7smL�׀�J�6��3�C���{��wYNǗ�M�������oߎ������K�
�)7���90�&�O��s��S
�۲鄚�������`
�Ի]z�ЫSo��Z�xe�����Tg�9�
�lj���h�B��~�~�4$�m�:U2Q�e?/��ڀ���eՃx���Б+��0H��������1���X=x9
�Jx?�� �iG�(��!�J#���y�B������"��!�ޝi����4m�����7��%��$�t��#,�a��A��Ӯ��K�У��F��؛p�VxTq�L��&]w�i@��3��p�3F@���<ε�I��'/�ˏ=�b�;/gѯg$���F>Ѿ8ř���kv6��(�<h噜,���>�¬_ �����J�� ڶAZvT�6�koK$�\���17zw�SW����I@p�H�/�A�B��=�(}�;D�j��7�ޗ�ݗx�O9R��V�}��\N�����X�o
�5� �Z��=u���._&Zg4S�{��6t�'�5���ª�`Rk��)��ت�[����9Կƀ=�}�j)70��*L�T@F{W��C�\���_G^�Yc���B����SvF���A�&������r�b-5����j�X�6fa�Bf�W�6Z�jQ�-��{C.[��FD2'����ܢ_:g������d|�Xa4N��G��y�b�\z�dP�I�o,�.�֠ $��0�J�zҖ����B��+�y<p���3�����ŅT4Ȍ�dRH��6n&�jF*�OHq�U�v�����|Fab2ms�*
�:�j���o5*pu�M4OZ��ئPo��^�S�I�5�(7���%�T08�A
���u��N8^S���3R��� �������]0��]�G���-���M �C(>M�a$Sr}���[m>�LF���(?�|
�+�n p|�|dI�N�G��U5�}T}���V�F 
��^�!? +�5�X�Q����@���;ڥoZT���A��?���´1[�s]��Y�O�M|/�&y|���Q���M�Z6�٬9N���#�@]wr���w����Uf%P�Q��R�j�#/.a���F�n��~��kK�+0��
�̱�@� [H�~�����̅��xoQt�*t��T��/3B5��&&�s���m� 6�;���қ3x:�q�Y4.�.e�Ts�=ϰ��B�[�(����8����q��;3�ퟱ��p��9o?�ȀI)���*4�H� ����ޅ�[� ��\�Ѿ�L��a{�v�G�YU�E�͇s���o��EI�A�3�m[vzҁ�tz��E�=�C�m��C��@�5_/�p�t�4����27�SE�
�`1�x<hs�Z��3Z��d0�ORD	�\W��.p�m�� +�����o<������ĨQ�s�o]YU`����yO������џNʐ�T��$�{�Sԟ}ǥ?<	����9h���Æ������j�as�@l"�����sDS�lSH(��
��LD�Xi�Tҹ3�-�bǱ'i�	���T$JA�I������ДK�?Ұ�߀p��K�/��oʡ�.%�V���$Fr�Os����=�TT�م6�5`B�H�k�iw�%�tԿ\��˪�Z�|lHm_�&Ҧ�����7.+�+��SnQ�}�E�����y�!�Bf�ؽ���(8��>C�����LT�N�K����_���d��wӈ3�R�-��k� �HW��13*�w�x������,�)�u�ښ�uwX����O���I&�ՎyV!��P���&+�ʂ\̩Mr���È.��g�u'?�ܹL��Ƈ|Pa�z���d��j�y���-�aB�4�1at�~���]����Gw) �ʇ�ʚ�z�ub�����v���"����P�cy�Җq�X�:��ɦS����V^V�E�*�DX�s'���?e����4qhE�@=�OV�Wָ�8r��weWn@i�4�C�|�+���[5#��-�P�*�� �T����'}Ic��I���q��̾3<��sR[Q+>�ó_�y�Y|s��:����P��g�:���g��tAo��SM����a�y�S�3K��]ͱ��KA�@�$����r������`�7v�\���+�^W������<W� ��5*��3��������Fn� ���D4bE���v�����p=�� >Io�JU[hm�h��c3�*"���=Au�Nڙ�t�n�O��¤h�����u��\3r����M�aY20����'�J��2�N��F��$�nm�(��o��{�D�R��e�%�T�Ʊb����l�M�#�oY�Z���X�\�R�w���T��h��byV�uJu��n���7�:��3d�ű��6o�F�{��Cg2V0,΍u3�����.cJ�}��lTJg⽼��ŲaDL֠��~7���"��|�*J�+�����i�(�cKOB�ly�|�]*�W-R�H0n�J��~�Zh[�ܝ��[�]<��9Y�d\�9G �>^S	R�W�-$�+�Sɔ�7�����Mz��>|�_O�0D'�o�2V�9K;Q�ɌU��Ȇ�o�ch�Б�����q�;-:'E.ֈ��ꍶ ��h��Y�+����G970�@����HFS���4�����b���G�V�͎���w��6�F/pR��T*5���p-��]��(k4��9����6�T�ﴑ��!��-�5��WJP������
3'���ވF�o���)����φ��E�ԚJM��yp0����9٤:�v�CI'^�����~e��O�:f*�����9���x�T�@ã�*���"6��[kG�O��,�G����.���;�g~�.Èk`㪛�rlw`�~�It��2��})!����'-:����Z�0����~�2��f�8���h�D���ޱ�����A!�1��L�����^����E��r�N������Ux��I��!�3Ji��?�T)��������bŸ5)�ب;,���b�;w�z��U�b�Z)�/bţ&������
���$��x�<�ap���24�&��o���"P�	��&�8���n�����xx�Y0P(�Ţ5m�ZfqkϥB��M�j����HW!JzN77���+�l�f���Z��kE,?yg>2(s����=�OЋ��?���f`t�-�g��o�G<'҂�;�p^g��SV�'���Hn���n�У�(�j�A�IL>���>-wC��7�f��j�=�7k�(���ٰ���*ZGq6�|6��-]�i���-K("t�]�&{��ŀ�.���i�2�B/��3�
�զ{��x�.ϙ̛}1L3��nG�ɢzɪ�2B o����	%6�A�/�@���wϸ��g�wS� ��-�d�L�&�����z��\�.{@w-EO���O{�Gߘ�^����u �B"ֺ'��d!�_��vce�ͭ#�v#4Cr�lbe��<9�����j�n��	g���A��t(Y�D$Rbh��������B0��r�5v/�v�-�y�)_���-YE��"t���ڑ���gpg��	q��wqۥf;n�h1Hr�h!�'��:�ϖX�;���<���� a3c����6f����6�t��b�;��~�l:˷.��;M��+�>a�ʇ�T1���_<�:��SO�S�f���Nr`o{t�D?3\�,�N�|�θ�fӜ�� $[c�	��6�
�J��'W��F6g>\F)Hv�1�6}�d��' �b&�ey��W���Z�п��&3����ǁ����˜���8Z.%ɕ�!0��p��%hG��>d��ˎ����W��ş��5�X�`qL��ZN��A�tV�ۙ]�J��-4	\�3S9j/��_�*��+����|VA���>�����iŒ����T%�Y!���}&��Q
W��*�1Q�r��
��aZd�Z���-�M��)Qƅ����"���pl.����� �T�< �No����h9~��c�ꖃh䵊j��-�ST3/��t\b�9�d;moI���A]�Q�Q�T���2ҮO�t�#��!/�׬�KA釧�ky]�>��y�Wn�ZB͜�-����|9a ��>� w)u`I��GN�1 �c��]�x�-o|r>�{�'),|���"J��;�?F��4!�`35�գ��$=?#�hH��C�n�2�@����Z�J�t�1�B���>�$�9i7�<(�a�q|���}��X���_�ա�u#=�K�]��Ҧz!Ȥ�./Ş���:���k�S���^��.k�=}:>�$�ص�y!��ȫظ���3&���N�T�����o@�6�J`����-r3A�h��@|�.�A������՗�4�u�쿼��)�_��,TR����2�s5�����~68�-}By��W�b_��5gLh�%�i��Il���q�����iDt�{{H���   ܃��2��\���9LفzZ��P��ah��㵵 �d���-����Rc3�N�m��Z����j��u�l?�ԗ��w�#��?ϓ�LZ.�0�?�C�hF�{�{f��d]-Í��ݺ�s���U*�Y�J!��G[��fȦ��������?Ö5����6*Z��ƶ����~O�t$�0~�����>�,��a���4��v��"2(>�||��L��xT #�K��_8,P�����r��N��j9��d�+�&�#�m�'�K�+i?t��L{�c�EP�K~�]��[4uu0�,��7P~����Z��ӈ�ڍ���C�J�F�%Z$i.tϭ�:(�6��k��t^��H�x٤|�n�
�!N�5v[	���J���͍��otJ�Q��Y��I���R�b�8 ���8/��~hui��aS�oA��Fq�����Fэ���g����#�q�1�,��w�0J�1/��Cvd�F��/�oV�,�%�=���@�M���=����5-�N��%�A� �y�K���z�_ �)͚[)nQ<L��&����>��ƃ��;������5\P�F���)�K�.F���@���_|�1��DY����'^�D�E�g}� ��ѯyAFw��R�J�#9�W����@BX�K�g�S��S�#7�p+!#4�t�/9r�o*satV��S���q�U;S�-��Ua"Vݿ�jX	���j���q��.`V=�-�?��!�*��p�Y�AN���g@R�i(X�~!#��s\[BG� 9��v�mGe���C�re(i#@U8g����7�륺T�x����b�n�ǰ�?t��鈑9B�`�Q5�ޡs�!u��Z'ͣUV�"\�	ҥ���i��2^�*TZ�Wo���C���-@+���ůR��T���'��v.�'�v|,��Cb�3 u��~�,�@��]}t{'?�y�sǧ���R�Mi?_3o<�q"���[��2�T
��@ %��%%��!��\+��;BL�n���Yz���䙕@(�O|��s��df�9Ẓ���!�q ���R��W�m��|��`3i�2E`����J ������b������P�V���gl�؆�<�/4q/��Ɨ ɕ��[��N&����5������ّ��x!��$�Bs���ޠT�,�V����q.�2��h�s~"�c�c��ѯ��ըe�ܩ �� �1��{�>{�먕��m��<'"�����nD�Ҕ4ڀP&�<�Sk��Hz+�ev��\�rkq1T�@f ���\`�c�R��èln(���cZ�Ԗ��WwJ���V�1���yԍ0�yP~��.���F�¥�(#���miL�/3u�<vzu���گ"�ARo�{�Ȯg�������>�Q����F��2O����%1%kʎ �W���|��z��cB"��\�G!��`�HR��CeEײ�@|�P�|���~2#M�6�~�I��G��������횸���Az3��y�7L�`�|�T��M���[N��C������qvU�g�WVL7 �Y������M,����EM8�-i���{��ܛ Ê㢲?���
�)�� �G��*�/��͹5�`@�k�[>�����0��qL�L�l�o�5��𕇫hu>R�ə�a<����Gj����<#D�dh�43n(健n7�&��+�*��i/o���!�m�jq�O�T���o��q`�oH�VD��AŒG.N�[W��(�
����z��%��M�'����ֳ*���b1�]r2��}������r��ξ����'gߚ���=F�7�"Z�sFy�㑩�u�X5��7!:���.|�&�i��E~u�/8S]��Ek��\�z�P������m+r��yػ�F<&��i�{L���Ԡ_�B��Μe2#�\���5��]����iH���LhQ˲o��?N8섢���8����xe2���k^~��2�@�B>��d�پY�+j�lߡ���E��,1%��^�g��GS���;���9����(�NW?[S�G!�v�@ߨП���/�@��>��U���+~�9F_](0W�������`���;��M��H�\���&j޴ցV 26 �w���u=|�g�w�a�����E��r�ĩ��ձ��<aRO��Ik:t�Yӹ��J�]�����x���F�q��j�<��\����\�9�>M�y(�f]�|hA4 ����4|��N~Gt�2e�B掎H:x�}��c�X7w9$��rB�g2HuGHT��C���`�A�Φ�0�ATx�������ܽ�0%�s���G��7-}�
ND2("�!�����)�dۙ�)N��6�=6ٙ%C����:��o��+��9���r�Y?�
���f'I�:x� ���i�zSޞoA���p[%�׆A�
)h��V��@g��6f2j*�d�O@~�Δ�P ����Tr�E��X:7��*�J�~�����f�Ο�5s�}ˑ�+;U���5�?7��
h���?D�õ@�әU��PU߉a�~c���|w�]�]�a�)cԬB`b�6���@me]�=�;}�*�0�+��`�C�q�d�|��N�^&��S�~�à��NIA �2�ܓ����+'<�2�N Yp��F$�٪�W��<i���Vг���7�ꥀ�L�!+�������<��ĶP�f�H��OR��|���?����*�������O`�Y�]�P�Re��LO<P�)5^�x>�w������	�;�0�$z��\b���H{���X��ö�� G��l�w�<�o������Q����[
�8���O~�!��lf��0�3��~5��`�zi�La�z�������5e��0��+���������I�F��S��tNb�ݏ�z��4�}�˿�HܯC��(��?s_��A|���f:#��e��𮉸BdDW�`6��8�9� ľY�CA���F<Gbz���X<UaГ�g�:@�� �oL�`��(���xU�r��
Mĭ�EpV�'�(W��������L��c�eէf��R���Y�.PT���|ʴ�d�T��&*��`|:�By�8�g����h�{ރ��z���f"��x
�ܝ���8���:%*6Q�\�,�Ͼ�,?���6 �6�Dl�Jd��kEHP/��ko�l����zn2�?f��#�=D��q4ς9����@leX�Vv���5��l���Ekvg���L�yÅ����l����Nq�Bt�"��_�r#^��Xo>2�p��a������tS�%u0G�A͸n0�
�.�F+J�Ƿ�O�]:UfPD�Gĕ,�Av|��]��z6���|��8��T��`R6h�a�vVi���n�0�2y���e���zm�ܰ�@,6��Y�<�q�����u�H@�演��w����2 q!��	���P��̼g�X��u듯�D·�[M]�[�@�#%_�
ֿpNj�8]��t�����'W��v���aT�J٤���/����
�7����CBm��$��Eb�>m�2\���J�ê�MY�}w#���.bzΕ���?�J��,��%?�b�O���.�箙���H_~�u�;��(���=�,��L8|��9l�w�־��*���4-�g�+�{���߲�%q���֓}��F�C�b�P�y ����rS�a[���$�"��A��K���A��"�G����IOB>���4 	:�G�7�k��%5ƅ��8t�ړ�Tw�t\��L��|��֣·]H〖y�^
�F�k��9�HZ�*�PW> *�_�k�=Ճ�>V}TtYwdv�2��FT���&8�H˟�bI%5I`�ٹT9�r�-R����A������1��Bx+�>K�a�,6���|F�v�k�V>I�p��/,>��B�s��08\2�
ئ¥�I�$� �"}���~h2i���Z�������<������)i��`A�D�}	!���_�]�ҍW:<xn�C�`�8ݫ��It.�?wOxX�ޗ�)�_�+89������ʵV�+��"?]�8Q`���<��J��A��/ƌ�
xiZ��N�yn�z�X�Qѓ0SޤD�S�bg;�(��[b���E�DS��1A'�Kqڸ�X�gq�D��J�X��sL5�gg%%�Rx	O����������߂>��rB�KHc�Z~Z��~�$�IP�~Y�Xlt���i�b��6��	���c����T!���ZS�v&
<ɡ����>�eٻk_T�h��b�N�݌�,.��uy�ԉ��m]s��C�B%&����)�m��֌���h�#<n��B�kxRہ����Gn�G3Yb�n3	�B�_�ׇ5�*����6�F��(l�#CjQ��1��X֜��谻���Uݬ�� ���Ǐs<*���^��Cx�jKFԞ�?�mq�k�K�`�Pg"���&�3	B�g&Z��^�ӣ���p����tr/�ޕk����H,�8yN3�F��Q,��K�>�|�a�|o1)�t�qӛx�������z����ʠ �܆g]�I��|q-fۖ��xG��?$�ҹ� u��ܳl�V�Jx�����"k��n�Q�A+ԭ�P'l8��a�e����NC�C��&�E��U˄;{��:����؜�=Ϥ�v�c+3�h��s���^<Z{ky��[��B['v�$IM��O$��a���Bi���qéQ����P)��X�2b�̫��յ�n�V�8��UQ%y����De�~1�S7`����M1mn|�pl�y`E����Ȱܷi~3m�X�F#��U�&�O1�孶�R+ftn���M`,6��^Xpj�0q�q������[[d�$>�>hp+� hG��&o�(����n̪�b��.	�2Շہ��ioHZ�=�a���2�J��k�Y0�S��U,w��bQ��2�<{I:���,���q;�@��yw��<�
F"d�t�KiB����0��y������\!��"질v�RXP�H�����V��gF0�m��e3m.Ϗ�_�	U�~5��*�xV�nw�s�67�P��T�t�N`�u;t��N�`V%�|��5�'��v}�7�:�4�p������{��p VJ�w�k����,&��q���{=#vZ�i�k4�������6#��E��f��ͻ y�n@V�:c�o�ު�V(��î[Q/�2$����ҏ�O'�RI�� h̅����{:Ib�H~�[�PJ�8фУ������w?q4��l�5,�YkDm��$���ʶ��1����:Fs�]�T$h�+��7�c����p>�5���ݨ�^�3�Di������ͶE��#nD�V
�2"��D>�����|{��ͬ�(��m�D��S��p�Tr�g��~l�Y&�, �����=���J{��Ba������2p���5���Њ�gw��{ !Љ�
��O "s2����2:��a������e��Y>��E�H��:�i�2�J%�� G�RZPz��x�V7J1�[�d�击�q:�X/T�S_X�]�ߟ��؇M�y�7%xl� �
��-�"���*c褾����9}��]E��Q�>����;�K[�FC���f�AO�]�x��j�9��>�Pr�LatH���Ugw�����\bБ~���?HO��<qx����`O�V4��'�s6*�#O`}޲�ş�=�Ww��hc�#ʘ��GŅ"��w�}_�&t('Tu�P^��Ǵ!4lt�D��5��[�;Z�{���F�uI��W���.!�X��q�(�pnCW��_��w)�̮},�z��JÉ�s<l�)ӑnw�<�� k���T�-5�����'�-)޶&M��#�u�o�D�|��0lS:@��1v�s��X1�$)d<Oⶣ�l�CLV�K�M�!b8�@��b���{�$U���]#Mo7Ҷ
�%0���t::��Ⱥ��2.�D^�B�P�œ��(�_ ,0	_k墽1Kܢ�X+x���iAns���8�(�&�q��dދ��P���Z$�����l�s.�ُ��_ʑ���4X=�@Y��Xh�o�V`�(a�,�j�k� ��Ӆ���|� 	�0�}`�M�����9��;Ue?@9P����M�~/3o<��2sf����j�����b2��u7ZYV�� 4�f�o�\��j;�+�׌�aJNl1�È&����[T����߱��2��yW��t2L�N��}8����$�@��u�����G�38���'J���~��G5R[�+��ͯ��R�vaE�=���/t�|p1(W�.� S� �*R�=�2����8�257"����}�/��?�W�n�R��n�t#�[^����
�S}���s��,����|�����|l	��q8�*���$��cm���#(NT��i���7*��m�k��],g ��	��W���-�'�@<�mF_��]�d�a�zm�1��=En�`!����:'#X3�~�Q99Y}/��
�V�r�_vu4mO�C�h]3�
N�4N�����~��'D�.H�9]>���RG�����ͷ�iR ��/�9!k�gڣ	��5B�����0���r���{ ��Z��z�6`�qW���y��b8�?��g��N��Qz�v[�K�Q�o&JL^! )��+�a��x�!ɄB�wB����q��� ������6�?p��c��}���FL�/��^N�A}6����o!T����Ѧ����]��'��RH�D���NdgZ��Y��(DX�ʡQ&�m��`ߤACp���JT�ؖ��#�s9�?Ֆ�
�8i<b@p<�53&�JT%���	�#KbR^�'ñ��T�Ƕa������1oW��Q�H�N��H�?3H����`c~�E�������M�d�W=��GN<p�q��J@���`ܯ֜<�2��)��y�#���Yr�Ph�F�>�o�X(	Uā~�pC�
s̱��;3&��v�"�f�a�@^N�����H�L���T�S�Z��xb�Η�ɑ,_?f�s��~!�,R	ԣ4��VR�H|d���c 	���5�obhDh��]��Sd����AD�*�׿�M�/��T)�*T�F-r�gw�ދ�K!f�\2ȧ)|iȭ�j�7����ip��6I�T�R"DK= ��}��F�[-cu�+�,R����`wٽ.���I~��L�i�/&�����flکE��0ֻ���:O=�������f��!�M5���(�c����%~UmL���剈� ��ҨoD�G���.�둰=����"&H��?���O���^���Ab�j�yY>�x��O塏�aoU�ڟ�j#Ų��!��pe�S`�L\��a �:�I�-���d�1�W��&��z�~>�?�7V����X�߱A\��ai��Xٲ�������_ٍʛ)�ݍ����X An�|#'�^��83�K�Um�Pk��� T9LD�B<�Ca6RӞ�CfS�Ɉk����� ��3!��=@��-�!�튳�U�]��m�.Gq�"��VO�s��p��I;a��KAk�f��~3<"P�z����b���!�t���}��k rXu*�=2�?:�$�_�#}|Ȕ|Ë��s��W?���~��'�{*�O(I���5��?��k�k��oC��xs���b]:�y6�;E�d�sE�̗��&�-=r�c�H�C�#_@���g�x5+E��M��^�݂�����~���>-e����9ͧ�,�B9x�ą�����`���z��&S!��N��B�p���&�i�Y\���%F����#Cyr_�̳��0���0�#���.�ә�T�DS�m��[O�9���?��$.�d����x���6k�1u�S����d�3TSv�w�cѩPϝ\�ˠ����N���{�(��p��y��~�z�?�m����{�jU�Бt�*�]�]�Є�Jk��FV��r��_�bJC���2��P_)v">H�������Z����^He『����=�'�L�8Q�Oz�+jK�C~>c�����G�2ވ5��_�d�ύ���?4:F��!���N:^�Ƙ��R�O��N>�<Ϧ`�g�qn� �"�K�3�}�F�qQ���z2��fy��ϝ�'�)j5�e3���%�#m%��Rs�	P�w#[n�v�ʎyѷ���9nJ�. @�]�+@�����ǖ;lq\�V;���{:�d���Ԍ,�I6#��΋�)���pWU䛓�w��#�����퉬����>�qj����k?IPp���M�|7���"{����R��]�
˝=�	��p�	,)�pqY���I�Y�����-�-�j�?��>�Ͷ�+����� ܤ�#�u���L ��`?��x<O��)��[�%��OJ���#t�(+_D�%k~	��u�a�3��ɔ��]���0�f3l?"�K⁝R�7!6Y{+���%�Ԗm�s���hz���
��e{KW�q�'!}�I����DAr+��m����H�ǨQ�t����:�U�5p�p��bv>X�	I���s"�:
^��~���yfW�N&9#H��r(Og���m����?�̵0J��f}�	�򍞃U�-�g{$��b��2
�e����!'��^�ҕ�H��IT��+�e%��?�p�*�ڨLSIʞ���J��"����Dz�]|�^Q�q��Ff	�H�#�x�/ya-���w��i���)�SI�`��N��mB
��A�w��#9��e��Z����=�y�:bǇ����?��I�^12pQ��{����Z�M��	�Q�������$ð�O���n�4���K��1M��V���XR$�f��gi�܏�j�{��a`Z��ٮ��b��Z��I�Lg	=CV(��s�"g��J�<gd29��(��"��:�͗�I�}�����8\h�����������P+��GTp�������s��m�����&<���Yvc���ّ�~[N�xr~�5��t���#�����9 ��zpk
��d�'�� �����2���0��>�C��Ϙ\� i���޾�fuƶ��������#[u� 6l,�?�^�p�~X
�;V��w���f +����>GMg`o%ʊ�K�:�1t������2���Z_W�Nʒ�{O�bÿ�ܥ��Ch ��2O��ymBj��q���gQw��|K�a[W�I��R���%ݺ�-g�`����d������h<e�"��������R�'�tUU��fϲ�W�s�?�+ā���o��V�(9�l&7T<eݼ������قԧ Fl�� �}���ܺP��#`��F8u�$|2�ĪU�������4i����Ƚ��
0/!�� �& �(�v�r�@�5��ҽ]p����O�#1�14�<��5�%1��A7�_D�-�Ɔ��
��f�,ff��r�B�۵]�?��5ʟs"��|���m+�޶?e�˖QũX1b�e#��,6C���F	�m��eHt|Q�����'hN��c&+�1�w�|�����R`�Q���̇�.f1�Π��O}ʷ�6���0�z�yi`�����Q��\ۻ��}�D5�\}��`"������ps��uR�ѹe��Fת���7��&�S�)���� �j��9��P�}���mC~���0S�p׏�P
¶�nN\ W���ڵ[b�ɉiU@���W�9��zQ�Gg3}DFp4bZ��3�T�����@%BP�����c�����;ŤU��v'H��ٺ��0I�=�"�O��7�P��ܳ�'���������Ơ�	G)����/ $�r��Sү�pQ���V�������>�ntD2[m8^0%2���=�\xrR�h�|�� �[;��X�A�ڥc�Ȅ�r��uw���
�ja��E��wg>1��Gfޛ����&_��N� �b9hE��(bl 8w��9��l�FŢ)�z��[y�iW,@�[�J�P���o)�J��_}y� ��^K�3��8pw�e�l��
?�q5�'4&/5����y����TEP �Q�� �ν]K��s;���T%�ssIbW� ���>,��/$��y�jw���,��*�-���G�%M�����k��ѥ6[����.r#t/�T,+�y�O�;Q���'�(�[:�"-I��稜���u�t*g��S6�1�3I;��T�k
�C��w�<:3�D-Ǡ�m��0j���\��;ne��n��z�2���$g�(_�)_"�q$�hl`&R<�6&���(/<i�KX�sG�V��D�]z��Iҋ�R��["�c�N�D�I1�� Ǟ��!y��A�[���y���c��w��ʏ��|�%�1؞�2<$c3�����J�<�oH.x�8�G���������-� '�0���~��V�Ǥz��OU����.�� �TʢGBZb'�0�Ӳ�xchR�ŨGr���_ ���;^ܹ�CR���˙n!:�sۖ�T���<�L0��bv#�(9I�� �۳Xyg�dT�3S�k��v���2�7gщ�`��*�����zY`�pV\���̇�+K>��+�'�_�юF�4�3í@��tqa�ó�E��(�t4
Ns-z��k�OfG�ֿ����Ӡ�RGAkH��A��N��[P�_�S�P�ď��q7��Û�'�u�-:�J0���+*B��s����|m����8�eγ[2���Q���K_�\5��I|�!��M�b\��M����|I׆�u$Lp�Pʅ;5����!Q�Iū�}���f� ��?ݴ�h�x�����=�NF�{'�IQ���T_��"�X�=:�'�#�&�5O�e( %�����q�猘�b}�,�J�������̓F�^Q:�y4�zgZ��:�hB�1�G�}F�,�@mh`���yW� K�BZ��J����#q� 5�O�|�apw��ړ���/\�n2���`H�!f���tة�3��lt��hk'��@6Me�>���/��NO�6��ғ��|��ϫ2]b��(����Ƚ�n��= ��re�1��݋���}��U��!{3]��k00�hǊ^!,��'%�(��;h>&�f��饩 �H9L�ʌ�ԉ�`1M�;��MQq`P4܏�qO����?�\���W>hO`$?[��Y<Y�i���;��A&�� fn`��n�Ҍ��k�b�Yx{�E�0g,�6�poPK�\�݌)�63|AM����'�F�q�p� ��Yf_�]�0��c_��M����
�p�2�P��jUxtb�c@��NIV�g�1 �3@	u�����j�4E q��ʺ�*T�H�����眙ĉ�)Q0Y�Wi���0*��{ǵ��{�?���n�	�][�g���7���ʻ��خP[�v�.DR@�c&Z�^�mD�͗�A�Pԍ;5���mb�)��e=yCs�YV�(�cq�G�5yIh��Y0����J�Wv1��X��]M�-�,�(�4`����L�kQ�9��X��D\��s���7+s���Z�V����,�v��{aE۳A;Q5W�.���2�M�92x�g��*I}��1�@����L��
6Ў1"	��g�V�D�# P/+BX�C�^��������@M�����'������<WS�V!Q%�8Q��m���0�W��_(�1�:����8� �ϖʩ~�s����$V��E�*��K�$�>�Z������`��xD��B������*���I�Z���r=�0����m�e�� ���-"^�_3G��g-�R�y����X�Ck7󪹂(gA=g�c���h���C&�g"k%���vp���N�:���P<��(��i%�N�U�m����\Jt0�T���YK�:f�� i�nu�NE+�k�r�m�;�=��f��E����M)������i״e���Hw"���14`��Z�@��s��S_B)���*��n/�J�V>BU����`u��H�3�7&��4խ�#pG �e�J&_��>#jQTtB@GOy�rQ�!\ټ�8?W�Cq(�\;��+��8�t*,1�(ELf�����{ydUL*xb8��OƇ���ϘWْ~�u�Ud�ѹ�x��ĒSȎV�
'�l9Tz�i�»����*�e��Y�xx��`u�g>�`�4�I����:[�k���(�VD��h=����{倹3o�g��0;�!�4�Nk�>bա�bw�����x��Ui�e╩�ڗU^3!�fr_䊆��ȝ~Rd�q,�6fp�'*X�`i����w�)w~F8����z���\��vf�u�a��%���f��KA�J�$ά�!$�Z%��9�/��9��6
y���;ECAW�V̸^�~{�"J��,�>	 B�ٶO���U�h�M#@t��G+x��!���]�^粃�=�Az��̀���l������������u���Y�9���\b8״��[����6�n0�#���;|���uܟw�>�(ᐲ����l�8�!6+�I$�sa��_�UQ�����_ �g�;Z�,a!�/M�}F��ۓ��������;�/�+'7x�gׄ��8��o�?�?V_�S���i�W�byG�5��w٦�huJ���ΰ��)�,}8���10���lf�5��W�P[����Ώ-w�E���^@}!i�m�N��%�d��` �����޻Øok�����k4�[�eH���)~:�q�$$�9,�N����k�o|�G��K�\�4-;R�1�X�*!�LV���}���??7d}��]b��V)ԿT��EiL��~v|L���sP�Z��v|�٥�w;qNJ�v��T�oR|@<�U�4��`9̯]E3�����M��y�hj��͍w����!��J�}��������옗jV��H*p�^b,�i�I�zI�*�-��L��� Z^�!��ǞP��#�{�VT O{�r-/��i�>������BΣ&��X7z�h+���!#cbс$}P\�P�#��aca��"�OP���5�`�6�M�`������O@�z�tEB��:S|���4������(��gg���u��1p�~#2�����~��oo�N������Ò)_��4��Q�'�b�^�@�q�A����w�WF�B{����h�x>�ʫ�31FR����O||�W��g��z�Q_���V�H푶�������f�<�ƛ"[}�u;[l�m,vD�w%Y�}�S��'s��z����Y��S�@M�PkA��-�+�\Fnw,��5�8&�z�O�x���汒�$�������M��G牚6 ��^m�q� �,"+矹`�k��ћ�&���5���O��E�S^# x��,��%:�lDi!��^K���4����7�1��h��Vc���Ry<�LC@Q��V�,9��o�ܝ�C�,��IJ�B16���!�:�P�>��M�l�h8��{����������G����Yi���<~����!4í��RE������ou%��ۣ��
��V��yQ�'+�􅷓���8�A�褣���[�y�� N@��f<�<�+������v�Eu:+e鑿�r𩉝�_�WR�ݫ��,ו��1�:'r2/5�3Lͯ�<����6�b����=\c�!�"����\kl�R ��UkT|��S� ��yt��(�&М�:�-Mׂ���V�`z���ψXV�T�����8\26������5���K���z�V|�#,<�wL�E������]T�S�!>����]����Y�/©<e���׭u�+��9��}��z��kJ
�rڝ+0߲�%�����Xj�<�.ࠡYcIX��j��=<�
�� )F]��2�kӤF8c�bV���ʋ������K[kڏx� . ���/��}"�Ƣ� ��I�7��{?* -�k�1w�ݷ�:�#�qU��;|�"�MR|�E?�b��������k�I�!s/~f2=��Y���n�?=��kW����fdP-��1�g��B���:��Y�У��P�I�|1@l?��:�j�!1�=(���[�C����pP���*�ذ�?�sII�G��T�&��'N��v.q9d�&g00��t&x�}�%.���(�<��Hk�mL5]k����i�΋��m�ҟ��n��Voo�z':t� Ѣ�S����G (��G�]��5�R�/3 ����[��H$ٲgRh�{2a��J��Kj"-��a�e���W%[��E���S��xf����[��i� Q�5��C���#:�9�]:����^"#*_��P��F��7:��<�\kK��=�0m�� ��L�=���9BG1�ldkճ�
��ts�������K�fZ,�(��廊C�D�,=�i�7#Ah^�Il�9˦$V��,&��OS��� ��~�1,�ma&�'�Yy[�]���H�G8�N��ǲ�b��lYv5Eΰj�sO��sM�a�����A���:�Z�1<K���9ۺ���_$��\�}�6��U{ˮ���'V0ܷun�K �Г>�(؀�Vo�L�v Լ��	x�=9|�p3F�)�	A�����j��Jj{�Gn|�8S|�`�4R��f��s�*�9+0�/b�G±~��a�s���a�s;������6���qЦ)�����&��Y��aU����Xt���ϥr��LN[�[�y-I��� @g�F'��&Պ�Ɵq��Zܓ��0hd�SDZY���w�a����A�'�{�˗��#yY��]뱿[��V$@8
���vI]�eF�Ի�F���b��ɯ���;��g�j��b?Zm����J�i^��Y%ً�����)q�4���Q����nuۤ��Ѭ�5�$r^�(T�6ēS�/�8=~3�ܖ.���r4��L¼/MR�P��>�����)򚙦d��Z]��醦)����� ��ڕ���7���ĔbM �
��>��#��$/��@FU����3f�!|�?Q�s/��`�'GJf@�d���������ƥmz����tc4��}	̧�����B&�O����IŔ���������f�6�D�7u���c��1�CU	�����>����b�	I���O�sb��������,�=c���φ>����	!�<����
נꅘ�����)!�	l_7~[6�Lc/��t_�~�
���ΛO�]�.����W�Q^U} �Ģ��َ������|��G����B�0������܋m,X� ���������C����:f���w"�)����;����k�kA �dw���fn���t��6H�96;��9�3r���t���1����j�;i��X��;���(z��1�&�)�..cc�PMi^� ��B=�������|�HBqs��7��4�p��ʰb�V��GS��Q�ôa��\��P��m��B�i}h8� ���ȑ>���,.�oA��%�~��_�su%/��([<4c�T?��(�c$he2rn��ݰ�I�I]��[|Y�/������x�'���/z@��:b	�[
L�m9��{_*��������]:�E�uH�s�o��la]�fbb�&.�����c6A.{����U���b�,�&=q
���߹�ʈ�Ӗ�%�2�XT)�:ܘ��)�ne��a�K`�.`�<�E�K4Ͷ�xgº�2�;�5��D��%65&��#X�!��t���o�R�p?���+ި�����<Y�w���y[C����(��Ǒ[�pG1"�/҃`�|Uk�N���";�j�*� xĽ��t��T�nf�s&[�����E�Kˣ�b�c���,p�����w�I���۩3_9&�ju���a��-]���i��"�B��sM?8��,��h6�~���� o���.��Ddd���l���0|WQ��u�R��~e���DK�veI��M�l�ట*�aCe"N�f�4��ɠڪj����CG���o�����������|ٮMz��B�~d�ő���0,n.��|��`��HC�'��H��V�
	��T��9o>rT��������8���2HĮ\X���w�q�	g��JjK* B?OJ�׃�x�;���ʴ����A�̵�Yq�f7�\�x��0�����Oi�C���F�u�r�l���"a��B�d��5
D	��.�g;=U���ܯ�� ���=�DL��xf9a�sh�'گ�[[�ki/��_��N}���Uɑ�!>�^|U�I) ����ɪ��$P�޷ f�I�0 iZ�W������/Sr�KCW��EX3vA�'-��?���	b�n)'�|>|�Y,��{��9x����GU8��0�����ϋ!�6��;��'7�o�.��F�r�[gͭ�V�	!\�{(�2�?M���:��GG��a0[͜0�������$�`��})&Rdr��^@N�+A�	�ɑ�"�+����P�<�"�Tpn'-G	Ӻ~O�ʫZ��Y�?4�?Ե~�)S"*AK���n����[D@������k���7 f;�6����&���S�F�PD-p.�2SY�F!��o{c�t��o�eý�q�yE2���n�+h��0�Bf��"�{��EL&��y%���t�����1/f���n U2��v�)m��[L�A����>��n�����ԘP޶���O Խ��(r�ͦ]�p�H.��`]P�@_F��TӚY�|�y4��.X/p�ߵ�c�W�h���B�bx=�� �]����ϱ�A���4Ϳ2�r�wAz�Z������6Ɓ7	ؼ�
ԚYj�䲵���z0n]8�L���A��P4�2��,񸘘�p�hˑ)���
�ɀ�]v>ԁ?lp�+GA�.��a�m+�I,Z͠g�
�L[bZ�Q.�)���l��)H����5��p*k�SY�ND8�G�̕�<9&�`�wL���u=sKFTJ��O&��|d}f�!.i�A��NZ��V������=����������NPo�os�IK�vXք��ut+>�0�N�q���e�l�v�o����!�ʡ�u '
���tD��$��F}���31�ge��0�Y��G������+���C��_���\�v4�����+�8�á�h='�^���� �Aj������1������d��çq��Z��
�u��TU��4;pA�v���F�Z
[F��S'���q�a0[c��I<8h����Ǜs�V҆�TEF�
H���{Yt��UÄ��:h��u+��5h���!��J�D�8et�h_2Y�l�c ��>�K�Q�؟o��d
,� 5ׇ\�ϸ�j��N�����@BV� qg��ְ6�6R��[�o�U؆\�W�] Q�o8F�Ds|���7&Q�'����͛�W�#�]�b
���L��㵫b� G�__R��kN�֛sajd����	Gj����@I7�#�P���R������#UX�zg���T&		o���&	+������o���>�0̅(RL�0�g�1���>[��r��tƐ}n�J9�R�d)�p��"�����o�+��������*��l9���y�>����E��%�k'���6^�B8
Z�D'�P�o�93ʒϧ� ��:�!#�)����+H׭��`�J�TT�`����<@�;`���vJ�}`J��iB���!4g�\F������6�R������HR`��Z-t%:�g~��Ň?�H�I�f�MW��iQ����7s�-�
Ņ�Z��J��)6��2��߶A$������ݖ��b��GĆ4��<�������z_�����2�-�.��[�t�}	oO%
���D=��bA������*�|�UK�����o����W���)���/�G�Y�}MT��j�4��`G�Zn�a�N'8T#dc��U�)T*y^)Ze�$��,5ju?C��	��1�/��Ǳ�sנ2B:���vx&⯖���/rc�KA�?�xeCj���w���$��9鑆�Le�}�d��d��P���[�@\bhZ��)��Y��g���� �qt��P��u�C�,���V��@����Bd��5D'곲`����?\��ڑ�,q��rR�.�����&|y|�pHW՘�sT����5�$�E}�=���;B�I���G����*�
�_�2�s9�ƸlDncR\�D4� �+?/2A�������*B��� ���ۥv�N H2W�tFh�ٗu[���12)O�~���_~��,���Y��C�{� �x��h�#��rb�'�c��uy̓D�i�n3����<,�u*�f��L����XSn�$��=Ǻ��gZ�t�,X��6`��Z�Am��hO��=bs�^-����7NA���g���tw:F4Ԓ ~�B�����y���7�>Ї��mX�9�>`z�f}ē��]%%9SO�@��
���Q~�H����eʨ|�h���\2�s����פ�@z4��Z%3��7<k������=G戽��:�N�(��!GK����F8V3ye�>5+�kN�	�[��f�e#�t�6eք=د,#'w0�tM�X;���M�Ot4E.$tx'S�.4:��͗އk����� ����Jz��5�E���V1$)5C��Q{���7�`"����G����^�6�ry�p���C;;@u���om/�	U������l�`�{��C��2��Vd|���!�Ѧ���ο�,%e�#��ߘ����;M8������{���׭�>��y�D�=sg�:�"�ڰ����	75^>�0���Q�}ϒ���
*��N0ؿ��,�{*�6ᑾ9��0�
�T�oX��7���Q/0fŤ1��	JфKRZ�-��wh�9W�{ݘF��M)siB	V�7|r�!�cЪy�m�-t?����h��a�"3Y����D�����0�F���#p*�e�E ���/k4����L�C�?N'��G���3!Xr�����)6����G�-S��"�ڤ�
���H|�3�RGW�+VD?;mΣq�&V�t�{�XYz�P)�\Ԩ���nZ�D�e���R��TuE1��ڃ�X�=�fw���rd� C���2���2��fb{x�8��*'͌��
�ޔ�x��� h��;����f�+3�n)�c���`����_Ӆ��B���؀k���1B!m��+�n4�c6��~ƻL0R��e�w����XsNŏ�ʏm��ϱb\��4�OҠ�Dl,���cq�s6����`p]ɭ��w��x2�m�Z	��d{�E����xY�mb6{׈��4h�{�����Z�R�V.th[{�d{���)�;+����xsT��{4��5��R�Ѕ��C��)��т�"�\[l����x��i��� d
��s �z��%:>�"2�A@_=�O
����q�����"8������5���>h#�a2��ɏ)]Nh��eэ3Q�� 审�ߖ]�p��8ž���:��N)˓p!_|�f�9�����U�u�#άE�+D���I��i�y�d�}CF�7���BO6iV�Ōp��M��c��9M������7:�'QH#Բ\��!Z�ѽ�,���Ͽ��r���BS̟��Ì��WW��6F�v;J�r�B)�*�9v���&�0����µ�U�5�%T
yb����ke|���5`H.~9u&�t��q���kI�'����@��ժ%�� B�B�Ԣ�PR|C�Rp��*rn��H�8��Ɠ��M��m�0.=���,7��,�M=�?���'%+{I�֪ȱ�gl;~+�� �<�Q��_�ɸe�Ng��Ʀ�4P�N�M���_�e�+; t�yu��w�"E;����H_����ŔfJ+ǟ����,���^;"\�R�	f!��jG:��w,�v��nHĤ_�؂�e�{^"-��^7-�پ�;3y��H�饗u�a�O�+uGߩ�dk�p$�t�T�u�h!0���W�FP�Ϫ�k��#.����ɞ@�]c�
�����J&��<�G��j�g���e�:a����@ ���^wzo$���6��B���he�_!�VS�)���-�ӻ>����#��4��l�T5�if+�~$)�����qq�Z
ܐ}����Ǧ�����8B�S|آ%�*5��C7Oأ,҄ö�HC������O����f5+�j�!���ĵ�l_`a]<l�����
����k�.9L��2���F��%ӷ�Y��xS^W7Y�h�rl4��#rD:�e�;9�3D;#�Ͱ���{TA��j7(��2�K�	8SѢ���ȎK �J����!�;��������p�T3�z�n����s��I��R{E����?*�GJC�_v�YdԔ�:���y����@G��D��8o����]K���cr����ߣ��H��[b���U�9t߈�����8��獻���G��U���y�\ �Ԉ1�Z/���['�&���Ju�mR���5P,�"�r¦��Bɚ����|�v�^S㺁�����n�V�'RV���� �a�s���.k6;ͪ�#p:\f\B�RM[�Mc8�I��\:��*�y�Ć�8�E�� ��[���A��g�n)K�e��r����G������!a0o��R�ֿ��ܠ��̅���3|�ӛ��hR^�&��?�F9����U?.��"���=g����"(�� ��j!\��+��JyI�kZ�>	�11{�L�D*X䣠��f�#W(h���C4/�PX�����θ�_k}5���9D�Umqx������A���sZ�XIi5\�ܷ��hr�5�r΀a���ԓ���R���7�Z&���@��-#-��>���~um�`hx�c�@vn^�ԪD���ކW��ɏm��9��^þ
�O��+
��l��Q��Ԕ6����6(j�wF�po�j�z@��U�,3m��C� _�F���Yq�S�'|c
��ϟ`@{:i�hS1��p��V��
�eR���l+�"����fwJ����*5�nq������*���" ��� �A�k���B���/wj!m�v�Jd��0*�p�!K���>.��1�ʼ��],V�a��
fU�NJ 
���&l����"l�����{*�AW5��
���Uo!ϬP[����|\+GE���QB�h�ٌ���� KJ��6l�o�쵿R������=Ko�D��ߑ��Y+S>9���י�Ԑ��󷊍���uz��ISXoAɎ�b��]/_�P������[0���b�Oe���<0��6)H��1�[Z���e- /`v:l�!z����m	�u2�̝��L�slHܚ>5k�Z��g�2#=چ���0!��1*b5?�&�/H@p=,��7��k��@�cs����ǜ�tϫ[�ӿdA��A2(h��G�h;R��Q�l࿽fF��7�AWώ� a�LK�I{zɰ(��sݹ�)��[�aw��a���-�����aF���R�;�8"���^�j���N<^���NV��N�Jno���Mu�,�+�g�kX�?�f�q7=�Y��Q#u岀�g��K';�\Xx��<}J�0�Kɀ�#��jk{����.���	��^/]��X���c䠾+b����)�Z��$�ܥ��2W���g3L�徛�(ѷ�P1a�mۆ/��G%��w�C�l�&2u�ǲGz�����K`�T.��
_�R�u���e1���r� a=q�,<�զa���;v��^uS���?�X���O��G�Z&&��V�Y&��J�ǫ$@@������:E���G�ق���-<��픣��#jH�(+��Г���:����+p�������Mg��=BAs4��9̾��Iʯp ��,�E�7=�v���*��������ʟ&�7�	��\���fV^)a�������|t��"��H��6É��Ɲ�+Z9��M1��ze��	*�kj#oY
��rL���^}'�w�������-����~��ꁔ�;����2�-'�R�r:�����V�>�#w���ԥ=��~zޛ�d;�M)ZGB��!*�}{�n�F^���P쪈���/De*���	_�s����wVJ�� ���֜�*��>��R�
�#�_D8�	�@��i��2��]��AtU5�g����h�_Wo���L��l��U�y��N�dADK�X�i��#5���;&h��RB�Qsd���O�L��~Fu�@�ꄶ��1w8��P��Ϫ��qp"]c�wh/Qn�&�Nm����-�N��<�@�����U�i�c=����C�J1�P);�q͑:�F{�f��U��R�9�i��~1Ʀ��Jg%�
��C���M7��hTJ��,��h�&�&�M�߿�l���jF�{�#�hy<��bޮ������/�͢r��V�'�:���D�h�=��&m/��,a<�ۘb<Ν�;�7��φ�	��M5�뙞���d�w��B�z\��6<���kވ�\����1f�-���5!��N�"��\�_b�'+�%��hk��d��>�v��J��K�'��®d2t�LK�mw���O$H�K�����,��R�=�SHs�`�%���T�wӻ"M?�-@�7iuK:d9;��2POh��(˻4e�,�R�{�~������el哏���-���W¿��.�u�W��R�2b �r⪖���n�N���79<�R�xd��ks�,���e!C���B���F��3i��Ĵ�Pw��s��n�Ϟ[�,eބ�SVX>�
�X"�C���W���&\��E�u[��	�=x��O�,P�ُ~ⷩ���\�~	�@Nz�DǵLs��Yj04ɫp6����ω+�R۴i��1�Z�i�ߊ;M;��U`�ǅ�XVي�3����TW���d�%X�J| � Wk�y��W�=�Y��z��ywp��c�����||��>_cذ��V�T������6ҵ���0�ɑF_�[�Jj�1l����+.~�eٹX�e�k7;�l�����6@o�wǼ�j)�Q��y�c�<�e���:I�Oԧ������%���{���0��	��ˋ������+��3�ꮷ�����+��h���(q�](�j�6�ٞ=��p�8\�䅰������H_#��^V���M	����RӸ�%ʘ���=�{����F���2DE�՗O^/��1OV�&�}������}�����'[k�Ժ=F;x�Մ]2�CqZ�B"rS� @��b�+�V����YA��#��3Y/�x�/��iKz?T&:��Њjw��o�q�S���R��U.e,���j=`/�\P�����mE����' ����'�";K��g����A}�c3'��a#t��W��H_S���ބl��� O)��2��*����a��bm�w���T�<?��b��sq�yg@JU9���Ο�'���\ڑ
�-z�iiA-�]Yv�2胟�FH[&(�h��3�A&K*�8io~�H�G�H�F�����8�z�p��U�S�"��>y�|C ��-�YP}2����.2҅� e���}��]͹	}?i���g���f^0f�w��#	�9��y���F&��	��\���dG�]{�棎H�>03^�H����ʽm�Tw���`�o�o��&�CK���!e��k��\+AM��oUЫ��f*�hY?fP��F�"6c�>��`��BمX����(��vl+���STAY���"���0[�HQ��Mąm'�̮E@���4ZU�M�%���wJ\��Zf,>�+�m��U5@i�_�i���x��\D9������������MӄI�~��r��Q  �Xo;J�6�W�#�ŗSo� �*�R��{�Ř�'t������u�Ze`�����G��ٌ��%�3�*���JlC���mZ7,Y?��=E߈��/m��T�Z`P��Y�X}�6�"0�O��-����d��|�/^*�;iM��t.���诩����R���[�)�w;�����I���9��)K(VU�!-1/��E��"O��/Bh��[c,ca6��K"��2��������;M�g��dJ�cw(�Hzbo��G��[
mU��D�u������\�`B�x%�ʜ�B����"�Ӽ�s��G`���Wy����#6x1 �N�;�2#_1�yܻZ��qr�֐�<B��Z~,�B���"���4�U�V���2��j�H���e?�Ё�7��b��s��锶�ע��uJ��33z�tZ�9l��P�I�&dC3O�%E|�@�F�Q��?�E�kc���0�T�5���ؽ}z�!f��"��)��W��X���Č�v�5sJ��<Ԩ��צ��V���ؐp�	a��M�āK,�p{���mw�8����̎g��=R��5�rwi�уdi��P�ç��I`���C�T�r#'�SFp�kk��g6��Ȁ�	05��!p]H����yR������s�?d��O�7ŬB�b�Q{�(O�0���)�Vd�[�:5�Gܪ�h�[j��d�
ܧ��v�i�c�������H(Q:�O.����{���RHI�{[�p�ɚ�h����0Xh������SĶd�1%�T�wqɴ�0�y��L��\3;O���Ś�����A�R��+�k���qعk��6R/��/����������l
���B�(�GԆ� �P��R����f~[6�����vڃl����	y���2���>\
�"�UKH��˓�z������z$��A@
u�1U���)�*l���&����=j3ă�Kl�49R~s����~+��9�Į��X��>!��|@��]�f�V��a���Y�ƶ"���[��M�F_D�?A�o��mJ��w��^�*w0�C��-}��!�2hJq*1��;�辷����k�"������h��=q`��$42�Y�F|�'G��y����l�4�QɱG�~�$�������f����d_��q��l�����:?�(B�Vp�yy~�]O��C��$�.�3�Q��$؟�])(\}�9��g��E��@�i�F��#�G@���F-KW��k)�0��n�6�&�=��� H�H��Q���н��Qi|׈_Q�*/�R5�6�:Z�.8]�����C���lwW��G�?<1Z?��	��jC�(S5���J(�l�f78N<���6f�'�j�i�#���υ����{Y��4��>B7'	��\Sj���� !5AN=
��'�G]Ix�����G�ȭ�V
��- =�'�{S�7�߾����MT�ْ4�kbZD�m��r�)�\G|��x�?�ȇg"_�����g�"016z�H�1C��2���R�Y�u����o�\�/��S�`y��X�Mnך"u����bw����2�@)R��X+��t���E�U,т/Y��O0Ck�xAE�g�4��`X�U����8S�#�J�:T"� �a�.�Rr})�N@��\�>�A����_`�c��K3�f1W�o:	nP5C����/0�{lu4��kp���#NAe��w��M��1����3r#���$i:f�d!	��i�@�9����6�ؑ7������'Iy"䶏�p;��o�:���߫p�X0�ŀ�mBby�ݶsm`E_�OB�OS�� ����'ǣ�γH.��9X�l���г��W+EDx)v�o��b~�f��3������K�ɓ�u
�I�����v�-α�̠4����isP���_*:l�zqԠ��뤏�,.����h��ߤ7�'��7)������h�
��X<��~U���zz(m�n�7���?���������<	�Oda]>�|s��#5�� DU@TtT�$ꗦ��I���eܲO�f����n �/����ϦB���f�����؂�.N�Zu����e��"}e(����u��k��Ҕv���iC�P��+;���O���T�#�tX�d�H��.�g���1-9�W�d�{
4uM�WRr���H��ñ��ux~�[t0:��M&;\���wr�rqn˴���	�<=Kٛ�q��)��]|*;eq��<b��U���P�����Uy�"�wE8,`�4�_ydm���R�U�/��.�B���^@�e�Xp�J�>��.){@~w�eD����!�H#�$�<+�F�t�&��{�y���u�.��0k�����7�X.W&�Z�����r�*�`Vg�c-�H� �}��	������d��`1+z<��P�Ϥ�������#\WX��_��H�� �Ϝ��7Pp[�#��Q��I�������"�
W*�^R����v@
��E�ǖ�)=֌���n ������8q�&m��C�%���Z��ڒ?������nB���7-�1l�'��G����='�Y+��Y�4]|A�O������;�4R�v��3��98��|S�9�%Y���FKb{��\��ׄ)w[�xhb�Ά�v������>��:�+���Bi�$�����L��bcr"�Ƌj��=_�.��W疨�$ҐNkՠ�X���9B$���F��#�H��\x��� ]c��V����K�x�v�亊����xƗ���R�p�z��Y�
+������֒��S������{�P�\��菠	�����75y��bI�i��n�����=G&MA��`]�&H5�g�硴��g��`�p?�o[��C�&4��L��\���@M_7�i�W!�D%6�5	;�+FP��L����ApK�~����?�݊������Fe��)����g .+���v��ߪ&wo�j�_���W+�sVn�GWSj,[��ܭ=C�`�X���k�m
�䂿�y�A^��A���#c��_Ɋ�wmi���>�@�Dz܆���pF=U�b�v�^�����ˢ˟d�k�����	�^�&��6G���ag1�o�=�f<�_¾�,.0�{�5iA��1�����,�ͨ�W�Ÿ5�f6RU��8i�>�.<�"�$^9�;��ִ&}�6�gA��(�߮KKo��θ�gB�0��f�(�j٤�pM<G�3�v҅�F츌��D��:��Sr��gܲ,\:&+q�Wj)��'��J�o�.y^g ��q��g�g��8 �8�^��_D����s��sE��HFҴ��<�����4�4��\l����ٕRG��s;�g��E팈���8򖖴����C�0c@�Ը`�s�-����K�	��G�'���gL����K`,ٙ��Rҵ���OE����������^����8�^��jG�iK�C>����h\�	�YE�{���2���qi���@���;e4�6�)�RlBpM�_YsބZ��Ջ�O�(�X(M�^��Ƿe-�����	���R�Q��'˃����JƲ����(�q>�6�l�\R7�c<��J㾰/�Qa���"��ǂa�xX.դ&)�;\�\�2���FA���R?�N�]���������=��t�xmu2.�[���N��Y=`�P�7�%��C�մ�f�:��S��/�Lc�K8�E�IN'�o��f� X�P��!!�C��ۯ�2��(��fp��1�H}�F�ӟ �w+JO]��wUF��U�
1�M<��G"r�#�\T�?i�FH��hNlp��ok����bA�#�Ξ���i(}/����2?|�~ ���b��Y�= -稖��򲂏�%)*��i�r&,7����T�ݎ�LN�8�8�ӈ8�k�e�B`�
�b�fl n����p��6��kk��B�wjb��X��6���h	�����!�`���p�n��ڰ�,v�YZ�r�-O�f�j�</�kKWm�8��!oJ�ud*hn����$K���W�ؙ,@�a-䚮��Z����j���r�#�ۦ���A���n���|���Z
|�9*:�#��M䀹3��|�/Jz��Gm��W����M��0A�U�CY�͜�m�\ ���x~�~p�O��H���rI�Z�����*6O��XQ�H���۳}v�O���q��΢#L��:�_Qg��%���wS��Ⱥ��m+��{�y<}�^�X-Ͱ[�P���1`sZ>��Ppg!j�K�M����6�",�#�
���2x�(֨����,���w����[8�����#f�S>�m���Gy]����{��7���r}��Qz]�K�8�Nm�x]q�-��K|��X���dr'�d�k8W��⢸YKrb����SX[T��a�+���x;8n_�"���C)�~�
x�)I���23�]���䷵o'X�x2���5�*`�C�yp�A��z��o�r�t;@��F��n1���M���1�&~�t>���XE���%"�#�f+tj��'t����^5�\1���7�L�iM���t!$����[�WQ�_?��ڦʣhK#�OJ��<%_[}ҙ������zP��fHl(��ZcR�j��@v��j�5�B�e�^��ɽ����9�������V멆��M#e��O3&\�x�-�x):��	z���W���x%r5G���)�~\�� �-=�K�� ������0FK���x��&�i�h_�E,�g����)�0��3��Qd���Y�3���?�-���{��#r-�[��V�ɽqPx�$	 ��`i�3�JF������`�¥r���=��N�"���!��j��u��~�6�_?c�g>�C���6�Z��tW�N�O��|Ah2�Y�7A�BEa a�ޔ��x�$��*f���S�Ł2�k�#��}y��sS��t����ܐ�j	��$M��a	�q��ֳ���c��I���y�x���.U�t(�l31�	���v���)�6:���B��*�U��g�;f ^(V�I����B?.<����4尉Y����R�oS�ΊzD"j�悸z}�=s��u�%�:��?��x�1E�>�M.Sn��׫Gq�`�T81	�LS/���+c���&�I�ĭQ�WʊA�?���'���X3hK�O��Q������)`[�D�]��~�71;HoZb.�������V��<}��?�nTm5.ROƵŻ:>�vCP�m�q��6&�8���\��]�B�19	)V��0t�p#㧉>������c�Rr�	�Y�����V�:�d�M�B_D��,[��?��I%&���?b#lzǘ���OA�Ӂ�y^0Pe;Ң
/�t �5�N Ǹ,�A,OL�ⅻ�vڶ\�O�v�?�eI�ݨ�q���c
���gd|������R��Lmcv��6,eBa��f�3��+��X�mJ5b����ڀ~y#�P�W#��h�v�1Zpǌr�J�P|�����VW�l��<vao�cU���A|>pg`߯VБVOCq8�@B�zvZW�(�a�8��s��2n�B85�E�-�$Sku%0l[5B�XJT��5���Lm(����2h��t��q���K�a��orW�>�Å�ʷ���0=q�G1V��K�#ȅ���u��8��1�rE��k�ظ�s%@��[�33���b���U~�P��"��8n�BԒ�}�|�OD��1۝��anxtHl0�/i^��i� y�F:����ړ�s-��ׁ3��	�6�����_gj��j���U9�LA����xa9���q(Ǹ���{����w�a��9�'��iZ�꫊��f�?��"���~�����E����{� +U����0��ï��������S�jWF��9�t(��Tϩ�\���y�9�����b�庩��2�9m�E�,,K ����$UiML��ئ���l3kJ�v�B���c��W�'2Mi$�4�	#��Rc\�˨��u��0y��9���`t�G����5~��-���ȫ�p�4�ф��XW_�%ff߱S��;�,�-�)fU�A!i>��@�����ϞV�NL�R�b�H��XG�jNH@Nf�9�C��9h�9���Q���KԮ��zU�G�6�:*�;�ru�],M�\�� Yp���{�d:�f�<���F �O�E��_9#kn>�3^��Z��2k�ˊJ��g
�:k9B���ȟ��l��>	�4���=��c�ՂX¨��~�J�E��DO�3�D����j�u�3��­���{C$zX�=ѓy�Gĵ~vh�p/Kw�tmz�R�ws��_n26�̒���^\'�\� J�Ҕ.�SNH�E�rx�t��:Q9t�t�C]X"h�H&M�:Q�-�Z 4n���8�9R��7b_:�a
�ڿ!�@9Ɯ�xB�\
)�U'��#P��]�XϿ�sAP�
�����w��l�ٿq�6��1���O����vЋF$1íF�(�V�N�*5�_������M�X7��_���/e��k�&zc%�Eܰ�\r�_�%S�'�X�\D�7�@�_b�L�Ov�����57�n=q<>(\ʠ�Xd ���(�i2;���^�� �f�MSE�_��=����Z�)�U�C?�P��|�_䥾Ԅ������#�<���7��Ɯ�l0�iHl%\X��-f'����O+Ws��AN.��I}������߸�R5BTtO�����|El�GqFT� &�ks�����3��%�TC�]>�rB�U��q3��/��	��X뼠뿿����j>/�{�A���^�hE��A�g��,l-�ɷzo����\vߖVT���7V�� )� ҭź ^�o��9�����e����긟_���	t*gr!��*N�k<Խ�� ãG�B3���*},�`|l,Zi]{�RaϪ��H��� f1GS��oo���>�<R]7���bؿt�4���*}C`��M�JH�dMi�\����p���wC��؞��o�94�-`�d�/C��C�z[�r>�Ddm��щ�eA���������$*�8!�a��Dʪ�f�:�|��-����Q�̓����̃�]�ʻ�L��˾U�@�la��} T��L�^�Ѣ�_T�N��j4�PDéN����BZ y�{@����M�X��X�֫���ܚt2����H�Y��i��d���0RLs�?���a���v�~�	�N��w���4��*į��߀�p��.5K��G��-�2�N�	�yh�-��Ms��-z�2/a����cݳ>�����5kS%
1��9���(�"rt��.җk�hc�n�|������T�s�4��g�g"���m�1 �}��i�$�ssٰ����J�'�$K)U��ݜ=Dۗ�[c�{�>�F!���Q}���T��;e�a�h�`A���)<J��,Uv�u1N����G��l�S�4��%�-C�=��4Ǵ.[J�T:0�r.d@��eTgɝ:�p9P��'�ɂ�o�G
~��e♀�%S?���hD����ԋ�䊝�ލ�dK��.�3���_��9n�[B�/�$9���n�C�%ܙp���i0�|������V*�9g�c^�?�֦sp�Ơ��)������8���� ����Q9�X\�!�\���5Do� P*7�;_�86�)��o- �ʎ ��ov��S�f=3֋�ܬ`��N�F�!�r�0�����}�PѮKc*l��8 �T�/�R�	B�����P3f('̈́�+:��������u�a��h	&}-b��Z}�b5����2a�5%�sU���J�k�[K쪂�xV��5�0�#�|3�.��/'W,FY�]�+�8��vR>M��
�ӟ����cQ�����V��Ў H!V��Ա:Q����m�L�:mJ ϴ�2�5J� �hsm��Th�u0��V��z��ot�Z����AL9@V8��ٟ���˛���l�6�u��n䎓.x^�s���/��E�1i%�f��D��u�vAM�t�͔e�&%�ub��D`I�N�0�6���{����"�]�`�ͦ��lxl*2�b��^���ՙ��:�^�� ���4����vi`s��$`��l�V`6�����.1�y��&C����}I�"�R��20�^��o�ۓ�����͠�V/�U�$q��Z����	2�¡p�0N�c��r�_lĈ�M���|��p�(k�)�Lf�N��b:�06Z���IY88�(:�k����|ܙ��#E�2��+
�!����*�'s�-�)y�_�f&�*��V��O�:����oq%�C9�`��v�����'A>�C�2S����T<haN�󗂮������8=4'������S���B�|-��<͍���S-ӻ�|9B��J\Qy?-ίq-����Da�����0tQNq�y�nÂWLXU�Cf%^ذQ�b�n�8�|��V D�cŢ>	gZr�2�~x�h�Q=?�	���>��33��7��ѓ]�ۏsI�*�׍@s{7잲-,<����K�_-�|t1�$H2L�Q�I=�\uH�j�7������E�Z��F��-NTT�#?O�c����v�**J�E�%=�b�W/-�A�W��ޛ�Vq�d����o�k��M�Y�/=˯���J9����?A�\FJu"����+Y���ay�B���S�{(1�x&=���b�z�q���Ŏqd�}O��?�NTaT��(��-��q3�H\� Ym�O�P1��DZ/����%?CYkmȒ�(B�����G�`�f���}W�'��3,��yT���y��[h�I
�� W0�!�Ԛ�LP�Rd<b�}�
��b�����=���n�R���>"	/�
V����V�wl����S�~�F��6���y���O�;$@F���+��<�%eY����m9��nQ�p����Tz���MT�ڍx���3YLT[,�+�3S\&X��=��ծE��jq�kj?&L7�9"��@Tɞ����h�P��K6N�t���޸�ALWVQ�$�L��$�Y�X��w�p6E�S�W�:�{�W��2T����_����S%�o��'U�a"��qH�4�Y�4r��FH���|=$����O�jf���\S�VѠi(�� c>���ߙ��*�m[���!Q�e���$P����Ǻ\��d�BBQ�C�P�'!�� ���w�S0���9�\6
cV�������u]��ܤCj:3
JC�ƒ��I�Q�\˸����cI�b;�mr�j�wZ�?��s��y�����1�&8ĮKu�?���i77�AI~e|����Pjɋ�i��gH��ŉ8_y�ς����m�AW�</��h��TR���:���f;���Sf7cմ
�c��<_��NJ\*M�T�O>#	Bp_�H��녫�S�N��+��Dѭ"Ic�A-G#ߩIb��G��9�w/h5c�y��	@����e |�W�s����բ?6����k` �q y�*ԝ6��ЪK:�{%���c��*Tk���K��$>��<��p�+Nճ�w7s�_�0���rh��w�#��g,=1��:=]����L�T�A>�*����a���:179�\:_S�0W�i��ɒ�2����T��:|�~n�Yg���]	>F-�oS��h�N$)���M�H�c�=$�����k�{Õ��pY�@㥳C�wc�w9HVh���Ձ�l��^�
�̽�E��]�@Qɥ[�e��5�"�vt�
XT ��$Z�Ҋq|� ���	��"���j,A>>.�a����d�� �����T=���')<R8o<9B��)�6(2��P̖��n���$����Xm$����? ��'���Jl�n6��]20�T&��J[ĴT ��٨iU�9��b4�	"{~����8+��P��K���>�������n�{t�Cg>�'�*0)�xÑ��~�Y����i����A8��^�ij�n/�S�nWf�N���T.}��
ҷ)4��rC}��*L�k>�rF��e�J<Q�փz�0߻,{�A�2��D9j�J�(�z���v��r�t�L� 4f��b�t3~"��w��Ā��w9K�9���:G�1{N׻�Rݗ^[�P�_tz���$�9�N�����<�3g$�ڦ՚�d��񉙹���/����p�Ļ�	�������B� �"�}��F* �Fɼ�R��8�{=̮!�U]i�Ԋ��J�n�� ���>�t�'K�����M�@:��bΆk-g�1�[���a��!�{'�:��Z�Uz� �Տٴ�@��tt���[E1��HP�#��OQ�bh�x���j�ݺ�2�j� */��8V	.��Vs_އ��@���4C���L���J?gJ>��j|�����u�+ߒ����j����(�^KT��9F:�V����)4�r.��V$��O�Z�3�N�E�ՒS�[�#v��a��k��y�����?g4��aCQzjZ�p.��PA����`>`�a얧 ��(�eg�~3z�e�-�Ⱍ~�x�%�tMb�U4�PK��:ޙ�B�\ ���8o,��]G6H6��SMW/#I�z�`8m��aOC���@�l�[;UX��uZ�\�EC���� �Q��S��N[7�L�;ļ6�3��2݃e��yPw]e�P}��K�D3�B�z,�X�v��mF���7�#�+�ea� ��&Ȱ)�hm!��~��'������%��n5�.6��t�{.0���D:��;��q���l�&����n�np�҆��a�)�_��8:8�c��3� �Y��S�z��oa�U� ��W�LE�\�}�Fs�����(�x`�"�W��1�q���q5q������mH8,�3C�|"���#baO��G��(��KGH��r�f����wSS��N��E�l����fI�1�"ML!Ql	�gx��9SG�t�7�� �X���W�qc�����N@�E�XF�G�+,�7p�����"'��0Ёuf͖�m�� �!�k���"U�ʫ5@B}i�d�}E�'<i���;��S���Bw?Li��"�d���%�B� �(��YV�C�(��zs��{���$��V0���ڂ�����Ў+o��P=P=+N��D4����#�X#�O5�QR7c���V�6����S��}F,l��gt�9���Գ`��8�A�b�e�XD�ح-��2'n7��0��.M[g����L�X���ʦ�w53z^�.-~O�{����U�p�����2#�R�uO�HԺA��K���{	?wل�9�0:����3�������8��h��l8�s�������jA������ы
�<1�D��xјSLsG�g�R�b:B�n�����Y ~��?'��R����Nz���P�%� �5��*ؖ�V�sf���kl����}2�Ȣ��P��=Z�Dp|v�c�$�X�1P�i��
�×��kk����=�<���#6kH
�3�t�YdUx��"5iG�0%���q�'l���Ǝ������5�E���qA�A��{�i�h��9Ѩ	vWg����8���P%�#j�.۠�]Q���4����1ŗ%{i���H���)I��Z�}�=a�cڕd☻3��9�؈�����?<��kɂÜ�a�R�n��AHw��M&�I3L����&*\n_�Uݾk`�=���P����K���[\?���֢�mt]��g��A:5��ޘ�Ŏ�L\�J�A��jߨ[\���{��ӓ����W�)M�v]'���L�U���l�&���$I�k)"/~�`�����ׄG�=�Mϙ���� .2M+%|�<�Y�(�R��Rg�ծ���*	&)̱/��m�c�܋v��g��O���;����.r�m8�%�z���8�$teg�P��
&u�rT���c.Hw3p��Щ���z�-�TNT�by,���	�@{`�y\^3>�U��?m۝�P����`_�nѐ��ڢ�o�\�I�\�t]A�V�F�ģK��=�V������Tv=�h�G�� (���j���������if��C�n)@�E���,SB�W/����Ftd�ȑ��z5m�]����Ec/,ǯ�@TW�t>��I�[ c����֘���V�W oj?���Ą���L8j�<iP�\��ZY�rpa͏(G��N^�x�?�ղ��y�.����,��H��GU�g��O$�s���r�%e�E|��m��)q���ldSˤ��(�jzYd���8���{�}�2�F� s,�R��-� mݵ�<�Z�I�r��
���nϊ�lK ��Rk�:z���^\��K4��(�7E�b��s!�OM?A�Q}�����k���^w�P�"�My���w�Yv`�z��a����X�5���b����kL���w.�/-����9��}w�&�]+qs��(�iT��t�I�Ye��/�-P���Xu��o��X��g�n�1~�0B=	(Bܚ"}r���N�U��=E -�2���@w"@���Y8��%ӑ)�NG���i�W�vi�:�p�؃퓒�`$���1�%�ӗ�zF�c{�3[�z���{z3��)�L��O�F��4V�:�I�S������lI�K�(u&�sF����WQ������Pf��t��2P��6�E�]�cgh�).2F.<tԞ8g*��[>�G�z|@q��>m��H"����Y>7G9+�����k�֕���'����p�@I�?{_�	�d�����H���֓�k�!�
P��t#"��[���I`.�A��U��t���r�K8cd���`��l�Z�i����2���W 7��e����%+{g�uө	��1,".�a�?9��A�G�J�s��j��:�]�8�˚���A�T��z.���1�gɍ�ix����|����ʵ��4��\ �~F���9L��������3[���ωs%�_|��f�Bs������k�j���.`F�q6�	�������Y9 ���Uˏ��U,q˛���̽������6�#�q��\�-c�]N��.՟I-�i�����zg��+.�S���~DN��LB<[|tFi��ݎ	U���>W\�S�����r��^)�r׾8�'��������
ݓU�z-� ���ם���f3S�7�C>r�"����݂AEѼ5G�@ ��̣�K��?�nM��O��W�i��T)��H}I� 5V�w��ζ8v��}���n [Z{]�Z���  �z!vʤ@sg�M�$
�dI!��B��ԊE\b�p ����0�	jQ�wBhP5�l,�Ɵ��M�<_�S@B���fa��zy�Cۄ�(���Q'B�v��q��Bx�>�r�|R�b��;�AG��)��k�H�7�}� 鱭W륟��>���]��1����Þ��"s�;���モZ�l"�~�6�2�$��Ȟf9T�Sf�bw*{Y�a�������F�]�ݬ0Zu?>��wV%�8����,�� �����GC�̒27���=y=�W��n��xƘ@��R᭎���{<a
�kлg�,��(�y�5}���͕]h�~�}��A����k�m���CjEA��H�K���p�p0�ys*�j��
5(>Wx���K.nLZ���Sѓ��*C�����!vׂm� �/�Rs�/�]�?���������R̚7�i��������z�F�)Դ�F;ޛԫ�\K�=������Ӗ�-(�/��k.E�o��1��������p>Η�yo-�,�����ɬYY�`�I��@o.�s�E�TL���z<���w�}�f{oT��ETǎc�_Af8L1�k4XM?U1Nt�O��9��a6E�{���<&E�i��D|pc2Jc���'�C�ɻ�m|%:��Q���L��h�Y�-�F�/x�z��yg_%6���7z�[�aT>3������𾧅��Tͷ[F�(��ho9h�ڄ^�N�>њN?n���dc��ȄȀS�"��$��|�=T�e��󩆻����� �P65���W��TO�!9	�5]�)j��?�^fޅ찉-84������[Hf�Caf�ȑ.�����@�ڏ�N4�1tl+�{�L�Y��QM.sr����߆�����=X$�G�u�*��Y�nhG1�!���+��7as�G����ٴX�8��f��}�x�m]�㑾��׽�c�gj�k|)S[�>��{�@�N4\e5��j�864�a3zS�
I�L(aw�e��v�,5}�E$�����m�'{�C"W�e�C�T4"!c��!&�q7^kǾ���[j�`��f4C;.�R������ [�
������Q
o���3����EAk)>�tl���hw0 2&��>!X��ܯ���C�g0A���L[I#lp�.��<^a�g�%����:>�p69��<�*��=�5(i��a���+�'�R���:8�ʈv�0���H�A�Q������_��t%�X#d��w̆�/�4f}@�达*_;/b)p͆So�U�����N���f���k��B�.�wl�ދf�����:V<F7�eI��C���#E݆9�/�GX���(a7hg�s��'Xa���P�h#�F쮙��W�ud�T�^6(k�NL��v��v%�����Q�`s�8�)ԃ<��n�j�1���4\C3�}D�Qc�Jy1���1����{�R8��i|�O�G�ø.F��@�Д}��-���H��W���B��k~�����K#�-H@R������E��v��� ��\{%q�њ�a�����l,~^���%Q��W�=5*@8lP�"��<�|���-\�H!��^�����O5:^xT抗=�t'�M ������7u��})�-�_6�Φg:Àt�ˈJf1f���b=�nB�P�\� ���9y���(�b'*��D��;I��٧},Ɖ�z�oK�V�UT'Z�v� 
i�� �	|x�E������},��-�a�-��SB�),�o_�?���
p�p2CD_�HA�p���[7>6aV��;����Z�N�ީ���Pk*[mw���:����y��V���+ `e��S�=�k;�ꞔ�ϫE�eR'���!�2��9�z��bĶ�#H ��pCˁJ�w��H���>�>-�A~�G#Z�MF*�������yf�mA�5�t��A���%^[�i��L�>���/6�sMa��8_���/����u%���
b��~{���i,J�<(�!��̭�PQ@�ZA�#�9�7 �eb��3��x��=�ضG?��p��>� �Q��P7F8�_1�/��uL?0���!L���M�[�o��� �B.� lE�)�W��NvZ�(�!"����T�7����'��u��G���
n9�m�
e�YA������v�4�@.��B۫��{�[�x!��Y�����5Lm�/�l�ڃ��s�r�
b3��|"��j:���<����1�^�m}.���s%�O\W�L]�?�X�M�Kg:X���}kf�䈸6��	\p� 0-^oc�������sO90S^���������YO�d/�`Y�v�$0O�����u;�� ���z�s�ެ�w7|�t��K��Q�ǹ��� �d�Û���	�Y1�Y�e�)	ێnt�,��0O;0����+͑��[� 'u�:��5Qu"M Dz&h�I�|ZY���Z��	� �����)�4{�RW�c�+~oա�}\CW�q�\�&�U�e��*�2���^��:;�ح�~Q��@�$�"2�O��������XBP����wP���/|����V� I�=�P4���;\Rl��9,�wh��?�����ƇdN��Ԏ����[���9[C�W�5�+��F�]�*���)4���d� �H�or�$�a��d���|�N���7MC�:��.���"B����Z����{�}yQ 
��>�'twլU��n�]¢b�PE_�\Ȍ��]�P���[�L����O�%��;�3|+.��ݻ������i&d1H�G���.�#?G�`+8o�F%M�i<�o�Ad�*+<�2UQM�i�����ծB��![�$~�Z����A�(��{)���L�6��w��ep��Y��Y+� ���B�ti�}o ����q��]a�޿���"ǟ*���/pp�o�)3;/Q�0��Y���%��R�$���F8��L�Z� ُ	�P���Hk��һ�&Mu�i֑I�Lށ��Q��B�>B�fw�Ҫ��eؕ��2Ē�X�]�;`#�c@�ʷ���6��o��N�s���~l�HU�x"D�>Nz��/�O�(���I-��ۧ��?}���c���w���k<��������s?�q �R�y�fTՃ��jn84��lv���q�4:�s�OSKr��$���=`��x� �6�E:����Z�.%�M=J$tJo�B�W�fK�~��Z\����
��ֵX&��Ҷ#9�G܎=-D:<R6˙|Z�Qm��tk�;�c�0��ծ�5� ��-�!m���2�����������av@s㜬�+'�![�O\��+�_wϰzW���΅�����Զ��+�,a���0U�Zط����_]Uip=�}�q84�R)5u�Н�	ܟ6�=8����B�$(v�Î�P�W|���z��0	v}���+i*��<Q3�@j�o�DL{���+DP�ay��b'�b3���^-��H��Ê��wJ�6)�M�N�����"j ��Ll!r4	/&�x��ol�Ƅ8|U�	f�	��$
*���"�P?#���ٰ�!G�o~�Y�	X��*�7�K��}��U�������x:����%c�y�r�'�����]�
�KFӊ�!;䗍7?��y��Yl'��7Ob;�����`�6���Q�6��O!��s��F��a� ��B��EQz�g��]0/�Z��bp׋�#�|^o���2�a�~'9`��g��~�0�'3��&�+��8�¬�. M��=�)N1���n��X&�A��(d,y�`v���=�)Hi��-i0:9�}4��j5��a.�\���j�)b|S���&����4U�e��>��a"�l�@Z�c�R&��f2�������Č��̎�	�e�t|+���/{nP���g"0 �`a�u̤G�%�a\gf�Lz��U��휝�[�9� o��n��1O��+~(�vm�,c����. �P��#6�?V���Wu���h���U�R�q,v�IO'Ј��Є6!��_��f�f����p�s{ϟM��};}3�+M$�&�}��u�5��ZQ��Gl����J�%�b���׀�0��ک��kO�5$׽�
�v��J�ѸUKw@�o���uO�i�����֘Ë9ժщ�IE�Gp�:��+�^�Z���)�C����"5���2QM׿I?��ɗ(��v�.��?�DM4�H��h�|�V�q�MU{w*�[�}XSܠc���O�+��*���uYQ[F��hV��	[�t�1���	�k:N*�n��m�wsTv�aadrqӣ�"��Mӄ���b�o�P�Y���̓��ƻWoO�@�7Jk�6NZ���h�V�N!�7��{ϙ��(�$RB;�/����)d�4���1����kEb�Y�^���.[�VB�>-2��r����Y!��ԉ���`	��IPI��@��
�Q;��w�?���3�5��D
�R�$`}��{:BkVV�}�B=�$�GT����Hf�m��K8D��P�������quʍ���z[5��d��� �o�E���Tn�Fo5�i}K��e#�JB3��x�3��RLʀ)�e��/��(kf�K9j�����:a!����549 }�Õ�f�|�.6���\��%��?3ⴳS`:�"R�}$~�p ���à����+�:,βf"�P�P�U�C!�8�W��:H��G��e��E���kM�L�W^ZIX[�f�bW	�sdsC.���$4����E�T����y��b�8O�_?�+6ٞ�Y�,�g�vn���مKT�+��jQ�_����:Q+c����w���ؤ�(Jo��M��R"օ�
�j�K�wcSQ�	���z�Pcf���G2w�r�T�թ����.��vY/�g2/�'[���k �g7�O�v��'�L�+<�̃�ßG�+	�bt;f��[�V2_KϮ���|�!F�!�w�f��(5�KK�69�4�g	N�$�W���!,�՛w��n�`�!��Q�$����Ǧ�JG�EZ���q��Ƕz+�B$�:"�
�yMxҎM�S=N�p�R��:<i�=G�dľK�I�����V\9G��7�,��_��fk�('\tX��?.<Im���{��Y�D	�w�X;׶�ѧw > �y�w`��ڶd�)��-��tٰS��P|2)rD���Tb�X_����=)(VH��l�>݇I�`I��Q���+�=Cq�s�Y(��W��A�{�-���\�"ɦZ�L��t5�[9mmL�U�p��7	*���2��<&������۶�`�W6S�6�蒡���n��Ýn ]Lm��������U �X{+2*1������t��r��
�x�W�������Un�oS5L�r���<J��k�;s���e�>κ 3W-=�M�F���&����&���5fK^X|�ŶbR���k���)#�}m���<����ޜɼƩ�	�.裞敬42�UϘ�\n����Τ�k�|���n�Ͼd���7j�x�3pJ�2\�T���C9��&g��N;�-�1s��4 �ϲއ/�k 6=��}�Ǡ	��A��O��_[���xp��ubʿٜ�y$
���4���¡b����l��vk�m<t��E�s�z�ʝO�S?JR����U��B�u^��>�h W�ض 㴷�z��5�DWB��}:���V���v�Y�/�����<��|z4>a8�ޒ����6��"�lm^̱���"��-�X3�@bA4�]҃��7���= �P:B�O���A2���GRb��I�:C�W��t��@#�{��M��J�"�wM���/~ۊn�-&.b��Lw
	�.FV�!�ΐ;�"ϋxh򁷞V^>��9�1hq���i���@�S�]�8��^eﯠк���j�30�X�$xèbu��Љ�f@	�R�K�7�wW�e�)W�)2�X&q{���D����|�����	�?r_Y��	o� �{6n.=�=���	�hn�Ӫ�Dv�K�.S �H��Z�r�yK�hIO��z���Cj�.��,�L�I.����nGX�9��?��a�`rG$�t�%��g�¿��_.؛'�uΫȇ��o��V)*3�f��Yʂ���ñ�N`�rp�<��[�j@r�vAj@�WW����k}�I��v���yD�yF���5�����%��S�6�r�O��ϱ�b}�&���%N%O0r�yM2�Q�rZ�q65
˥#�H��(��!Z��ɧѭd�MkH(��08:��ҟ)&T�y�(��=��T#76G+>^ጋ��\r��������h�`��Zp;%���s��A@�!J�\Ј��h)�R0ik�w��`��btw�� BC��w^����#�R�vI�=+�jƁ�Y@i�s�&���PpA��u�3P�H�m�wXo���轈wA�ü�A�X��+m&���aŏ����T�%%���:�i���vu��r �X�fqj�{CȀ�B�ząJ hj�PzY]����:e%0M�Dz��:�c���|O�-\K�W�X��i\�G������w06������$[]3�@L�s�,CI���k���:���U(8�X��#A�X�uZKa�Vb�)Z�Eb{��̰zZ�}bE7���m`%�A��Td���`������W�ߧ�ǘ�G�8D�k�4�*?ӵ١-�k�$�Ϟ��3sm����}���!��K
�F���v$�+�zD��\3�W�0q�Z�M�W��]Nt>5{��_@��XF�2Oi��A˚c�|�	�.���Ŵ@�tf�^�8f�0���~�w/mʆo��Pa�뽷�29�1�����U�χO
RXD�= .��F�ESx12]�"l5��
��	��Ig��2���U�6���%b�����oN	�Xrۡ~�H(��T�'s»�x{4p��T���YI���E{����O���.q�Vf�ij���P2���"����כ�X-y�^0�
Ra�C�I �/ ����b���d�{��b�>�XfP4q�b9�U�E,2[@�)�z��fv:�A�(d4�ZP�ѿ��r�8�?�t�n�?0���&8�5.v��13/���)�*�E��?��o�B0v2��o����M1�2m�bS2=B��"5�1Nj�$X�t?�. �p�T��"E6���B����X��ո��6�N)��K�bB=r��:����kf۴~u�V9��q��e�D��aE�,&�"U$e�P����J{|K��:.�o^��4_��}�\6s��j	��vD XȔ�qvÔz!������&��f��l~���R�tmKгQF�����˙Ŏ��/�H*?��a�"sґ�yX��;
p���ؕ1����q��h<�*<Нw�o����hK��f��CB���_����A�ľ�z⯍��ǖX��o���ћY��{���*�4�)���϶�K�:IJS�di�� ��hZ:'v�Aӥ���a��V�PT)7��{��>
R�L%��5bh�>c�`�� QV����6�Зeǫ�Xr)�åC�T���V����	yc��v�z0g�(R$� �X�Ο;ͷ�ź�[��jٍ ���ǾF�I�J��Z臦����E O�A�����&���J}1A�1��y�g۶�����.|���bI��	�?��( �鷆8�f�ŨƋ���@L&bOW���~���E}�"��W6��KQ����͓}�},H&�n����dhޛ`o$��������l�V(��7���Xd �l[�z]�+1Q�w\p2���z1b��Z���C	�xqX���ԭ_�����?m���z'U��ɑ\G��kx�z��NW�ګ���7#5ѮM�~���Zd9��8�l d�֭=��Ew��?�q�R�e,��@���wX+���l��+�j��tN	�9N3�;�F�t��X��\�-+َ���'��{Hx���"���N�Z,�Gu4��K��
K�!b_N7}"}�,�( qʋD.�b�����D�U��N��A'/n�'�`��\,�m�����z WC`L�/pJ
�Q&x���58�R�NC�8s)k������*T���s���b.q�؃#��S|z/��ny�+hLN�G�qym�A�3R�?���Z�H@`���A��|��<��8�>4;�X��_ޏ�"��,�g�K�Ck��+Ք�Zpp�！�l*�s]�<Ï����hV\��䈙�r�j~��笑*s�)?V������,��U;ػ�n����,��$c�v�}��.����K�A�t��V`_Bz����[ Z���9� �����\&��PY'Ct��H�(�춱ԴS����Ew��j�#Bu�$ĸ����j9�=��x������YZ��J�W�8��#1�"�rP��:�a���eާ�U6���/�-��]|*N��}��r��E��Z��� C�N��Bթ@�A��L�,�q<�.B
���ǽ����:4�fU]��q��HP��U&v>����� ���C Q��j�x7��k�i~K[d�lE7�5��m�j>9�i�o��ݤ���w��_n��iְ����-W�m-�	�^}��x	I ���{��}U�'�5V�K�i���6Ф�+��°�������.e���i@e���%�][�ʲX�)V�ռh���+>���ҹ�N�M4y���#�
?`�M"�=_�����K�7Wo�):m!��&����xoW|%N��$v�\��GVщ�/A�"_�}���9�,M�8�։�R��AO�AOQ������+��'n��Ɛ�� z:���1�B��]eG�6�2�ֺDZ\0�i������ŭe�����D]c�܍v<�+J>?�|��/E�����4wr�:�Zp�6^���9���0�o��.�!��<�����kJ�eB�c^Ul
�toE��E��C
lp����(�7b��Hj�3;����r�2+�܊�`�� �IpC}E~�=�PO]
��pԆ}�<E���(߅<��R>0��?T���a퍮I�"&Γ���[�P��>q6�
5J��l��Y)���ᶻ}�������#\������`�&�����2�Ӱ����
�S�NGN���(�h�&���&c� �eE��.,��_�:���g☃�g�z�.y�\�x{�5�G��ֱ�h5T�T�h�r�m��T��_Ӣ�z��;`x��A�b�̂��^��$�T0q^D�&��n��/T��=��y�.'d�c�F�iB��w��XD�/6�z��܁�����k0�������������� x�>B�q��3ĠT������0����R0��\�-L�JYj�L4��a=��mCA���[���&	�_rJKቘ�t4TB�S����3�d.�Ј$�K5;�fS�F5z?�b�YU|�
��ƈ����Q�;ܦۉ�Bπ�[%,8�ϫ#�]C�M��=�����R��� ��:E�v�bS!mB�ϿD�\z'����v�g��}�����%�>��~0iU�$�1�Im#=#�p:(:ͳv�D�F�[!�m�h�j6_�n��PA�Ģ:�����UCY&�����4��S+�5qGK�%�I^!��6��3� g�V�XPv�|or ��s���`�?�>�
JfvU<O5���E9T
����� ����h;eo44��f�5��e~\��u����U����)Qo������A�V�k�nK�j������N����:�CWk$���C0��\��O�	-�+�1��������;��Ih��.O!�
��ng;����^"���ޒ����Deٿᒭ�P����v��NfT0���@`��@�;��m4���2��V�`�`�$�o	�|Bz�S3��{ʿ�p�P���m���7Ȝ���)�z@��Z��[�y|`�h�r�P�-�Pb�٫��m
M���.bx�[SJ �u��3��H����4/6��귂��w(Φ�V�����e_q��w��
Z}�	����e�a�U��Y�{������տ��h�z:MS����}�^�N}� ��NҔWĵ\�����F��ިe?��#UQ�,'32�j�R��Joj�l�oI]`��UG��f�����H[��]��~=�e�589��xU�0����������ʧ>�����}�������6=�{R��tHBS����0A����2I ls��yIl�N�̶����?���gXdc�s�b�W)A˟�8�b��o�0b�> G�ը�$�$֭&�ك��fyy�fT�#��B�ۈ�xX��}�.����>HZ�<��qN=R
�y�eDJ�wUH�G��_4�u+k
����b���]x=�b3F�[��p�#83#͏qECm��jTj>���j2o�� ��fWRG�_���a	�p��[PƗ�M
\{Pٽ��G���Nw�C>�'����N�L�_G�2����3���Pu@�A�8�u�C���[3&/ׯ�����m�N���#9T�����Mh�s�[�ĩ'ۅ��2�P�K���yt���S�2�J�pu���7��� bnFh0yז淢�z�� ��L+xm"^�i-�*C����لQ�o�u�#���CI<A��]�֠� 8s9�13��Y�Z��->�:�[�̵a��l�Ssn�άe���WS}�m�P�����P!L}���p�^�IƂ>d�GS�r��ww���#���&�`�����R=l�t����w u� -��i�`��G��E�
7����:�ģ�*�G���i����12_�+��!�����	4�B�_
\�o<]�;�ΫOZ���Bjb�lOOa��'�L�t�� �O�����\�i��H�Q"g4�W�`]T��VlTCn�)��Z��kv��K���{��ړ	���,��� �@I��R��?R�.3qN�����}�
��ޚ��ZB;��|Z�Dol�5���'@Rg�	Pz٭�nx�v?�ɠ���AwW�����%n[��v�N���z��������lbS���R�����܁���������v������nBϥ��Ʀ�ؚ41��_PE�aeճ��J��SHK�a�%�S�q�O#�� ��s�Ǚ(c�`��$�:��wֱ�7IuZ�r���&Hls��*�UoSȦ�h͐F�2���V�#'n/�DJ}���r�yɳ����~N�+t%�v%�PY�U�"���n��\����[`3,7����W�?��Q�ݧ����]�"�b��CwfAh�7	�{ؗF.�i`��X�+f[� cP7� �}&����XRI~��x&6O�R�g+<�[���o��#�?��W4�)�%:a~.r<�;�� ���v�j�������N���R�I�AX�:�@+g'�-�p=��ߕ;D��\^4��Cu�T;|���R9���8n�� ���<�xx���G\7�W�i�����]w'�չ�,�i`oV���dc!�l]�`���'jS��/B�:���tM�
�9/����l�aZ�<�:�Ӏ�Q��!ng�.a��~ĭ��$�,JSb�p�;��ϛ�|��p��n�f���%�3�1-�Aa.D<����F�Z�hM����ϋ�f�t6�g��.smw�+?�i�i�AoO�Ƀ��r\������`�*��
�튟�IL0ȒC��U�Ҧ���Eh���L�ʉ�E2���
�Al'O�%u �ӭpw�+�u�:K��}JH3ki��}�
$/D�W�������*�эl�.�9Nc!w��x(��<�=Z���h���_�Q��k��?Mb��F�7`D�̖{��ӔI�� Y���f�6Rp��DJg�ًϴ�*^��6��:����}j���[̿�P��z��L��̭H3�e'�TS^�%����A���~R���Ô�1���Ȗ��0�v4QA�-�(0џU|��M܋Q��_���jː��26����R/
XN�������q1!������]�'�(C�\�W�Z�L:};*�5��Čɘ?�H~0���?�.ADԆ���s�\�]�J�;dO@e:���VܥDcQ��m�7q�O(��}/�j�ǥ� 	���q��B�i�02\�f���h>���_3��_��sl�T�D�z���+��(�9&���Ƌ-�N(J�J�`@͒�n���S@M��NJIB�QlF�ޗT�.O#h�Na3(�jIՇ;�_s�~�b�YG�|�_/�~�X�:a���g��˄V���L������IB��M<��?[������i�N�Z�����!�!-,��'���ؠ����h_��V�Ah��G�#x�ϏX�'�� _�����7��[�3:�dQ`���6k<!� O��G %l<Q�ê��$]�&+������6Y���}�S��yظ��B�O��/LU|���0շ�3>�dg��9�T�~m�1p������f�l|-������u���?�����(;�:�S�d&ZJPL��
~��9��o�;�I�#0!��.�W�yN*�}Uo>�rBG�Xx�(T�0��cŬD�U9B�G�qF����G@��}��=�}z
�g�����_�J/�
�fP��Bj?�=2W1,���>!$>N6�G�臓�S�_��\�tN����K)�_)�5w��P]̖��ȯ�|���Y��IX!o3���D5^��[D�q��G��Yo�S#	��%^�W���a��9_�f׃褩�;���xi4��a��k��y>t��o���ȶ��4�R�+E�^y�C�[-��������E��W���J<�)ϭ �3�g��gD�%�z�ZZ�u;pc���U`��R�ܚ7?���������!��.VE�-\D���}�E9�c�<�5v�4H��.A���� ���Zhl;���B��.�/]c���%^uN���B�E1[�VOᆨ��ў��w�y�����>��l���%n�B�/�9��3��i��b��j�zl �y���Q���E�W��p�������`�9��Ó;1�@�ˀu��^�,0��S��/>6���Gv���j@�Q�h*�w���«�./�N!E��u�{����UjJQc2���� z��Z�c��kJ�(���)�:%�n�r��1H*�/�?���h'�*Z�E*Q��nJx3[�yh�.$�2�-�І�r��]S0�|G�y0L������>rx �*tA9�{�����N]�J�PW��Ǖ��8%����4D[C�����hi�9٬�(�n�u�Zx>?�x}���ccM8^��N�K.�R��$��iUc�Ӏ�1�fm����1>%}	����X��#e�B�p�j,7#�[ra�؍٩v�Q\D���6��!�m=RG�4#y�k�;��)%
PуYp��8�<ݭgjr��X��ڌ&��(P��Q�`�<}�C0^0~��N�ٶ��ʏ���2�ƿ}ƫe�K	i OZڑ�h�[�����-,T��nT������P���@���w��jy�Tq�OT���R��=���_��;6X�4'�uxH�lC�`+���_It������tx?Yd=������d���ye�f!���H�@I��Ya�e|]�<6���b�Y��DDW�C�D�~��ȡZ;�y�b�5rT�����6v�v��F��9B���n,���ӊ龴�����O,��B�]{�NG�u;��m ��r�a_�r��������g�M�,�U������6�]_#�CcG(�6�E�j��T��TEj�;,+I	�c�_<�v�D�^��E޲��sq�"����ܓ@��.h4�ͅsZ�%o���_�n��f.pqb>��iS�7��%��f�H��Ѿ� >� ��T�@VLza��=h�p1pH|7�ة>��}P5Cet���ۑ'�O\q_B�1M܍��l�e$��H� ��ӣ��Da���G����~^�J�tb�U��1�~ώ����!�A���"�gT3 ��F���M���"A��Go��_��4�7h���{�/ؕA-I[$�q�G0����X�c����.�PP��!��wb���ʮT�1�A����;}�l���.��Kf��Dym>��}m�0��ݧ��-�kғ�@���ݰ�JWJ�]��]H<�cC�M�vHi}z���Y�� ���������g$\��Wbj2&q��W��I�����Nm��L�}��Mm�(���~p���v�t=�ao���v�~��8Ӟr9+�z��ԯ�8-h[�V���GuC�� �&p�VQ�.V��g5���?�@1&���j��ZP�z$`8�e���r��3*FM��k���
Y���e5�uߡk�Q����w�?X�߄�=7�j$�������oI�z�ZS�L����Ө1}P?��*ѐA=�K�w�vLs�Ozw_����s=L����'ߧ��:�#�Si)2^yx~����S�SrƎ��`s�aw���%�'J)�+���-�A���`�cYPq.��ƳJ��D������)w��هL �2�Û��nz�Bi���[(A�a�� w��V��Z{�⽽�}�W[Eß��"Uo"���_K\��@g�G<ֳ� #*�S&9�a�/�2�lQ�=J�5�L�1�R�!�Vzqd�Jk��bo��z�f�p0j5�@	����"�Ϭո�P�De�_�����͈~oO=�`��
B=&���u���f��?�&㲃�zA{��G����
�b+��!@V���m��x1��P�[Ù������S�
_Q�w3�@���"��uW�l��X*�� �������6��bIp�R���K%9�T��85�̠%���K�|�6D�s/b-Ya;��=�:�x�i��>���h�P�,��<�1*�G���z�ϐ��}�
�Şz�	����C�C=\|]F=���üqf�5^�б�6P�k�8����%�і��'�S����M�>���V����~u��fs�@�B3A,�_�jkǥ�l׏mP��y�zs ��
o��*)^;�8�-z�q~�c��r5eK���-	gPA�Z�:��fN4��mtx0� I��jw�i�2�#K�>R �D�Y�d�F�����j2^p�7C㸜_F�	w�/'B�p4�|��(��2��`��]���t9��y�𪭩���P!���8P�DVy�z�E����Q���*-sy���j5b����۵��� EYv����V�e�ݤ��ḑ=��J*����i�\i��� '�����@��|O$B��@��>��Dq<eO�ƶ{���-I	j��yLEO����Tv@��pw���Fv�XJ�?��U��-dT-J�s������K�tL;��ɯDC���X;��I;�o�h�>�7E�s\^(��w�P!���GO�ʔ:��kK��(��"O3Q�=�����7��SH,��EK�Ekx��`ꐃ���'Rz���ƅ�_����_�=�R�"HA\t�����y2��K�B� {�����h����Eq/�pVM�Ε�"�ځ�����b�M�['�M�Y���l�(����gH�z���{��)���?k[�HL9��F�������f�����<�"��R((hޑ���cr�nm|9]�8�G�|�����lyЉ�������ZZ�b�E��Cs�j��j6��{$�z�����7��@�x'�Um�z�;$|o�J��0�Ģ��Ki�̵��N�� �[(`�`h���q���q1\��a�mwr���	1�٭u'a�Ӂ�.2���j\iP�ˇ^6mi�'}�-��7��ڞ�x&@�V��b-�h˹�o�Hgp�4`{��"��?6��گ[�/�i/�kOe`CR�6�q ���Sxg����R:�\*�m=	��/�g���X�A�h��g�@%`��Y��nQ1`	�k��K��O��ؿR��%I�l�D�q.BA5w���ղ��򈔝���:a2g[����}����@3n.��Nށm��׿Ə,m�	 S���7q��Խ�0�
گ���3U�o����UZ "���!�Wl�`bz������E!?�*X� b
���X���,mg+S������� �Y�9���߶A�Tr�`+r�RG�^�Vk�����<u0�<З����h�Z{_;9��j���D<(�����j�鵜��,�T�����f�����),��	�g��4��U�7�A_�B�Q�4X�	��,�D�gE����ڂ�_���?X�����X��c�l4��G�@����8r��o�{�Phf��	�X���"� (́���ul�G��9+�ԟ��H�-��k�������@
�wwA�d��A�\�i��l�ͫ�m��ӊ�)G;�^���N�(g��$_��:"$!۱�y��w}���{������>�a[�][��L��MQ�� ?TP�-(���y
��R8���NO2"����]�G�9�4E��kU��H�'kM�[T��	�%��c*�����w�m��|�B$�1�,q���b{j)g�_K$y'�G��I��\�~p^%4�X�@�����)Nb�Ȉ'�$��*$���0/l���[0������T�ks����3kL\l��=\�nȌtDS�E�S�fאx��}g(�?/��m/ �d�]7ci���	������@w�|hu�]�Y�C�|^s�ԅN�[6r)�~[�W
�����~�b]�&���8H_L���Ғ)�so��x&�Y�~�Jޢ�Z]FSM������i݅f_X7T�y�$��"� 
$pN��� �5������܊�\�\���������Uc�!����r���l~4ϛz��J��0I#��٧h�
��t��Q����!>cS��s]��g��?l�z`'��2�|]$�D���x�P�C����!�o -⤌vPNv
-~h��vo�U�[dD�=��*��o0D݄?� ��c�;g�/[������%n���C���x)`j~[�t%0a5�6�O,�-��!��Z�"���f�D(d8g>e:�P�@)�
���洭g�������ڠ�{K��%S
��>���?a��W΁�
��Ru �2���`��^u�e/��2ȭ��2̣�{I$9�l�v��:��ND(�1!"o3{���y�\�rU�5DQۓ�C��:]-�6l�e<7͗�ȸ�!�c�d���:�b]�A����Ɔ8U�#
�/�FUw���FjO�8Y��f�A�������@||��!Z�T�ZYd����p�t̻�D�F�0���N����đR����p�VX��#�	k*ԏ�~؜��s�"��	]����+�W6�(�w�"�ڹ�8�|�OmF������Ƭ��}<)+:�R&�|I�)½�q3�/��d���|�v�+V��e���`kv6�f���K�>�
[��-�v�{��ۭ�@�[����?ęt����=|B\�n��m�?L����e��� ���vC|����}��'M��o�c�+h�����v��ƙ�)%�v]�ؓm4ai ,��O�ѴS2�%�R�XK�J�p�{���
�T�8�1T|��nB�p�TmT��js��;�Ӝ�b���.�����p@�ウ�z�]���%�/��-tn}����N���J ��~�k�䎝{��o����o�r�(c;[�dS9#
/�a�
ꑚ���'���|�*�*�m�s�ŧ�@^�h�|.��?z�jY��@����/UKW¨�N�"T�Z��e��1�K�>�8w�[P���s����6 ��(	���lq�w��AC	r��ܸT{�J�����Ahh��w^��o��4c�3�)>�z� �D�f�B�+Yr5o�� ���v�8�1����ӯ��� ��nC�\+�����zS$��9E��vB�!�
�;t�_�����>P��V����
<���eʮ�X�cM���lT�E?O?|Mo��F�jO#AAuv_84uTvT�D�e��-�\F�PM)D���2k膞�m�9�9�1����_M���'�=%���WJ$k�y:x��,������t@7vq��}�x8wVVߓ�g���3#��t3'���p�]�x��G��ø��6�✨��\}�2��/>���oUl�F����m�;p�f{���|�X]�7X�4��W�{H��;�j�*���pQ�stZж>��T�3C��%I��̔<���n�>��X
���͏H�����-vQϟ��_���O�
�!r��B���?��F;z�&��<\b��U�1F�)���UwY�8�����B��?�zO��)/�j��D8*��1��	2�_l�y�p��;��i�}�"
�b5���p/uNsC��U�����׌�����ayr���1wu���w���*T]0�O9h2��[�@M���B�iuʑX	!B�>&�⭝y*�!��3�F�}���[��^��Na,؊ŢBf|�&T���2G���k�1�(�o�ضVazL��~cjg���s��q�=$HU�}�z�D>��2�����}7�i�@�  ��U�AN�f���^�iU˼�8��R���4�����ݼ�ި� ��㥕ʻ�4Ty���=���:��]����e�2*$���|�d�&�M�B����2zg9@a��p< �)W��c_#4A@C����<�Vt�ϐ��(=��f4�3�r��V:�u� �*H�efAIu?�{^7�7����"|Ң������=�61@��}�L)��įN� aI{���E�!p
���ڈ�³�2|l�է��J�Z�2/��TyC����u��W����C%Uzw��I&�1��m�f����H��R����:���D��Xf¨�q���������聠SU�t%,L�+"=YAD��N�p�r�j�;' ʄ+�_��B}�����t'e���G>���[q^�u�^�K�ex�6�R������}�1�Gi�Y^�}�>8=��p{��u,ǯ���8v�	VW\I��$�0b7��8��{]y��������Ǿ��{M�`6�կ�1�4׎��!H��� �O�+<:P�^�:���Sj���|�cj�J��3pIAb�-w�C���Ǳ\!TZ��O��Uo��4����&>�QmfiO�:�K֢�Q�A�C"�mԼ�U�,�Ќ#��r��5��Z��/�[��/��,�
�����So.<�����SC�GubY��QP��eȢ_{����Ű:6u+=�a�HC�yl�ϖ�;Wߴe��jp�7�<��mF��������,��(��T�q��Gu�n����QaX���* �u	չR�j~I���^/�LxH�o!�����4L4��Q��M��3.|��)'�*���*��Qg)}�ƨ�!�kd���Ƭ��c�?T�z�١$X�M�Sw��3�!�Us�4:�ռ_���7_���M�TD\X�%�Ϥ���
�Q�U��k����x������"�_w�פ:�+��������m%�K��E�����;�7'��L*�i���������7�!���8[/eܟ�>Z�(�5N�@+Q(C6�}s]��\��E,��$wP����u4�}y�~��$DZεt76�KCZ�3g�bV�7A��{�Gh%v
Rmǐ9pUF��R(�����}i Ѥ'9�o��w���5xj5�4T��l�w�2Io;K$%S"�����c�N
�� v?�~L[Eg�=�n���WX�����a�&v9l���µ}T��_Ͽ����	�<5���	w���ҫI,޶�\��e� W�u[7�x���s� �~E{Z��T��s�]��>��`>Z�ᑈ9SS 4�2�/�,���,��oJ9@�m��6��s��W��{U��qj���4��Too�u�C�5u��GJ7���aɊ�v�#3�Fh Aج�!���Ș�2���?jt�4}�J)̌�m�Ć����~�B�v�C��:��r�=e�9˙�Rd�F���Z3C���8@J�x �Qj��uS�f�>�!ƚ�k�u��������^��BC��%�Q	c�E�AW��c�pgX��r�B����GL������G�&���S�:r�YgN9:z�
��>��J+���2n�� {��Rw/�x�}ګ���m���]�;p����� ��r��хt���`���lV�˥U�!�HKJ��]��� �2ߪ*O��k��{rw�Cײ�d�h+�d�g@C���ʝ�O�����`�$bW������E��omK�������J|�v�);F]�5��O��)	`+�Ǳ���R?\��_8�oǶ#*<�$�=,1��$�dc[����h��8�ӵ�RlŲ�&ZE�`�H0�\��f�hV��Yq��[���@V�����z��L@�Ո�@�������2��K�\7��g�߽����VU���1˃,��%�LI��=Y����J0r``FݳG�|�N�BI`nT�Y�[�c�JF�4�?C��,�$El)"\9�F��WL�~E���m34�V�����D�'�ǻ�ނj�@;��'�?YL�xe~�K�j��{�-�����J@��Ɣ��$�;f�]3H�����1�_��LmZH���O%��RڑZd��Vj�±��8���H�>-=e���nu�(�3�t2��Lh�@�Ti3�VF������t8��:����V�n�����f��׭�;���q����EU���3���Jh�;O������X���R��"����D�M)jΊ�vc�!�S��j�pV��dů�j�T�T����-u�S��=^��2C��d��do��Pb�[2XXɵ�a�ؙ��*��'�����1�H�8C_�˴��Ȯ�Dg���/�9}����G���,BAZ�Aj��l#��+��^+�A��̀��LZ����L��h�O��iBD����_�	��z���:2���x����*���1
�B�>��H�7m�a���Ӈ���ϸ�W# ��k���7�x <��ǸX�zrr�~)���IB��i�2h���RaԸc����b��)5G�p�����g��Ѷ��83���*X$��(g�-�+b.B2J�q$R��j�^���9�FW�Ƞ7oo>#TL�6�nf%��L�:L55�C��#h:'֜T��Ϛj�#*�H��!J)/	����l��r�~�����1e�� ��7��Ben�#���z��b�d����$�x=������Q ���w�aܸб�9Dr��?�z�!Q�#+L]����.���8�m�q��G�q<����]u.C��Q���zg���H��C� �ۅi�PXv�t�7Ϧ���sz� �i����ʽ�y/*�����Jh�u4�l�yt��^��ǡPŭ�!���
*���L*l��/M��E׀��R���}D�N�%����2�-��T=A:#��	D����烐�{���J��3��oj��R2N��f��:��9�k+��$;��Qp'�Eӹ"vx����e�j\�x\��ӌSi����"8�bri��ď+~��D-� ۪�	�,K��d:�ްk���"Oz}��8*�ls9L/�MD��.�Ձ;!���ݡG�O�(��ځ��d!��4��a���~��u�P/�6X�� �\Cx����fJ�՝���ԂCZ�#FC*(�%�5�M$�w��q��ԡ�}P�I��V�2�g�]G�b�*"�e�u\rkN�2&��aX���-XC�|F�]h�p��::��\6�<�d&�۱���Mj�L��A��QRË~]*�Y�����1�k�d����O��r������y?T\Bl|Y�4�����\0��r'��X�h~g��[��`t�Pco��ȍ10㪫A��.bۼ���Ϻ�N]=9Zu1`.�;Ji]maϚ�?�`��`��O�����t��0#�(��[i- ڨ���[�����ݗ2�1���V���{�띪F3i�Zghe�^�x���B�\o���=��%��r}���Q�M�Wk��dN"��n*/4���p5�VT�EH�@=E�w�Pq�H�g
RK�*���nH�ǀC��?$�}�1G�ސeU��\<>�*�<@��2��-ƁM��k�@_�v� .�� �|{�V
+�Nbc�Q�3�I �g����D"޴�w�\�˄ �E ^B8��/�����Txd��;��9H�&	X.��FJ�|��C�MY&B$Gs0fDߪ1�*I�����=�P�ט{��R��_d�Kt�{b9:�Tc+���߷,��-��ٌ]ӐC��}A����D����wćR�-u3��Y߲q�S��X�����sQU���點a;g<Ԙ��t�Ω[�8,m�3ú5�$/���!��japU��.������qK{����]���?j	V�?���*�
��l�[����(^a� e_�̓�܏gk�侚Yh(� ��qF�-�T�2|��P�����F�!$:��e���f���r�0�ҡ��[�����l\j�h�t��1���R���"����`����wZ4Sy���s%~��e�����a��J�H6��.V��D�I�*�V���f��X�2ё��fCM��/�U��|X�T� �D#ر��Zo���LW���c��?LM���I�u3��T����G�Q�i�5[�����_~�Ii��2���+@���E��z�]G&UJ���t�[ך��p������V]��Ђ�渳=���{{����!�ۊ$#oNW$)�z+NO�����h�CP{��k��̹iq��5v��#�Z�$�z{8���X�'�TtG�ءJ:�}�r�\�`v��7y.��B����]��}��bڗ~kdK��e�~_R�b��z�@0W#]0�#������BnBF�#\&��w0�5q���������Fu7C��uū�����j��R��)�&�KC�<�L�d�2>�`QVk�3YG��i\jE�ZSًӅ�v���'�8:OmEC��j�=s^�+�.�gQ���1נfee�M��^-|������U�JiQr�
��hL�$�6�u�c �{��K�ݮ��=�n�#�.�q�e��)�_��ZI�)Bq����|;���4ϹH�ձ�M|o��\�#��K��Z�"F��?[!��~-ma��R�7��W�u���:[��YRL%�9�1��;�+����=TY�]�'ޗ��!*60Y7�ݑW�����Y�D?�X�т��N�/�>�[29�W�;�� E��0�Z<�C=�W�5֢?�q@���^afd�զH����l���Q�`UȖ����@��:.����Z�I9�㷅Ƶ����ﯛ�?�_��
U'`�z��l�b%�5F�a=T��μ������%qj�Q ����1�ӿ���o����#Q��=,�����|�"��W�-�f
>=���T��4l[E8�G�g����<�HP�`��0B'|4~���f��2�.9�iů|x�v�3,��%}�AM,xA(��(=�1�ٝ�鯆��w���'���<����L��L�e���?Z_�;b���Lf2n>��_��[��}�yu�e>���@Vy��T�{��Oԍklm�ׯ ;�+B/���[~�b+�p>��#�N C@f��I�}�\ �Z^�������p�i��|�^�lo���Y��^:6�̪������$ܰ"�,��?��-�
��令�JT!�#"���qk����:�v��%.P��@���O�b�C#��R��r�����(���\��3�ԋh�M����o�7�d��y��s�����y��A5l+v~��D��+�=WĜ��2�㔒�L��M˰���;�s���¬��љP�-Tӗ�x�(^yl���/5
f�.gܑ�J��CuS[0g@~/��5�p�|�
ʀ���mњ�C���X�T�3�?;����/.���<��j_�b�NB�E�^�ӀY�Z�~��a���qOEiÊ��0��0���(D�Tf��IˤÏm+C-���s��j2��@��r	��Z[��jĮq������8Η��F�
�.	�IU������4΂��M�*s�p^*�������$�S\{n�a;���Ӆ7}���K���̠�@����]��i�y��&�@X�o��n��8z��_�F��}M.m����="&�P
��9:�/ V�Z���[cr;���X���Ɩ
	-�����]8�1Q�Z��!���E��}x�T;x��|z4�r�pM�F_J�1����杖��W��'�'H0g��0�|XY����!l�����K�t*�o�I���#v��A5�T �m5��h��§|)ۙN��Z�fE�E�X���˽+j��I)��/n[�����G�ɟ:3��S��z{�sC�̄uv۪�k/i������eE��z��k)w�Х�eo
�w5��^dgO�-��P�d��m�,\�����7�u�V�T����N��x��1�'`�a	��G���Bq��'�O%B�*�	�tmR��Y��eA=y��G���%�I�V%^u
18ޒ]��$ិ)�x��X�XU�5ȝZ�rUt4�:]��3o��,bv����^�C�� �Y��Y�h�w�m���E�&�%�@�R7,��-rh{s��B�}�!Ʉ:(��a���V��/����S3@䡙���`���F�q�-��2�����j���RR#{��؂Ҭ3&��"+f"�b��|3+�،_-�����Y:H)�/U@J{{,�Q5-x_'�ζ�9��j�4S�sF��F�O���e �JNR�t�t�2�@/@��	�E_�����6"���n�
j��F���%Y��b�ks%Be8���q@o�_�XD~�/���U�S[�������"������Pm��������|$=Bs���� I%�kL=L���8���M� ��44�F|�Ŷ=�w��Qk�}r.u͟v��b�#�	�A��d!=  ��#xh~�S$S��r����S�z�v�L.��{r�o� �?��,�V.�{�)�]ٹ�{[|H��S[ܔ�Ɩv�v/.^	�AͰ�&]V�cy�>�C3�2��+�U BC�l�V�vk,4�t����֮��w�	�`���p�O�4�P�'�p\l�pL��O4�5ժM�fE#���@�p��9c��SB��-�}����!�׀*���'�UB��D�!:f�!�JJ�7g��G�jM��DpS/��`_��hz͸Y�1������@���+��őb
Y��0�)�z8�𦥾Xw�ؾ�� �l�xFak����V������SR��)!��(�`���fq~F�R-�$�2q��<k���}g��y�������ka�H�۬�4F�Q���Ϝ�滗���7 �R=Zw���v�p�'Нr��_\־�֩D�H��.�F��ir��%�9�R1�Ғ�[u�;�x�t��\}��Č���逰�]�Y�G �sJ�xg�֐9�q�O�`���#�V`�^��*���m)J�u�S�a�-�_UԬ!��'3������o�G�(������m�x�z�]��bȊ������r�7=�ՂR_��f���j��~�A���=��L�#��ýt�<��4�N�0K:1���
#�~W�N��F
���r��H5�\��8�>^�p����--ZWmK���%Fإ�c�6�ר2��~�a�XڀO����g�Pa���ǈ�Ԛ�����d�N�9e�
�u�Μ����!���oŢ<��~�>�zUm3.58豯}œ�ȓ��#PЂn]~@v蠜7�<�l�l��SX��|��?S�� W��O1\���K]�;I�[/Y�ӈR��N�%J���:^��
��xW���]��>�F��]#�Հ���s�MXO)�v~���
����M-����4�"| �C<��]���F� �13��)~��A��}=24���X̬�$����iЄ6����F����̆���0\���wL�7�����D��.�1�/���KO�l�O>C�7�
h�j���F�3�6e��P����)�N�y�Y�q���w��u?2�>LQ���y�5W�a[fT���O��I���^�5�UW��!�z���%��
G�6�,���۫,�gL!}j�/�žo�p(�^d���]c��ǥ�[�2���ڲ�N�&�t� 0¨��р�w�������~}�1�F4�9�ꌮ�`J>�Z��y�?.k#�7[�0��bc�77�ZJ¸'KFي���ܼ2��?�R<��۩H�f|}��A�_X���u5xK��y�tl�/��7������u�G{��	�SK�[�� 0�����E����7ܩ�.�s�t:�ZK4*t��߰�F�>z��a���\��*L
t'xY,�@H�8P�[*�N�	sê����y�d�$"$�q|�|n:�L)��s��	GN�g���8h����S<_W�f��ʫf�n��?Y��׊>�zn�Y(&�9aW�;��mG-y��YUjK�Lk���I`���v�l���d1�@��S��
�� ���f�j�|� >J��q��\8�ok. �[�0p:�?bI��.��ԕۡ�Y�a=O
N<���.��bZ�nPF�W��s��,�$�<`V��_Q��`��)!7���}UEo{%ј,��r�U�%;ψ	E���>�X��E�wm�ӧ��4�/��X
�$|�7����t��Tl~�$�j�T��cy7d`�P:7{���u��LG;�2�"H���f��k������ř( �`!�b�A�d;��eh�{J��؜�I�r3��sR3^0V�!Ƿ�e�M<��3*�+��藮�������u�T[��娡0�����GD��,���.���}�s}v_��L��D������UB4�\n��@2m�sj�T^�%vK;E��0��R��<�F3�/:Q)�����_ט[/�ͦ)ޑ�C,�^@�P�T�}�����u���>L�D�VC�P:��i:Y��U���[�~4:"h:��"_�nF4��aw6~�|��N[�nm*hQ��v��I[��E��J����)���j��x�Y��R���l��~�Os1�}nXN�>��#�/ ���$ �,|4UѢ?⽅0�=����z����.s��ϷV��le%ڿZ��R�O�5v�EOg�-R��1��%���d�cu�/��!c	�9�U���A<�96�������FDdu�|)4��xw  �����E݅C�|KL�\X�p����^����4�O;ƽ�7��Ҁ��^�
�1���j�GOJWJ�=�w:�r��j��L�z[�V�{B��h�yE(���0��G��W�x��gG�kG>�M��2��&�Ъ�%NˊbW�e��/��Ȍ��+k�R2`{�S������.��)��-�<��.�a<�A�I}�~JՑ��D��WZ��XZ΋���4�6��n`~��AL�����hkǴ���lR,��$n�Y�J�Dj��'RI�]Yv�tM��������V����\�����:�;��dZ-�[lw8F[��>yN�B�⹥�B�����N;��7�f��v^M��L�c_�6�9��^��N�pH�V;��_מ����7��ڍ�JF�0B�^L�g�&ȥ�7�%��աysi����uS����<!��Y-D��(��̖nu�0uaN�
��x(�]�3z�SO�o �,?O�Q�?y���@^4��s����F%�\b;m#T��?g��a��FD���2�S\m	Y����"kFQ���L-������.�Hw���_j,;�T�t��Ri�Nr��B��4�[�'E��T���k��ki��/A5,�� ?*|��-v�ǒqY=ne+��C�]�.34_�a�xgi�1�{G�H���#���6e�*�^�uyQOi��׏���h���%h{xU����6q �.���q��\��!�m��nfdn(9���/h����)C�!2	@Z�
�˄:��1N�0�3���C��3��$ N��蔳�4|���:!(杸K8c{ל"��$Z��H�����_�?T-:c7�Nx(Pז"���?�năw���w�d�<PhE���^w�]o5�Dd{�0'�A��8�k�7�c�}��ŧ�G,���E��Sƈ��	G��������=��f���w>�(�_N�����$�0���e�F�^ln�l�Zxo��W�b�Q��U�#Q�R�����RY2�GD�"��aP���
2�7��z�p,�E�Yp_����`�P���{�#�6q�R^���U���	��Nf[�mz�b'{7�	�l�l�j��������aBW;�b<�M��h�Ť6�}o�o��.��vf��YnU��hS��Fe�UWm?g�1Muq�
e�E�<�M�n�k��L���C�ƕ����vʴ�ھ��G�yAxZ;It �Dф7�ƅ�fY-X��W�i����!U����bv>Fd�֥�R#�d��b%?ea6���q�S�=������b�3�RX}x@p����2~���2��MI�����+׺�9$��Hя{û�{gd;ֹ�*.^m��	�����	bI�x��}�u!������#g�O,ڣ0h����g��9�:������ �����ҊB��
�u<Wa���iͱUAP/J��J7�q�PHu�D[�جnj΢Ѥhx�_�A%8ff[��lr*Sn�ws4[����Qg��t��[ 0�YË��y�Y�J���T�p���7�C�&���89r�}��m���:cw��g��3�9��D�24�����%�aL;�=6�{4��,�~=���i� (�����W�Ow�
St@�����k-�#�us��MT[��|j�E���3q8Q��R����u}��ٔb*R���,���C����U�+��Yr�?w���ʫɦ7�e�iڹ��Qm��_P[n;|x��];�����ߵ�p�#�&�̕���u���?��7|T����0��dY�f���皘�:��Q|W�_�;`�^Ϫ�'�JM��v|s�tzt�e&]�����s	k�'�_�z�x�	7�gUS�ї�G��ڭr"*�g�U�'k�}0�ʖB��!�nb�[�M����G����,9ԍ���P����v��\ˑ�uSJ�ƫS7�>5)5���9�c��2g�e�E�����_3V�O�/Q�L�v�ēu�&J�7�^��P;*+���Q�����2К/H@�:�DPv�R��1�k��b��~�~2N=�$'cb����}��6$}U�*k��o@zC��S����+]Yc�"
XYx%�N��,:�[�0*�H�t��A������}V7��4	R5[ũ�$q~�'�V���IY�����M=v3��AL��A��f��7����+Fe����X9�2�s����՟��:��o8g��LP�=P�3�څ����Q/V���h��!=fY�z���K�`��J��hn��NES�zQ#�Y9��I���d#��G� l�P�{T9A��F��E]���b��/Dxǝ_����5�DJ��9���q�|t4���;&=v�ɇ����bS��𕣶�B��O���a�ʌ�ы�I!՜}�/Xu'W%X_W���֗���n���ۧ�����9})6%a�ȡ�����d�I|s��eџ���h)�c�e�R,�PC��]E� �l�����XlNN�Ug�Nk(q�\��Q�Q``R<t��8hy7i�L�y8��� u��.��7c�G�'l+u̙���Ł!�qu�`ŧL�	ː1�I��Ԏ�A��,ޅN�t����Hw���� xg��.��F�q2�!sBP�:���~%`S7/�aGh�'��S,���ʍ׫�h
KP � �,���IGe9�y����)����!��e>֠��;�Y�^q6�P�[�����ǐwT�V%�ԋ_bM�(;׌���c�GV���Q�W\Zq��Y>2�wv����cI�m�_ ��u�����滐�����i���O=}�'P�1"�:���Gǔ�@?����Ր�_�	b+�r�K2?��uj�t�s����";Nù�>6f�j�wp�%B�`H��}r��6c�����H� 0����}ꢧ$���T"3��>B_#l�$q��~e"��H��O��&0h�U�jZV��8���<��`���c<���r�Qr��zH�@�g'�����!"ń�_�-����Y��Φ�͞ʷ8;�e��V�΃߻T�(O.9y"l=�O�-4�໫��Q�V�'�U�#���~���-�$}���u�N�> d��V|�-X,��"�Ŏ\T"V��?C4�{]9s����&J�^?��hhe�'��L�f�	�ժ'��᠕V��nV��t]��e����+�`ס����) �sX��1����kZ�?��	��@�B�R{M���6'���#SnH�Z\�]���
U9�`ZG�uNlR5���\�\e]�qQIӑ����#l+Gk9�����/�Oɧ��R2�2J�����2+E8�'�X��;�'��{;&J��6��2W�a^����=�q�h5��z� {�쁵&��լp��Fu!��5�SBGϞ�����'Jn������8=Ж�T"���=q#���G���_��#0R�#��I<��;N����B�4͔��~��>�ˋ=�E)��y���.���5$����M\	��G>@����\1�(�9͉������x���"Z`�s���*-Ԕ*��zb�0���ډ����`�Z/xS�ٕk'4�F,d��%�����*���L_K\�O� ��c���J��,��(b�ˆ�3q�����`-`�$��h ���TD�PR���݈.���)	Qy�s0��S�-{�9vjKW�� �����G�؈�A�B�{��T�CI1P�&������� 5oo��ְ,)�a2�#S�W�5�����Sڏ��Y��؍>6d����������K�X�]��������Ǉ_�͋ ��=_=�\��y6Z`*�#/�'��-ը
w��t>��ilJH���7A��E� �F��5z��SN fG�d�!������.�˴�f#Ϛ��|�e����w�%k _�c��n���a�u�X�>�&���[I��;�����cF}Q}6w
�^��WTH���R��^�����t�e���Q�]�c/>�n�C����Hܓ�%������u_Y)���>�mG�-�������q~�:D$�Z"TJJ����0BjB.�I���F�A��+���gt����d8�zղGͽ?�S��� �	j�
7�\����l	r#à��^��>�$&�97a�H������{�����q\d��D
���� ��!+�Aי��U�ӗ=�2
��L� ��*U�y���>D%�j�$"��)�V�R�M����u�U��(d�{�D47��W�3�ui�\B�cu�.k���́��_ �M��sz�X���HA��NhS�'��D{�AӘ��h���\G^b�K;s���|'�%6��l�e�2RsOM��������z9��B*��Mx���!��SL%M��)���:�������x�6��S�eL���=IW<}��)6�o��l[�GNd�o�sa��&�7װ	�<�%��5m4�4�������"Y�ލ�g�1Y�q�3T�\�3,�(�]�7`l����$�����Ћ4����l�����W� �F0͔��1]��&k�@t�K������y�O���/CYXʥC�D+4_V0E��KE��y���d�����Q�۽CsJ��Du��.��m�6�#�|�l��ڹX�}�	C� ��k�����ƺg!�$-�Z��3��[����ő���K��y:�.�4�3�m�/V�8z��VY��T3�+И��{a:� 0đ0�3���9IvՋ����*&����l'Q�:H��͑����i
ڭ�^Oq�� ���\�{�s���Π췫ZW��D|ȅF� �>kRN� ����mg����P�TR#�֢\�Č�IF�uԓ��h�#q���0ٗ�w�Y���5��|�a��Ǫ�I��-��9��7Rq�i�s_�����
��tg���t��}:w/�B�/֢"=�P�f�-����گ�Lғ��pE&�m1��<��y�A���'��6��$lǀG�zm�b�a����QP9�����������ii �����C6{`Ը��َ�u4];�M6�Q�Mq	�C%���X:7Ő.XlO��o1�a��~xݮn�T �cvAJ-�2L�|���c�X��Ş�-��[J��`^�H,�1���V}��Թ5U�B� �k�^��〙}�}��B(���vuh���N�� "ޯK4�PtX�t���XK��~LVK�|ߛ���L�j襯`RR+'���s5'VWQS�X��!�%�x&���Bw�,lɇa��2XSJ�'饮����+���w=�]����R�=aT_�T-\f`�<��7����(;5sM���4�<$�����"��ucMtϢ�*8������ع�8ڟ�3K:L��c~I�@o��*��DA�?n��(�kj�ץ�N���.�j &(�z�u�����M�F ������y�ӻy	���C����܂suH[6����Yy���+���!:;y����Sh��!x/��#{�=]����藼#�)���Eg�M=�D[�_�9�ǌu�32��_���(x�W�[ED����V�MpO��/��
"����½�!�о�RwA���E#r5|�����(Nݤe���n�$�`Q��6��>t-�2���W��H?[���؃f^=
a�])�}H����T�W������
-���޸'2'���[�e�jZM=��V���1@�=+��)�l�
��'��\MCDP	��;�zn�[�@�q��!kU#~�A�0�H*���4ܟ>}�M�>"S˅Tቭ���FCm&�#�ah�	KF��"K����q��w�b4n����O(��4�Ob�FDKHe�/Dx>�������]�����*{����Qƣ�=�����_=W�v��΀��)7�|JxJ܋J��.ŞdA��zPyv"ZXI�߮�~yPko\U�--O�C�U)ݘ��̛�p�}P�a�or�'����|h�4���IYF>iM26
#����E�q?I���֢�}��Y�]�e�n�/eT���
�.��|p�T4�w#��)�z�c�B՝X%����J)=�e�w�M���Ɯ��~H��螓���5�����u��9P���QN������'�z��D-˓��Ӵ=��/��W<��,c��vح9�P�����,[;�2��b���]I�M�M� &��^�^�ߢ�l>b��F2�3��	ͭҷ���c��f�_)g|̝0h�}t1�l7 43���$�y���wq�X$�G�?������.BƔ6@x�f��O{1I2����؛�	G�-7��jj�)�U �?ݳt>�T��^�f��@S6�o^�r��!��+8���^맛j�I&�V޻���E�SzD`uY�N�1	�T��]�����ڇ�-���HM�	����D�.�[�2�dQ�������~�����Pbsl�q��"v�R�/q
ˎ�����\YnY�9�ף�'(�*lɭH���r]���	���S�=��J�o�\��0�)��%�67V;"�U���ܒ�0�¥6dP')��Iz��V��(�J��J��q^$�E��RZ�^�����O����'���ɷ&1�[��o!�$(0���dͮ)���D�j��s��$��������w,��.HeiT��uT�~�å���0�Ykh�з#�;��@��{�y,B�p2S���ٷ�a^��i�]���L���F��֌���?w��N��Ѣ�?�=>�nC�A��ީ����:�����Y��Oǂ�\��Q{��	?~ee�C$B����#2�T���74|���ye��qT\D��1 M��]8�qѲ�S��ߡ=�~m�e�/XnC��G�H�x�'��܎��k,��8�2kԄ�� q��`m���㹼-��_W�@��!*GQ#돘s�d.�0]��"9���v 4܋�z��r�Jb�9a���i`�N��}lđ3Cف+G��C�ŝ�,���)�d?�k��^�^��K�14�׬�]Z��Z���Z��!(��EO�.r�j����ŗ \��+��\j����V�#�Aӳ&�` �q�)����A7Y/%)�9���2q�.���yEX��9�U/�7�KA���ൺf6?��*�%#4�JH,h7�7��	%�p� � :И����B?����&�.Ƕ�a��Hԥ[��N�Pᖶ����=��5��/:�1,�_�����O����)ڊ&�bZ��݅��$���@d�(L�Q�)uG��q%P�P�D||�_N��2\&��w1ׇ8{������Nn�����Ob�A�E+�@К��2���lj��䵏N?��{C6���2V<cͼ����715({�YdU�ޟ�4��	�²�̅��?���b���.V�,D��b��(j��_��~$�J�ȡn=� �x�kv�}u5ljX�Z�p�����S�;���,~����	�41�a��M��}]QC�f>&ۻ��̜Js�,ov�3�8�m�须O�y	T��㬭2�jۈK�`SF�$ '��ø�����hx�m��DJ�kʚwٺX5װ�R87`��3��/��1��y�Y%��7L������.sݹ?��7HN,[�7�����9�h�pzG� ���r��XXi��J)vIӏ���3��I�F��oX�[]��X�8c�"���%*F�X,�:��V@�4uȟ1���z��TǙ��$ �3�-]I�Bq�J����md�����p���f��ZM��c�������b�׫�I���������0V�g��R���[�����L�ue�}fV��2;D�|��rh.[Hk�)�"�l7�Bʪ�X]cQ�	p�M��$f5c���@�f>@�ad9SK�p�Ѱ�|��U��w�F�M_av@���L���RS5�n1�A�`��k�
;��S� ��D�Vn��!Mi�Qh G������Qʩ���o�鑇�,�蔔�c;�	���kl�H��P�4�P+���]�����qLU�ė9'j&5dھE�{�s��]�}F{ë�q�Mhf�a�i�1�5����(���xq_���jĚ �ˢ�o��^��_�m��y1��!���J�rQ:�}V v�Kz��n��5,o���9��M0��c(��<ʎ���%�6�s�ūB��Dڪ2�u�[�dhU����]�=q�81���Y�{��_��`3�S���=$���л�
8�ќ��;_�����.G��I1��%nip�А�֭�x~�P^M
Ӗ��9�M�ʐ�V����Pտ�5uq~ 瀞'"4KÚ��2�6z���%3i�� 8��ְ�VY%-���0��q�J��wA��T������Uגjq�`<�"g�teb��sP_ �{� ���%�o?�	��<n�Uݻ�C`'V�S���`�Ͳ��#U0�P&>j�Z^���VWl���-F<��$����*)����gN�4� J�ƺdC�D�<u%������9ύ���#������.�ϴ@� ص<����I4QOf�n����>i��EKUk�!
t���t���.Pi���p�m��L	Y���so��`h�Oj~
�����7�Ъ��v[��z�%��Yu>�-�I�P�i�<���Ȯ�8�G���ߌ����coR�نI�eU�����Q�ڶ�L�x7q�7�S� �vA��b�{����ټ��W;�m��-��-�6���;���Z�ʑ	�*�k�n��l���Dq�?�S�\P?���R{c�⮅��-��E�E�RQ�Nv
%��w�j���CR!�c��,f��~tKA����J}.K�d��1F�49�?��	@�k�b�.����L���H���(S�Vo�Gn��{x�Z�j@��+�6"���uኞ@A�qӂb�b�r���S@]-�+���\��*���'~�o��[,,�� P0$#�Լ��mm&��z���s�������1ں�L�4�5g_z·	a<��Xy�r)$Ԧ����IAN��.�^��T���������	S��D�M��p̂W�7&? �XU��3�r��A��z�>�f=@�§����v�%BMg*J��ig�`����J�Y�t�]�AM�-���-ѥ�;O:D!6���/��*����#�~lo��=	��6�)�-s��0l;�Jx��a_��U�i�d�+tT5��]@y9�^'�u�1��[��郙Ms�^��O3�G��ⴿp�E,^G�UP�%��bk�Gz����y�Vp~#&��%�������}�vXm
�="+�l �m������V�Y� ��n%4�����l��c�}�kZN�ȫL�ܜ�����t��7CD�A�U�L�4B���n�k;&�H�`7�y3DŔ���r�|��;,J6�)W�K�7��]/��2%��E�Dj.�Ikc��:?t���m#h��Y���B���<�-pчdy�K�@����9���S����T*���h�Zd�٤�����.آ�ն����h,].�>�mr I�
ɶ���><W��W ��:���"M��鱙�����O?D��A��@N����^s���}s��(�SM�ጫ�U���!H�X�IKF~�ƈ��E����z�SD��n$��@a��GhZǈ|��Xա��īr���,���/@��H"K���+�6�]��
,�=�u�"kc��2da�H�������`������ax�J�S�(�ƪJ#�,�(�����L�N~[4�̚':����&�Lt�-���8��X_)�󁰐E�|/�g��dJh��d����pMJ���>� ΡllO���K轉�M�$�4���A�ʭ�!I|{9l4@\�3�����\�c I���� v�/� ��i}�����(�QI.��F�k�d�k�3��Ԋ�bF�]���%H��#Ay�o�1���o��$��OR��]Lf����2��C�ҍ��s{�hT� R��@�-�mJrP�Nɇ��!S���J-]��'5b�#�lO�${�>�p=Q���pm�>����i�~ ���Δ�<��������Ȩ�!*7s1�q��3Ã��N���5�<��f����C�����@���|4�z�u;q�N񿰝d'�����%��k��W����!�?/W������ӳ��u����] ���䴗����]+ڵmM�XZ�&Щ7��~�����ƣD`��V�����Z���G���L�D�]�5;�>��>�xn���k�o�+��Q�m��W�����3�(Z`ߩ-H���F˅��[��]�[�H�=����7�A1����oٌ쨧>�9���ZkL�JX�8����`�3��u9�)�TaάV6��#��/	O��U�)��q�A�����s�6�M��?}F4�8\t ��ؖ=[J�_A?��;m�=T����Ԯ��������0���8`���Pb	�e�rHP�@0�a��$��k�1�" 
F���GkpU��n���U�L��b��}�#j�m��'����ˮ>�N�I�)�i�0�2D�����G��G���d�/M:������Nq�k
�b�S�_�q���M�Hއ�g:*�SX��2�Z���?��=��)ۚ%O!R�qN���{$��Y�aԄ�a�Q7�j+Ǚ� 莮�[�ξ�HO2I�r��$�JC��V��
� vZM('�}'�(aL�xz©Y!�]D����=g]p#���q��6� T���'��!�o9��?�UQ���H$�����C��n��%0��W��u�a)8��3�_�.��fLj9���v���&(b��@��}C<���\>;R�Q-��)�8��Dlv�^�(ݹOS�&^ND{�S���l����9#��2I�\	�'w2'U���.#<�E����SOxt�� ���k�L`w�k��7>��zS�8�w��P���m1����:���%��7	jl#�����Q�f�t!(B����шB�e#����8�������	���FZP4t��~��<�bt�|�{�`����SD+�A�p>i�Iѻ]���iwLn�l�o�R|2��<��<L�����W#`U%�\��Kr�L��ӞD��H���������*\�L���Q�-Iy��=�nXÏ����r��'@�0(�L�ڳ%|}���䊠��|<빖���=p~R��ݓ, �vC�7�����&��*Q�u�d�9Z��d��9@2ˍK=)�Z��(o�R��;���4���Ղ:�K�Q�	mL
��}����-Bg"��nbz�%ǡJ5m����$θѝ��`�F��7���.�&�(׸3J��<G�qiA͒�7������g�hgtϚ-��U��1�r���g�����#~4F�Ӗ��_�u�M&j��լ#���K-e��e�f�G���A�]���J���Uҝ:���m�v�S��
��C� ���/%�-	pBOA!�1���x�ױۛ  �Y�ݓ�+c�|��*�aE�N����'5E���d��
��#Ҏ�]N���ܼ�d�I/�,�*K��.���#�n ]�F��ѽ��Ǆ=IHね��>m��lY�~M\rF�-��s�s��	��@2��u� ��wS��ݧ�F��C�	�wS����)ջ�j��W���X��,�+���3Ɲ�))֑�f�e�,U���a�,^���ǸEM6V<}��O5y8���'T�z�'��Ɛ��Ym(0�r�/`�5`L� �@����ZNV_��Bߺ����5J�#���^C:})K�y0�f��S���ↆ�ܟL<�~U��v�����qR�C)����%6��W�in�$�+7�G��$X�������3&���ߊG@��G���wȒS| ;*Vmn|C���k�Y�&|�σ���>e�â|}�:7b[�p��p~����Ob�!����j��^�a�I�ɮ�[X5���I%����I]�%�H��z�8S�_.n+��%�n=Hg���V���z&���k�j"�D�v[ ��R����}D�,C�i�MB�e��Q��l���ot�~�Ԫ�3qɑ�6��x��gT��u=#�*�K�O"�M_>�vEm�F����s�gG�W�]�3�8�+��ׂ��� �+�4�R)����K��˂��D�[	����Hݗ��H}{^k�?��9���}1��/r`di0�qs�/*�0������-�l���}.�����`SAr%��UP��|�b�#m�� ��_{�ݳ5�x�O�`��1�H��;�V�ᴨ��+S�9�y�q�/�Ә�S��1&�K��i��|�����\paS����#��6�İj�E:B�)�t��/0 �ԯ�-wϮ:���i��m@oj��8��j���N��
���DwT��z~�-�_�[N/���	�s/��T'X�!�8�D�Q�jwӐω��ę� �n��L��ψ;�#�����"xp�[O�Ut3�v��Y/��kv ��	�ܭ���w�䶃�m6��'!:rm�ԊR����*��9@O�_h���%{�J��vh�,�u,Љ�%���N���zy���o4�+��zd^�Th؀�%w����Om��*/�O �m�H�Z?ⴣ��\�oV�T�R8)d�Y602p]�cN����9_���������t�K*ZMsv����xP��s-�T���A�U����7�}GS�f�-
ɘkaG�м�������[ѡb�հ�j.����Wu�H��fx��hfLǭfv����	era�P�1c?�uЇƸ�gƬ��*;QǏR�x�?�=_�p
x����6����0��l �M�tѶ�qk��s��������B_`�,I.�{뮵gv�6��"�{)cf9g�z�NW�)�b�҈_���m@�b1o��;%�
e� �E>,���M�B�Ņ�~�����ΔE��}}��t�n6����`��D�����ݐ4s�F��P��2����IB�AQy�����)��Klpj3>�{�
c�Q���نk���ĸvr�������$�����k&�w�.ڒˀH����FOI 	z��X�}�.z�0A�+	Sf�lݭ��*��Yք%�kf2poh�M�
�U!�e��(��ߚ�o0?��S�`Ni�}
�ؚ\�#����ᷯ�hK��߉!v��t�+��~T�I8u�-`���o#MI�%�T�$����1�?�+8ؠ0"ù�t��H�f�D��	'����`QtC���~�jy�����5��^ʤ�	qJh�фh���O�w�_
:��tU���~Uwnl[�'Ζ��:��������Ja��V�o���y�f�v��,��J{wˎM?�8#����;T����;�/&�j�_��Qwggf@��`�T�g�T�8+�	5��%����N�5������n�o��b�j󀊛;��LA'�ILE3!��oa�W�������/��:'1�T���*�P?�v,1��a��S����I-��)�����������x��Ic@[t�zنb��� %���,H��y_�K����H8����FׁN�7�V�H\�fBw�r�͹|c���J#i�M#2��v���xʏ`$����o�؂;t��w�fEGc��*��/I,e�[}�HŃ�A��z�^j�Rh_���6!�E&��<
k��I�h��'˃�7�����q����X��%E��7�����l��rtƆ�[�X,���J@ץ)����t�[�+��!�2A/W�پ.Z?�P �>�2&�ê��K�A񘩽m���T�z��:"e��!���T�~�rC�s�XU-�Ϲ,@�c[^=�)��n`c�E�����ƍ�l�4�+R�K��
u��K�/W�@ޯ����F�
uS��\����/ߞ({\D+�5��n6nh�����w�a_�a�Xo���pѸ��m>a��! �[�:���uv���@���}P���N0U[Ѩ��9)��Kv��Zgk��JE����2a���>�'����%nL��&�7�@�re�-4�Л#.**����s�D�֭荁Ck��l1��I��Ms�>���b,����'>��	lp�I�T�ح(%��80з�����%�
]��v*?����nI���2F��>[2Z�j�XO����: �޾���]$�����D=���D�P�S�-�+��B�5�Ʋ�*��Ff�ʠ3�?�>�2���jN��q��a�B�����mj��H�� �z=@�4�<�IV�d���PNz��ʠ�A)�"����xH�0^0��M��HJ��Ic�;�G�̃�YO�H��D����t�}�(MCml�����A�.�Q���/���68sc���e������[��J���NJ@������1����I�t����y��_�*䌷�U��JB\Ia����F\�T�2��N�f�oP�8 G/p���kBt�Bԁ�������@G��9�B�y�Z�I������`�j����<�昑�(�?˭\`���Y���A�_h?�b1�7�z�@F�ʿ͖o�4��'(CC�����`���)������;M��xp��"�[2a&l��S&�GVr��O�H�j�O�4(��V�9�a�Z՝K����hs�������ԣ�T��|�������~��5��f*�隚��$vLD �O�ݬ�c��9HA�f�ICV�T3�l����v��&�跭�l�U�UBl"�X��֝?�� ���M�A���$Y�I�Fӹ�iM�f�����X���tl�ɼ�9N1#?Ηz6ֽݱ�w�'t�㐧4[�O��� ɚ
}�Mu�_g>&�������X�c�M.=K���$�x���r�F�S�H�`��W�lw�������Bh$��@. E���`||��33�os�͝�[��%�~��ZD̡�EV(c|���kPu.������T�k����q?1��h��#Cjv�=�|�r�.[�U��HK`��`>�Ỹ��5*Ei���3�h�9�D/��9�m~��6��I�I�>�1��b��-��;�yM��_�n�)Nɗ��ZinoL?��&njdY��3=6�����j�渚��,�=� �
ߥw��|�0Tf��Y��~υg�/�Q��r��"�8
B[C��YM�pĩ�J�
��yui��sp�+�cST
AW���M#�^�;��MG{���f��_A�ɍ��,�?���B)w(�E��7e,
 )�$��7�45�����z�R*�j����U[@�~L�T�P5C�j�uR�MQ��<�U@�d�;Y�V��+I���kq�T2K뤒��T��[?5���v1]���g	�c|k\����M�7vs���u\�g�m�Y�9gjǼbZ5�B<<����'��*����q��
���9��TnL>�٥��K��廞�����V��u��%C��^�/�uFW�|��%i<o�ͤ�u_5��|nҨ�=R����!{S��Pu�'�v7��m�~x¼�Wڶ���YP���q���{�4��VP[dG׮��˄ӿ6�&�ĪK�;.h�)��8M_\x�78'RS�Y>2TmI��8���FY���ГI�A��UD8Ѡ�$*"��vM���K�'���_�(Ŧ0-=�P�� t|��m"��� �����s�"�G�4�[��S\�;$7n��d��^'�㺫C
�I��Y�� 1UA��}���M�V�ā��q76���٢�x����2]�6J�L��]1�=nv����������H��:t�ƚ��U��f�P�WP9Q�)�h
� I�����ҳ�:�XG�l��s���s��5*�)��=����z$P7ߣ���D���z��(3^����JJ�Q#FT� "��!dʦ�P���`uw:�{�e5�lu=b֭�W�<#:Y�d6�i����P�
��>!C79��zye��̿�9 �Lk�7�֝���Tz��#�@�x�%�	��FR���\�ᓂ%�uę�a�b�};p��ܚ(8]rő�J$"�h��#Be�J��g�*�jE>$E˨['cw�V!����J�*����,Yʸ2��a����h��H��f�,L�	����H�(�I��CI��gH,���5�|N�&Ď3"�S��1-�THӾ��kU�v�JN�p���;��[���D��z
^�c ������&��Yd߶η�=���k;�t&�ҏ[ U!-�Q�����P�E�3&eգ5�G;�!�E��*7�v��QMBۈQ��?ڧ��c��GX�B�|KpJ��JOi藌_GS���%�o��O'N�1����r7�f	EiB�QBTܠ�yU�%-H��R\�=p�iΊE��gdS�� �R��_.�9�ʩ��sǧ�*��=��˳_u���q��ۤ�{$��s0�]j5c�7Sz�sʆ�"7�9��4�}�#	H�Y���P0մ��D�Ge�,�.����~
D�ī�K�˚�5��k$�!��dh݈�Ӌ�a�"s:�w����O<�G*y��d>;gn�^���!I��Ov0|!^�kt��4���1��K�1��-�[sEV����;�6t��F~ڱHa��өf��>(�	��FH�jx?�rX�V� ��g���V����Ǡ��L��8��
Cƨ�8~� yMG�ݿ7<Ë�5E�?���!�aT�u#���"�e�R�s-�����F�b����2�2L���Zc�#V��׈#A��y!W7�q����Q#�#��.�z�l�[K���p���đN����ㄣ����yb%w
f�&���G�{5�Goo^u �?��`��M�z%U����x�j|����6U���l���_<�*��y�Ϣ��U�K����Nb'���I��N��bSp�%r	�WH��'���}����'���_]�и�\1G<Į�SH(Ʌ~��(v�P����o�P��p"������a�4��*X�:��g��#X�F�r���p��1������zUZ9�g�۳��Px��/� [�b��Yf��.b%=t�@n��%����l��ȱ��4�ӻ�I�j�s�<�^���#Q�u0�0$�T�4^%o�D4�>3�SA�S{ˊ�^)���r���+	�z�q�.�-�*K= �m�fO�=��E��f2.u���Q���{�Ǒ�ʷ�s�!f���p|�m)��mH�bv�I�KtA��9��� L�oV���_�y;��v�߃\��y����YS�g��A;�Ex�Mr�|�V)�y�Dt��q�L� �?��ܡ�s;��_SS�T�ߺ��m��`b;0m"��n��P�sC#Vy}����{;V�k9� ��#�Q--��c;V�-8������#�:	EL0�9��Z�p�0���;O�a̓-�aФrA"҂��>Y����d�c󦩰w��ۖ1���XQ�/�وj�J��X���6�#�� ���02ߣq9
��P�����sQ�&��%��u�2>��&-�ϗ凮�h|�
C�(���tք|l
�M��{�|M`�?�v�LpZhڬ�(�}G����ŞǤ>C4(W�"�V/Y�L�+�N\n-}`�S���J��L��B�I[ُ�2W7�4(����^x=ntLk��ߦ�R�xr�Jx���w�b���cB�Ǧ䡦�����dm�3���$}��S�_'����Xy��f����n�jj�y:�>)Ts�xY!�q���ۊ���qG��P��T%y(V�'�U�oWU �1o<妟=g:��	`��*��;m
�0��`�]!�V3���] �t �8�ˆ=6��5@�i�
�1ư�b�Fk,W�/��Æ�6H���D���W��.@QCb����{otj�'��_I����7��6IٱE�ڿ�*R���+Jj�xܳ�P82�%��ww.�*�k}���ܚ<G1�bIF�㹵�s�E1��c����"n���!R��(������E�+�0a�)�ɋW�ȷG�^xbL���*�/�2m����|���?Q9��j�cv�95��� �2+�d@�"�'7�K��M�I�BG&�I��+~B�� ���C�z1CR�0�)��u�����脢r�a�MA$�g�^<�G���I�<N2l�� �Hl���܋ ���:�x�~�C/�#Q�)��B�'ӗ�r���=�����;s�["��Q�ת���[��W��:-�����b��/�ӎ5:�N�i>K�a	0Î8���	M���\���(��2N���"q�z�tbMB��$Ib,��x�擄c��5�6����;�Φ_��	:��V�k����y�ɑT�����>2{�\&�5��!������ECE��b�xV�V&HD�4e�^�.�]��X5�
S������l's�!\���*��-m��l��r u�{!S�΢0B󧙴E���鑀��)B+���`Vy�x[8�V�M;��q<%lT+yEP�E����R�,`6�hL���vضI����dI�SGw^�j�<9�3�-�����Y<��1��G`�&�u��G�m(0D�ҥ��3Y���"���}\7­?/W�'C�#������Y�W�ߍ��Z���(J!4��!l�h�d�� l�Q���_�PN4��GH�x������c��\�UE]�0��Wi����e�Q@�O7Ț|��O����ȱd:�D�24Ul���|����^�3G'c(t�;�#�s$�"�j�Vr���
oD�d��!��(�;Z�ژ5�9��eD��3��(NKm��.�k?�I��<!�Z��䀒bE(��>���,��V��p�<bW��~>:���=&}����@;ee�c`A����ٕ�&�ʣ��k�C�����Ǖ��Ȕ���!��
��f��=v@��}8m��kQ�փR:\�AN�c�Y{�D�m�͍��&��85YsUT)X��Um/�c�[[fp�o i�2��RET.�Ց{��5�a�ҕ��];:� �;k�t�Yft�W�$��y+)�o���;�܈T6zs0k�*o����0��˾��YiP�5�]�	Y�Kv*�V����6栗�#9������d�*�	a��3s�k�N| 1�3	GqC
DߌY��� +��Q��c�d�����}����j�i{�+��P5�.�w��4�0�؞��#���pP�7�|�!��R!�v����𚅀�^�B�VQ⇒̉r�Mf�JE�"v�ʟM.�p�o�P�B�Ą3�#[ֿ[^�:��e�Tڲ���˸/�72�p�M^"o&����I~{.�>}d�����ɬ����a!�Z:���b��&
��%J�������X�%~�<�8Uwn��]����B�-�U#8p�j�d�-�f��?�Rف�њ��hp�܇�B��ۮ������R���9ɺQ�$jd���ב��M��x�5R�`�����ؘ0,
����E�'�	oy])}�F�xM�G��s�o"䙶�����\�������/e`d<@͐C�Ή���w���(k|�6���U����44����'��wA�2hqS�wa���(V���Xqo�gY��Dҳ^�>����������ia��R��`�8ֲZuF)<���;#9Rg��-v�nA^@�� ��w�o��F�H�H���40��31�q����tJ�~X��,�Pi᧢Ӎ���<�H�@(&��©$�O�-�G��O��3�T%�Q|^�^L}q�s��ˮ][�������[u�KUA�E�~�%��������\�	f���r���:�+���*���z8%���s�������Z��(;�>yl[��ɩ�[t��hd�}�d��\�"�m\��c��j��m��*�_�*�PD�I9�E4�-��onU�Bi� / �a��--��QD�t��M�{�%0�M�gH�0)�9F�݋;���D�u�ӏ����8�w���=����B�6���BcI_zd��2q���Nw�t�O��ͱ�JMJ��Oe��(+�6�S�Z��{���r
��Ef�B͈��a2�.>���C�����B�XBg��N h=��5ٷ�BS�V�1͐�؉�x�� R�O���H��Ǩ�J�{Q���k�S�E�<�b����QY�rrB����'lC�� ��N��^�A�k����a��,��Se��/b]n<��K*=#_����k��fC��\�N$� ī�V�����y|�_�c����twX���礌5���
aS�X�+���)�����j�J��H�����q�OBv�Rb��L�LAzz-6(]Ƹ�������Y�zs���Y:�Rh2����Υ��?h���
������l�w���`���l(O������C*�]<���]�GxM��"��>UyW�$چ���t<�KU���t/��� ���ޠZqn��}w 1���ߪ]/ͯ�\j��|�X�D�v3��ȐG�d�:�p�`��co<���u'���YT%;ml3��~��A^��/}�=�q�P�o�}��Qӯ�=I��8�ĭʡ�b�QO��v��kZ��:�겑����wH �_�iӥ�A^�R��r�_� X��bx}_��A�^���nծO��8��}�M�]�^m�#b���ֽ�B�Ipy���?�/o��%�ą0S[3��,B��0d��L�tGÛ�nM�
�1t��s��5���V�*|�.(` �U���x���[~�ߎ�ݦ�su���|N�!:$Q�1L�,���V��H��kx�}�.�q^�����@�[����pz��y�')0�aNэ~5\P����ڒ�&�q���o��?DH9���`�trS�H\�`�8׎�b~qm�����W���O�L����Lk�}
l��,a���)��]>�j�-({�\��aސz&�ʅ�h�' ��_�9G2oM ������h6�8p!,�j�]�t񼗁�K�v�Rm�鐣�t��/v����8[U��`�'�+|��m�W5�V4y�e�fH~��r�&��L�N[y�CJ>J^�C�wB돻��h�a;sk)џ�&q��9��~N��S�l8s�yE��y/K�lɭ�}���)n�*9���J'�S�O�!�"0\��IvI7��Yu4NGګ���mf��Hwq\ր�Σ~���͔2�S�/�M"�_J��. /Q��q��	���*��Ax	M%�i;5Pr�(��EWq��ᥡ�N�\)�y��9
wFR]�I]f/z��]�P�	0���$�;�p�ܼؑ�P_� }yQ�p�ۯ'���MF�@4��z
�M��c�ύ����[N��"-|��G�������k)��љ�6|�K��s�G4I�+�{Ψ^"����0C�mM�dq�9����S�b�������:K}@@A�ਂ&��'��r�T��ᛅv��$���4m:&�u�th�`�i��,�Y��7�fV���,��ϱ8���[.i}∵�i�S���R�}|0���#����N�]>`E��Uh��ie��5ҍ9���G[`F��l��{����.΂}S�xx>2��F����H��9���2���mT��	�%St&!1|�
%���F�N���E=2s��s~d�zH����kqj�����|��0iEB%�<h��Y�HowA����z ��+��"IS�+��sNh#��$�}���]V�L9u��־y��81،��6��0�M��q5�F��]�,bO�=�<GDH��+�]��zv�	���������I���M+,N�Z�V���m2n"<^^#����Uf�d�ݫ[����zz�m*٢��t��A0���Ў}��-���������y���>��(�f��1�d�k ��vu�#���d'�˖�1 `te	�*��t�я�����Ma�+�|4���a��\Keɣ[�8�m+��avc�g�H��"��x�5�-L��n�Z֨px:Oh+�=36�9�M��ؙ�wmsWK!�#:-R��_�h�f�0Ĩ�����f�Lc*�,��c�4�h� �ُ��}T�N�w�Uno�h�ۃV��@{<7�C4�0ֵfmV��&ӯ�|���n]D��[f:Q� u���,���g�:zT��q�i\��W�q�V'<���|v���Z��!�!Z����o���	&-�[ͰN�o����]�� )��2�Q(D݉N�p�PA4��V׹F|��ӄ��sk�W�V�ܥ"��b�D��>w��a�"9௼�*�R@/]� ��֙I�c��f����1�Y������V�k���� �'�M��m�����X���:�mFsG-vǃ��҂��K�7КQ�c�P��eI2��b�9��7�K~�������>O�7��\ �^U]_�XC��r�� -J
�m7֜I!��7�Jp�!Rc؉�|ҟ��e��+b�f�$Y���)��eץ�Y�KRqɥ�n�{�&5�BM���bT=��[8�ۋ"G,6b��X���H��.!=����ҦE&2���^&����xa�$i���;��Њ�Co�Q�S���\ԄqB�����D�#ZV᰺��[�y醳c����>!e�er���d�[8H�Ư3�M����^c/�U%j����9Y����(8~�rm}�ڲ?]gx)�G��	�����f 	:��U�7�8�A���@�P��,p,Oa�ɺOWuiX��h��	�����:�e���cv�O+ȫ�T�<�F�((ro*�m��/zoV�-%�w�NHf�q?F�ӹ��l�6	��?�H;N��ڙ�?�9��N�2�C[�A�:o�`r[�!���EQ�++�XROs7{�� � :�׎�h��c�[s�#2�s�-��	�|5`[��f0$�������gw���G���ӧ�J����B:ܢ�)�R:��{�̈́���m�Ъ��y7cL�s��fY׹�K��l��q��Jk�)-
���Ѓ��c6�P���w�NY�s �U��^w�/w9Sk^�9�x���A��#P����������#rTC�d�pQh9�ul���!����j�Xt����z�������nW�?P�[��^��Ӧ 5uDwB��1e,�2�݄g׼m��zf��#h8U�&23ǃ�c p=�fxtcb���W>��YP��V��1�S�wg}Ѡ��)��/}l�������U�#iH�ڮ
������5��m.HR�x���Y���	^Jm�ԉ�oxP�	+i���V���c��1i]%)�L��f���k�sE�J2�n�.��~&�/L���GD��ঙ	|r����\��T
��m����� �E".nlj��ճ"�]��X�+
Y,���F�aV)�k1�+�y9E�n=�@!CZ��S5�	���߇�XB�QI��cZ��eN \�\�I��������,�X�Jֵ�zv�b,�dKR`�T�]�,�!~{\�5k��C&-�#�.��p�+��9�v֎��h���Rb�[j����Ə�*2��@��~k��.wViV�+1N�L��O)�lz�7M�+�%���B���8n�>�=����7�-�S%R$]۹�jNܐ�E�j�j&���R��F�&?���X8>��U~�����Y��4��K��4�n�%M$�>�Q�\�4��HOˤw���Y��[�I���_����/"�7'��ք���5V϶3NŦ���'�ѭ�x���A��j����u#X����.6e7[R2�ة7��A����i���zL2������eģ(4��Ⱦؙ����o���`��<-[=�K�ّ�"��}�9��0GT~@ᡣ�a�G�ЃA�$m�����h�B����Xf�Ǡ�ji���p�Bx�)�cG���걎4q�'��
����#�{�G_Xi8?�]i��z�H�Ŵ=���_xz�w.�w��铳t�=^�V]tg�F�m��`]TnM@׺�G�Ȁ�C2�]k�ҀIf�!aNS%��kj��E��j���[T1�J����ߪ�A����߳$�m�znX�9zh���at,�ۋ����].�2���F��Ewy"I�D��Ī�������E��N��oJ��wX�;�i���@�s��|1]昵fޥ�S�������
�H?Φ*w
,���-��#*I�9uc�v>^w -*�1�����$G��P���5�r�9k����V�z������[�^)5���r+e��".���v'�m!����-9n�rP�K����J{��̶FG�{�hh����t̜#�6Ej,Zv�#Je��mr����Џ;+A�ύq�ǳ3X5җ 82��V�������t7����¸>I.:�;ڸ?F�Q�t�zB��x�����+e�*�5k.]Q��-e�[[b�4 ��8q�Kn�9[Z��W��b�"ᪧ1k�r/�;Ӯ`�_ګ_9�Y's�ɲ!�®�L�}��u]��E3D�=_����pY������-�s��������iC)?)kg?<��ы�~����`C6ޡ>Iз!cD��9Ӳ���v�c����������g<~��[k"��������ύ�u 'N�b�}-��ru��FF�Lw����~��*�:f�9��U���z��Bhȧ�����'�(�A�ƩQ̅��(�0>@7'����m�k�:�)p�}k�g�	\��
��X`9�A���Za�}�Hq�tؤWNv��A�Ap�T^��3�<@�ΔB$�@�ZF`�� ��3b����:��-ʩG�X6�i	�[�i�se:h*��h�7*y]���!��y��	��g�g��k�{��*����g𧓭~��Y$/o.~u�X&�"B����ZiL�`��ە��@�Y�YmZN����V�ue��N`R�)錣t���UЊ�3�� g����)rfX�
�%B��ܕ�k9S��g���J' ��^���3��s�ƀ�X�Tz�t���Q��������n�_���W��W-��Y����� �3��8�z�S��� ���*=R�}J��_g�S?�-Cݑ���Y+ʅD3�r3TE�6��)���w\f��΃�l�߬n�ďS�,^$ f�}�ߦ�!)P����8���]����vҲ=�C�U�A�����"v33����߁�n΃HGv�I�ս5Cf�d��D:76(�5��<+����yJJ=T\d��2�M��C��n�G��S}ߛ�ئ�z�ڼ}�"��^-�S�̯N��n��=b���Y�7��M�z��'��ڑ���AGC�s}_:��^�Fڞ�8�ǒi���&
�a�Ar.�᨞�v�<jL<aՠ�;�v�S��h`<��5\K�lSX@bD��a�v3oN�]���0�U����~o��ϩ%C��/����'[({Q����
��CWG��_���2ò�{~ ��a���2�z�y]O6f�G�'�����\�ۭ�Њ�e�;�g��:m�U�)]Y��'���i�F�'s����rqw�&G��VD��p�a7YZ:cj%�/�x�啫O�8WS��� �,1�����&qMN���&5�;	UA�ƛ�gYxG;��r^�uD�fRK�1�09�5񶿙�
�ٛ ���8Fs6@DP�f�M#�$n����§Ȅ�>NP�ݣ�8��U�����^����2Nע�Ԩa�%�_-���ȉ�@V�Ӆ��oV����8�l��' =���	ӶƥD�����c"�qӌe3%�:��8$,!r��z��d�2�������Q% iO�	�&V���;�Ϟ+��;vpH&���ÂV$A� O{���^�b��f�W)��_6�;"/��ۀ���z쵽^2ze#�1�9g�y�I�:�t�0$D{L�KP����$�� ^�!��00�V��iۍ ��4}�c�e��3R��7��Zg���
%�� rZ��l���ʸ\Y���N����c.�`�nZZ��+0�A>e�n��3��GZN?�%�#��)��&ݳ�ȚS�q����d��Y>�M�-�	v�m|��A��^}�BK�_e��z�_l@8�n2�i,�!ЩCr���=�+�,��FC�"=#��)�}�E�+�'TO����Y	�v��<�����fn����^�d���*��ofE�OP���5����¡Ndt���tܿ��x,��Aӆ�I�{�������8�Ya��ə6�jr��	)���*������קࡳs�ZE��G�/��ג'�6|�>�UV��;}B�$z��l����\;6)G�08�����u�9�����"�c켯H� �q�CD�A`�+��t.-�/��J�)n.���tv�/���\02�׍O�2J���C)��U|��(YZf�Vo�f��?e�����r�QVL\��NN@�����l8*��%L����!FT8C&�5�9�Q n~�)�g�YJ@��ʥ��� ���!����ܴ"��B��A?��uI�������;����M�)
w�`r����ڤ$G)��� �N��Ѡ'c	h�$<8-�zu{�69=.#?/ǚQtK�OW����5w��V��ޥgd6�CU�{ą7�_��O�����&�'����)��ۖB�_Ӄk���B���٨� R�f�jJ&�J�;�0bY����5�ş�7��O�޸)����o���m����X���
���j%Kv�ͣn��MG,J��5��n�%�-Q*��6���HA��G�D���^4��b�	aP��=pV����f���	�����>J��-�D��c�l�S=�"�[s,eڲ������g��X
�q�L A��� ���v���_�U����(�Q5�w��YD��w}ʮk.�_��xux�l�M(��gQ���bw�xE�^t��k��g~�1��kb)�V�(L���zc�����p�GM�Ҕ��iuS�퐉�)���'�~�s]�a:>��Q	���Ƙ||��[��X>%b��T^(���xM� ȞRx�Z ����k�]3+�_���]Ga���4D�p��6�`3�r8���{������~�AC�uZxT:�H��%P\����vD�.1�Q�G��Ul;<T&�ӈKj���S�Gg��(�ƛ'�AD��6�2M-/㱲�'�6W���ĥ釖;J����$@��B&Q42�k��gn��>\����?��*i7��X���3�v���4鼙��.�%hYK�4'5����"��d��{���u�*��ĥ�k�����H��_q�D��S0<(:����� �s5/�?���{p���;�A�A���@ٱ�E^?�*��3��'�&�u��a��I]'],��e�a���}�H���[�3�d!}�z���1�dp��k27�%p�_8onڙk��y��6+,	���$�46���&Il��tv��,ݫ<ȹ
�N=�ܔ�=��a�S�#՟"�F���<�}�+��л�´Oɜ{ul�.9h:�v��b�
��9�򟋴�{0��p7o2�q��ߝ��=�]��y|vG�tl"�Ȍ�K��Y�Je�:r�}��kQ��4��a�YB��M�0�Bn+oLxƅ��(y������[�7J�]^�#����<;��
�q�B���]�Uil}����$ylqM�������:D
O S���Sx6���)qe_�sF���K,|U��
����.wgz9�pr���#�;0��T�㽾,?�a�r,�?e��~���Pd{��cQwa�-%���r4kt����u��D�6�r���>�ջ�1���������R�_��N��C>.�ѝ������������e�QSo�+�h�R���Wϼ�ߤ��l�E�_T�D�9O�˶��r8���1a��D�D�sS��2���4�ķ�z�;O�v�Y�R�$��H�e�*�5�<�~�HC�K=��h����X�$���&G��K�l��w\̮M1e�����Y�5�e���R;>r��.P|��x�$-���f��L���ܼ[S�R�s&�MB�F����Ad�^������*
ೣ1�s�/����Ea�K��KWMf�x�}��%�>n���K��LJ��w�MJ9�C����9|�]%��=u�F�fh��Lƞ�H禉�˯%����7�m�G�]�vKȲ��w�+�Y���E���*0g`�А����g런4����ӣ+�/da�(n W�	?	�Bnm���`h��N�ei�*�tJ�ܖ/�)�R�j��h�<@Aoߊ�D�ש�;^����9h_ۢ��Q��� �V|m��v��A�h-��ܳ�x_���wwƩ��hB�����>!7����0���[�Z��8nP?�EUQq��l�y���b*�a��(ˈM�
g���m� <���}^�⤦g�~�KT��C��6%7�p�ٰCU�'��?|�N_\�_���Кo�����U�P����#�{�c��ۦN��RՐ7g�q��A5�-$M��V�
n�yT_
�v�#�IS�
�&��K5����]���诔��_�n���;K"ᎄ�ǩ�O�=�%�-�[&l�
1���աʥ�.����Y)n%��C�#2�B��kߧ����;9�B���]��j]�=�h�!֣��D6H��Z�bu7�"i��q�A��^�Oߨf�X+l?���x�6�yl`+�����[�g������8�"mQ��]~|����Ɖ%��x8C������&j6�0�+���B��Õtkl������f���
ق�y��
>8e_V93�X��-��ļf��u���M�m��	�3�u�Zx��0���6':�'O����g;�q��ל�픺�mM�Qt��nBA<�Ǻa��3F��t6� �8�D��m��m�]ߠz��L�޾5R�0b!;Y_��E�3��#g�YG�d�Ek��(�&�i�C*���`V��Pڝ����n�[�+0z���hg�$�C�e�~���{�	@�n�~�?�߄�v�$��I�2��Z���=qꖺ�����f�e�c:��^m���:Gܯ=��~��� �\H��Hx������0(	0%DX<�q�O��}9�}�5q5����K��4U�F\w�G���VK���$ganRЫ<����2�}ck���b޼%�d��!-�H޺e����5/x1g�=������*�?5e5��kl����ͼz�u�};�h
��������O�/��/\��tR)�h�$
�@9�{�e�Ju#r�f5����f-J�ad�F_<�ڑS,ۗyw�,�ǆIp|�e5�yjĦ�v�� ��3���#�f��uO�����v��ɳ_3L��!_:fu��a�$�S��� _���d�� �]EkS{[g�]�������研e��8T�� _�n�a]��2����:T]�l���|p�PiF���ѿ�aY�o;ls	�[� �p�H�;�&hck�Ջ�Xg	ٖ��p����[+�dv\��j8m�~��jȼE��1f!1-#���~I�^�Ȟv������'�G�Н����yh�u[>��ZClZ6��7;��&+�20�����B<������I��Ö+��9ޓůV�Fc��eX2B�0v�9�>����qV�b،�a�ei��qYt��s��8C�����e<u,���r�=;A�l�K*@�����x=�oGN�ɍ��㴚;��s?�b�,ܡ����`��M,����{Ϊ3z0�H��^��Egձ��&�����/�	x���~����������N�u�GH�T��1YU���٦:�?�oX�:���4��l����;t"�{G  2���}��n|�Q�$Y1@��*�����JV"~P�#uu:��J�&��ض:�;7��W���e�=����P�ب�<B��+X��3K\}M)~����)&��K��u�[!�E� �U�5k�,#�ׂ�ة!~��s^xS����`���$ )b��|��u��U �f�9��׋4�Tٺ�W�H_{FO��z�d�T,o������0�zq�8�c[��WI��)���H�x�pA"cx�z�̎��k)ϢP�$hG�w5���`�O������kr4�ʄ1�#i9����X��ه����-z3�ӽ���]�K��Hm���W���.�yt�V&��Q�_��o�6����l%�.�!-\��I	�h�f1��J)�V�d��b����K�k��!�Ţ�O)���5~�+���H�&+ ��Iȕ<7t4���Y�JTM�����Fu�\$���v��W�<Gޱ�Iֱ��c�"^r�lL�����dDqs�E'�2k��~b�`<�U�6%�.�vW�S���`i�D����
 ��X���+�sD���>j�%i�� 
o��I����A�[�w1�|�En���ZB\,�=+��u���;�y�Y0���H�jK�"����u@��^�){��S����w�Wg!��Vq����7�'��%$�\��ôH�!{8��o�R�O��g�%A(�r$�C��x�%t�ٟ����`��"#�P^�J(�u&����_�h��5�|�fiW�ii7�l�����O�ş]!]�"Z?N���������Ι��6���ll����],�A�D�rOˌp���n�-�ݺ: r:,��D����7`e��~H3ci&�0�ֲ`z�"��o�RJ?�bnCX_x���<FA�SV���,�xn^��2��\G�dT^�d��{aE
�lBh\������P�>	�Jt`6��#�Us�E 	���^�g��j-:� t$�u��Y��[���͐��0S�]�dL�����$�g�%h(\e������r�Xr���*/>�䳐�:��)��Y�y}��yQwp47�i�o>����N�Z��K���د�㽤����\�v�&F������Է���<<��5 ��I+HN�+�p�T�;gD��u`�_���+ ��X<~��B�[!f�i����Q72e�R�Ԩ��a���nl���0	��Uӄ$�Ȟb��~��Y�:���wBU�w�6D��LZQpS�d��56��[�ڻ��,��cZ�� /r���f^��V�#S��j��w4����p�)��=�±?`�e��f�����B����WF#k�%�a>Of��ܹ�א�܃$Ҩ-�l����LN M�:A��X�/y��{��'o�����3�M3rZ�p����,1����z5���}"����*V���f�m���p�^ޭX0f+��9sd�����Xr��L��ޤD������Ţ�O�e߀Q��щ�WC��&>N�-�n5	�#�Y-�>����`9�!�y�s�������w>L*5d�@��m��`\���.i<LX)��`�i8�C��Q�V�H�|�d��$c|�B{�Z0#�j�j}�\:�f{3|�'yW��EKh-�l��%d�	ƨ��`m�yF�wtq�>h�ܮ!�4ȭ��$ge'���g(��Mp�t�O��p~~���x���e��}� �'(ۀo|�d��Ӷ��$%x&^�1 `��k��G�~>Rr�C��F��?u��]08�l�T�r��B���-J-֐�~�d$hԬ>6��~����q�򅷨H�G�x��S�J�|�*�f�z�5�f�3r}Ƞ?�����	��'r���MĢ�����d@�ꞓ0��!����Wə�4TZ*�N������ZRi�b.�xs��]�\������D�Z�e{���C��:`��i	G�j�Feox�O	��#������<WS��ޜ���)�of��ۓ�r� ]/��G�h64G�2�1k���%�7���'�^ȏ4"�g�\'\0�S�����)PM��0��E���[�"�Q��zb���;j�Ӈ��h@�xc�6�KڼH� �Z�����ü�^p^7C� ����9䡷�Ħ����'c�P�R��I?ʽ_��T�0�����WH����lf��#�(ޙY��3�i�wQ�?K��$��K����h�A{6�����'���0l�z�B�T������hx{�5'v�
�,����9ĭ5��P����ggL��rB=	��ϊ�qs�5j�;�}��_ȇȥ���DK�nvgl� �#S>J �8����-����}���+��G��&6{��\u��o����8Um���m�5p�ʔ���g$ۋ�R�6Y@6�A!YWiՍ������a����3u�ߩ�1�=�5� 6um8K�w�� J��-�@��X����!c&�d��OT�/G�0q�ɾ��T��ŷߤ��Hal7��R����iu4[�b1�1A<}����ܮf(�b6{U���CD����F�}\�΄[�ool��ʑj��=��ML��@%�s=Y�Oi]����"8�����.j�Gq7`�q�~��ֲ)��Y+��0u�F�d���(ݮ��.ɊW����{��K��S��~���d�nQ�ц����u:-�/������B�R�2hA#�<;�x��K �y�jA4�?C��.z;�U��7I�R��HŃ�.�Y��b�ȫ�f����qe���N�ك�7�S� ���:)�=)ZU%E�M]��D����"7�Or{g�RѮ�Y��F�{Pl��؛�gs��Z�'�/�Xู��e���uJ��Qk��o����!�%��*s����gaj#yA�T��\����[	�bC�arw�q�גsl��%�'|�Ņ�f	�7���ZO�UR�%mu�lqK_f�/ +E�����o�B��2h&6X�:e�Ғ�׫���k�L�m��ks����`�����2��!�����*��.�'ճh���=�c9�<,C��")�j�M��έ�w��p��~����`l@p���B8b�@�f�1�e��
��_5�]���s��m���%�B�ɀX�֚|fZ66S.A"D���"x��Af��қCs��-P��[H�m�%i=�z��-)�Ά9��cN�F����Db�KZ琊m�]���$����\��X�����q������=<&����i*�	B?�w�Kp���<�����XY�L��>O� �5�f1��E���i$m��� �
�%��*6��2sUe��ҩ��`	��N����E��uX�z�qJ�������'G�����)�K̯4#���}p������|1���|�סs��L82R�bW
�m����`�y�h+Q=9�M��/���JI�}�Lj�[LB�0]��������4���1�<d@F���G�z�����Ț��h i.�d�v��=i�1��R�?�i�ױx�-`�\Mx��t.�<,�c't��P�.����C n�b��ƌ��6��	��C"B4����9yA����ٕK���u��*�IZS�<�G�?��&�
o�9ģ*�N15>v	M�!�%�;o��"�x��P�n�y���������1<����[�3�������%��._#{T��1�݁�ZȔ�Q;d7�tS�J$#o O���lw϶���j>��y,�)Fg�;ҝ�4��f���>��.��[QV�+QU�DE�BE.#�P��AI֘�
�� ?�����;����s������32S,�GS/��n��:��!!�@��䜢� ����I@�f]���yn�ڴ����-�u�<I�=Z��0���xZ���2��P�a�L% ����V ��@��{������c�]]oI���Ǯ{R��F�M�B$�;�s�DY��^�ێ�=si�s�����+W��������bnq�W��BO,��0�ZR�1�B�c���T��li�g�NHJ��@��!�Bm��~����e(+i���$Պ(;��:o԰!�
3���,��S��2�@RG4���+��	����	�^[��P��%3 R��4������/T�4�(}݊��6~-x��P��1�y�S"Ԋ�-����'?����|$|Jm �+í׳�
%�QE�Y��/�*'X����}-fwT���j��Z��(s�`���B�y�{�/��|�k&Rd���^����|t4�7<�$�8�3%{Sﱸ�Qo����Pfe#,��>�4��ңK_�8S.�F��3����!�O�R��۰�	���
,͋#�8`����Sf�9]��7T.2a�uX�I5����=Ya�>C �@U��h�V/��\���R�ZaVu����N��1�n��=
�ܮ&�(��\���_K�����m?��ӷ6)L��"n�I�wK-������K�^�υ�=S�	��èƯi�R72�c\(>N@0�����n��t��d�'t��/����E�9�6�]���h}���˃Z9�se,��We�"�E.�]��n��� ru8����JN�g��j|��b��Е"D1;�� ��62��@���*4�����X��"7kt��@�6��No�SP�i��@nH�ޤ6��p�'R��ۮP\\xF�Iq_�=4��AYi\�Eel�hw����AQK��ϳ��x��S�bo�ٮ̪�J�N/��Q�7��.�QZ�#'�ץ%^�!��'�Aj��^p��s�-�,�P/ͣA��������������2c�� ;ɡ7�3H�<�TS�$�0P�]6�=���?�p��*��ʳ�>���nq���H���1)��Z�����~�ժ���,��y5���Z���M�Ϗ�6�<��5c���v�����ǥYOt��ˠ&��mKXq���>+U�Wړ�&�d$H�v��|m�V���p�2��/# ��J�չ�Qꙺ(�!Ӻ�4�b�S!��AY�iB��$�tx���� �PS����F�"��zwp���d��������j��v U�d�~;�QR�#��W!���#=�|����p�j�*��d[�"�����R�X�q->�.���3��&dRQ�CD��֌A k�[���?q��~���~#�p�W �Q�𞞻�6���,��%��uͬ��ݱ�7� qt�)6��ui��yZ��+xa5�kF���Y`��Ͱ@'�<P95�3�ͪ�����P�uF����nBƟ�qW���=�k�l�/E��Q ߴ�j3*6�� ��s��YEw�#�oF���ƪTU�
x��<�rI�X����-��t(�&_)������7��i�2%m�H:\��ū�2WH�2���U�h�;�m��L�H���x,��d�D�ӱޜ�;��1\��x�P����[0��Hyq	'�[�s! R���U����ك��Qv���O�@I�JU ��7Y>��v�?2ő��8�cx�a�5��=��k�2a$�LP���`�`�[B���Y�C��>��
t,n98z���@Ų��9�cVd����_��`P����4��� [��՚��<�`p
�٥3�ð��|Xin��@6R=�h)�|#��ud�d_L��-����P�9�B�M޶t�)8����Md3Ȃ,����x�� ?Mj�\j��3�%�"%��VZ�B,m�a[��ןK��Ŝ�n~'�a%IH'�����mW���6y,i�o�A�����/��Y>���uH��S��EgC#�w�^�"��Oқ�?�8]�
�QF�'B�����,t᪐:����38Y�^�n"Ӥ)T?('1���gNPI���I9Ӛ�#?��Ս��zI�Ϙ�ƚ,����W��1C��h���f�fBB�|���pew��v���Ib�Ο�z{�u�ܩ�'�K��'p/�BQ�m��Yޭth�&�O5�[<Vz��BM ��3d�}���Ƒ�à.���"�<6{�1W"Ɣ0	�"����j�P{W�ڸ�g�=�_�w��$A�H ��=-m
:0ɯ?_��`̬;�Z9��[�8�X�	4�-}�6|�/+VRU.'y�Y@�u����)}�B�N� ���G�5��<� �r�g�B�{�}�)�b����SB�+�L�[�M��a�5uC�>l��.4�P�����q��u��
�;�8�nh��8��E�9SK�^f�N��
w9�dxSt@����`�#���*(���d��������ݭڝ�o^��_�F���r (��;w�?��P#H���i�����1�=7�~��aI�4{SZ@���:��X�!ɞ(C>�cp-�m�|�}v��`W���$����6d$�b8�Bh������<ϖ�i5���7Rd{�0s�Yj�ذ��ڴ���Y�%�C|���-�4��t��BI7�&�X?�!|�k&��t���!S�W�a�
�bA���ˠϛ����%�D�t��(E!P=O2��B����v{��)B��h�
��?�0U�pKۄ�N�/�Q[��$���F=9{dO}oh�T~�����@_D?���i+���<��G�.Q#��6L��o*�٫��7��H���&�6��~�;���yy��ʔ���Mµ5�a�'IWM�:�4��ݘ��s��9�`��*�ް��;Q�H;�:(����!�pZ׊ZǫfږPn�����Nf�5���hD)n�i��p��>ʧ'p���XP�%��<����UD*�cd;yھmz��U���KϮq�֎i���.}Ig�A��G*�(L����Tl��;y�>���T�Bs�4e�Ѐ?Z?�'�D ��d�{|O1(�&���?�s����	p:���\&��c�ء��m�<�cdt��QoQI2�PQ�z��L����4R#F_?���e�`��z$2��*=�~��A��EX'g$g�Ug�.ëcNX���2�0c4��4�˫�u��7�2��c,���B�"�X"pv�bK��kIA��y>�,W�����+斃[��0/�T������ra	v<7�mq��� cy
�?��A�'����d͜u֪��r���0jtu�dO�]�^�L� ��}�7�)}y���if=��[�b*����6٥ �;&��ʹ��U��h�����&j]d����f����.�����p�a���LY�k1suG?��қ4	�릪��|A���_�l7���������w�y.�L����U�`NK���d��j��_7x�]�_����N��WK����b������>�X_k
ȷ�d?1.�yp�1��扊�j|:~(4�a�z��fض0Wh 4�M�&�<b����CG4B�����Жc-��;��؟aBI�tB��c9�pc����6�]�n������v�.��_�HZ��#����Mz�O�#K^P�uouusT�vn}�w{*�L�r5hJ�_)_/��N$$XA%��1Z��{$�F��:�����g�E�h����k�x�i�'���m��~����������S���v�v{�;����OI��CK�7��9y�q{Bc:у��.�q��5~V�v%�.n!È�as��Rx{M8�U���ܩ[�y9`�2���ǛY��h�M6���K���uX~���<f�s��ًv��tE8@a&ʎ릣j�U�q�I��Q�U\�'m�=ʯ2��������/�M1n�HBL�c!b������Q9F�J^m�V�`wS{tȒ��@#ж�˗��}vKҔ���¹���\���%zv���ڐ!ߕ�-�5�NS;�՗����ͧbb��)��`n�A%]���܇����f���7�e���eCŠ����P?��<��x��%� ����U�H3��G�h���T�M�*5��M�=*�GN� �/wWW�a:��¶�[�&У"��9l&���=[v�l�sD�6T��Ww������?�I� �'�G�Bv%#X�g���w��)�z#��0R���ozZR
�/rIA&�"�Z�Yi�����σn�c�3�k(3���-��Gf����=z�gr��6�mų��b,�v����@`WYV�ࢴ��� !��=
�����3q�c@^���j���b�]7�G@w�ɺ�!2��	FR�ŃXw(*�__���,�u�3K/���R�tt���MRA]�Ӟ~����	on��� !��v��e���Ze"����@b���cJK�d��H���ܡ�3dQJ@�t��K]�A��2x{ۉ̸z�����0�
�׊ol�60!Y;�}�2W>X�?-��}����p*S��n<���PQ9���G��a�I�}�i2�p]�]�{7�u�G�؜P$?<R�780[�����S�������+�~�bZ���U͢�����2�̢' ��Y47S��iy
� L{X��&o9a��i�����G���Z�>N������O�շ���ό"Bk�Q��l��C���\�_�M�@�&�x�v��/d1:�!���@�p ��4�ܶ��/{��v�5!G�6*%/q��|��OHL���7m���W{#�O��}����?-K�x�!k'fS���5�(MR90�PL��piP��I��s�FFC�17"�NVKE�6��-���dr욚�t�ҙdčpc8�?(�d�t"�� )�Y��[���b�1�o9k?4?�f�� ��ZW�u�xL*(�<����'f�x������%_�o�]�T�NS�6wk�|�-�#xT�� ��u�)�ݧi���]�c:���8��:�e1W�RX�b��S�T3I��KJ�8��q�Xo]�Q��}��߈)�ӣx�� ��P-��h��)��GC1���S�.uI~}��.6ű.P3 �2�@/qH�n�ғb�6z�.�i ��M ��= r]|`��|��7�Ey���1��@� ��}���Ҁ@.�xe4���W����[�.?���Qd諬w�=&�>�̠y���_]Uo-�0�@��M���;B�t���X��=�i�@ �Dh
�O�v�uC��g����b'�I�,j3�{���IOz�N}����x�S�<�A��>���}�8�XJ�!+}�#y��.B3m-�Ji��0�Ԥ�5�/ϛ\�b�0���|q��Y�8���L�-��1n�cN��M'LT�4�:s�<o�=%�v����TQ=�H���s���T�a�9u$d;��d�t��N��=�{?0R�A}��U����>�X��I��+_�H�P9��#�7¿�j2|�A��zHic���ɸ�Fg�6t��8��(D,cI�s �ڊ/4zx(��0�C!��sU���[�
�̎R#��k-���ꂲkJ���H�n��A��3�'?�r3�\7bhG�	b��� ���z��7K�*, E�Ъԏ$�Ұ4��j��8����x=�z�T�
��i�0�󱼁��dpU^�ku���~�S�lq�n�K�B��� �,����{!psG<x�g'�?sH/�$���}�7����{�a(k_�ujS��ŋ�.�i�&����rԟc����b��Z�N��x9��'�7�_�����j��7�X0]�%���C�:n<���bp�1VLY.�8�����2�  �孕z�vN�0���ĺ�Za1'�[��Q~�Q-z�ÿ�_�����d�XCy.��tS��.K�%E�@���x��vX��+ɓ��Vj�tV%�G�Z	}�/a	�]� /��A�7�V�����츆�R\>��t��J�����>%�l��yK�ǅ�~f��*幬׌˴h�[L� ��.Ww��dd��.�\�!_�*x�%{i�Crh0�/'�˕^Uƾ�.��_0����4a2���dh	�ܤ�% �}���A���?�P�A�C��rD�4��z��� !��A�<ԁ����%����c�:o=�7��RT�f	ۖ- �k����j1��OM��D�{�̡�,~b؄�)�|�QY�l�X�X��r$pp��	퐈��!�
�h���R4�=�a|�/eΩ!޴X}�����q@�j�'�"^[l3Im���'nÜj�{%�R�$1�"������= �wC��1��(��G�<GӁu���V�-E�P�ؓ[J�]δa��7@4I�[pMʿn�J��b��Z+stoM�(�]��uw�a�ЫgD��Q��]y{ĥ`t0i�>xt��gLG*���Wpy=(L��Q����FE �M�I���C�6d��Bw�Aʨ�`v:��ȼ�x\�t��AJ����&�)��{鍺,[o,�*2�ݮ�{��[��V5�'[�;�[�*:��Ի�{t&�;;���&8]v�V%d}N�uX����f��d\#��Z�@��v��	0Ux,�f<� �����C�gz�ǌ��P���R��E~8�-��w��T������Zo���R߁O��(W7�,����r\^w����w(��;�p�Yp���E��yI` V	y���ĸ{������
�A:$��e��D�'.�E�H�'����]b ^�3Z2Z_�%��΄u"`E~�V�k��Ƅ�1�ٕ�xmZf�Z%���"���*l����x՞?2hC@j�٩�'@�ڰ@����:���pwv9�5L�ֆm�B���S-�F+O��-ە��0\�]0�s�q��T1�,��`ߕ�o�Ç� ���^�I�f���t�Y�`Iܪg�ސ+�кϔϦ;$^:�ׇ�y�Z�1 &C�����\,�Z�eo�A�/S<?��������ݘ�<����׶y$	���6������$�x�D�q6V�~Ǡ��y�> �KJ�q�����c������E-�� �/�gW(�cI9�.�Q�e.
�(�^|VY��/rV-ue,�"�3�������) ���"�H�{���F����.���M�x~��P�	u-����DO:6��x�qY���G��a�׵<=K0�wS+,D
�����%D?��	�$h;����E�T4��˭�6�I쪊ւwV"��}S�˚��x����3�,5�ʤ=dU�1���t-n%2w�#�5v�����iٳ��[>Jc���F��7�Q���7����%�8����� ��d8��6gcx^>X��T�J�dĔ�)��,�,����x$1 ��ោ2Y����"���K���Lg#�cd)��ݨ�OᎵ�\��k��aʹ�=̙[��09��c�K��p��=��ۏ�۪���:m;�"�9/-t�f�h��+dX�ҽ��W=��eҎ	?��b��Ua�������U�M��TȽ:�S�FBrc��&�u��؛!5�N��0/v��V��O'���8�?�T"�=纯6�3�F�W��	��7N����d%i����������{K��:��k8#���<�O�Dt�~���7��^�HX��R| A� z��}�H(�+��aAI��tK�G炇�{mYEm�d{)B/��r*��q�{������iv�[�o���,��j�M�|���xY0���A[C�=��e��^�~}���gJ�i����e�76˒�Y�Az���hb4�k�u�l���;��ū���o��>����A&a�9AH��Ԍ�Vv!j5��N,b��!#c��d4tLٔ�'.t5�p����7���՜9z{���2y�����vq�6ṣVU��� W!��K ;ɥ��r��G�����9��|U�A)TɘY��nt��DZ�5|��S�u��p����	�E���P��"ʒg�f��-�4c������00c���I�'U�����a�N�����:u=���G��d6�w+E�F�|��P%��"��S2��@�����<#K7�)�l�Ǥ��୓����$X$����[��ܟE���>���9_�]ۢv���k��P�Uv����C2��=|��b�e����s�#�B�=�����L���E3"�$M��u�t^����$R/��$iQŪ�u�3+�\����$�u�L�EM��A�U�)�|ԧx_5%j�9ҩ��������o��8S�C�c3�뿋ԭ��;�Q�~7W��X�]L�>C#��@�J�X1	C�-N μTi�����Q	-��@|��챭%;@%
��9�������{���˨��1pŔΒժ�����ц)�kƏ�"ii����� �\Zt5�B�K���)[�|���u���x�1p��)1Ci�ñ��>d�Spٶ�F��^sJn��;)ʴ�R�Xr���i����-S�ȖTu8;���:�q��Y�D3��s���"=�ʺ�1�3�w�Y�,!�:�F����2;�J_g�P����=��ќx|�R��W���V��������d)���!b) ����q�H�,�;"���}�_Q0�~e�e"w%�����5��D��kJo�?P%k��/	�Gi��jl��z]�6ŧݭ���͌�e����7��x:��Ҿ��3�� |/	m����rX���K�̇2���/��8c�|Ư��ӡ��e�wP���%1}��ew/��U�1&�~�%��b����
J���S�``N�q#��?����Zԏ!^��c{�;�u�P�f�,'u�U�x�K��|��o�r��oX�57�$������/��6S�p}����<;{��o��������\m-����6�e�"p��g`��U�8'�������J��A��	���6���q���9 g�~t�S���sg�.K�WC�y��	���2,>Jwa�����Q���.~�KA%(��v�����?�T�g�G�\ �En�@%�dS��0�OL��3��L>Aa��<C��a`���!|��$�V�h,r���B~�(�"���K,���"oho��S2f-�8J��v�އ���$������[ˏ�%�W�գg[���h& 8����׽ʭ�d�E��[��3{�k b#~˝�[�)�Z�r������"	w�<Z7��92ި���/�����}>*ڂ��u��`�6�RW_�g�s:?�G����Q�1Qi�^�Ge��ƣ�^�sߪ.ӯY�S����}$��f2���!���s#��E���j���[�k.�P�R�y0�M�\	!o�����Ì/�S��P]�F��D�t)�M���N Wj�@�}c�I�U�9����5~�w��T�БijOS��+��Q�iD��۹���0�)?&��V���$��f��N��v	G=F�<��w0S��œ������V����� g�km7�x嶺�-������O	~�c�ގ��Q��366��uN�A��+]�����h�q�T6��vF��%��ј�!I�����q z+J�� D1�f
��Y��t%J�ҕ�ZΥ�>�E�R{�N�<P<�w�u\�G���0Ȕ�=���A���.CO	�2ѤT��+�s��=�Z"\L�'��{�>�=�$O��db�Lpb��+�,��1[���(���_��kHWR������ڲ�d�t��p{��7�)�+�"���f��5�����֏H���jlAK:6�av�5Ǻe��$�.�k�f~�<n��o�emYb�ǈwcl�ʌ��,��I��ŰFa���%2��n���rpÆ����@�ҩʃ��� ���m�Bz�1����
�r�<�48ԴS��������_-F��TT�qg1 v‖�7��o�*IF����.]�@W��nq3+VZ*���)!��n��@�n����8dKe]�Ԃ'��-Ń���5ꐪ+ ��m^J�2�5F�%�|�qi�+�z�AO��g+S1�C���~�?������QpMoi,�u4�Wn�\��H��K����$�?�7u���������P��u�H�u�X,����?� �h~�ǫCb��΁ȘA���?N�MO �3�X~�]�R�l���@��rI�-tR�q),]g0�!�*�acxj��Z�U���[ʚ��hlb�HT��?�6e��Rp�k�q�@h �*���F&�S�6��U�����Y�6]�,���R���wv�.m�L$�>Z��Y�Y��;k,ޛ�$5�}���	4�&�T:� jx�3��uY4sq�9�$j>Q�k��*�!�Mf���?�(�^��Fb^�ֶ�b`֠>���c�;�"�����5����&-��$n4�Rp��tӚ �U�D��!ǥD��F���*n�I��ʃLֈMZr�H򍨳
�/�]��a�pa
g�y\�+�l�W��V$��n�Iy�Q��Jni��@=k���?6��	�'�L���w���ȃ�Gf���?ƚNCy"���a���@=�=�F���;|���r��ӕ0!�rڍ&CL�^���
��~>��=M2y��Z����sΉ��.��Y·"�Td�]n��9�k�`]���hq��K�ڔ����K��wJ
/��(�ү��(�r���%-)�@� �zz�B�->�WE;�-�R�r����t�9V�SO4iJ��Nkh���\ !!�[�@Mg�qi�<�B��X�Jr��}䴑�-^Z�h�LC�N�<�P�S��7i��K���G��Vz�4�9]jފa���֠Gɺ�o�]]+��	��
@lq�[MG���`�a;J��Y��`od~s�%��1Fw$�s��7�6������.�8��Y!s�ׄM��۞���6\^[����O>}h��B����i��{����־&Q@�6��
��C���x�O�Dt�i�9�ˠ{!��O"�f��ů.p ���[d�E�}�����)��*���̆[��#ә �U���2���U5RtF��5OZ�n�d\��ƈ�����f��[L ٬.H�zH��T�����ʰc���U"{���;rٛ��&Nk�#Xq������qXc�%;j�����d7
d��U�Ǒ�FR�(��ۋ�s<�nc�[�7�*�n��.�+O�Z�Ӓ��ԃ�JK��m�p�FU|'T��f|t��S/=}m��bp5�\ǖ���F�C� �E홺x���ҟX��!�(��E�Xz�:uU��F��#�؂��*���,�c��y?��ދE����aa�S��:�s��[F���Xu��$�g��*Wǿ�4��O����S�+�~=�S�����>����o�x,
���:(�]8�Rr+�3�� u�tڎ`���ze@v+D~�|�HT\��X���ʴ"
{$I��R^�g@\�g�4<(�����Z��,���u�S�3&ߟ���9b[)��7�n�M���Ɂ�����I,(���%S��PA�L �j��5Z�CXdѕ�q_�'��=�#�nF�76�& L���8&?EX}���R�~M�!'WO;Qɺv�F���J����\�����7�b�	� �B2v��K����H�uB}�j�!��j=�2�o�9%j|N�=�b�1+
Ѡ������aU�t��N� ���R�`ܖo);�N�� � �Y{�H�	X��8Y�=�h��<x���"
hq)VQ�"!#�}�;�蕙�	Նg�"�l��O���a� ��Wڼ�L"��!_���d��9ْ�{
� �"��漚܅\5=���>]ђ��4��6��M�yu�*��x����lM!SX��YSu�5�v���N���7N����f%�f�1�c(LOqw~Z�bl�Hب=�g�aԦ��>7���L�M���Ϯ��0Z�8W{�߈��!X<Le+Gdk��Ay\��~�`��V b�(\�y����#6g�yyt��m��uG*�/��e�j������5IO���6�(��(i֎�g���	i1�r���Y�e
�ϸ����Ȗ���i)�et2�C����.��4kN�ä&�r�qN����P8��6�p��"�|��r��H8U����-T��Z�ʽbR�yGb���u�
]ڄ���$ e��~�ra��r5����K�Co� �c�tUŪv�yB0���-�Ԡ�Uƪ��6s˭���2Z��ЦEn���o�����h��hu�1�X�Έޏ|k�z.&j�\�w����Z�N�lǫ��sX���O�5p@~&��z�Az�}E$�&쩼Q�	:ff"��:��Z����]ԢN�Ø��"C��[�s`�ZL����m�ڧ���ߒ���
�
V���,iѪ4I�����	<Ԭ07�aݟrM����5$��q�# �L(9D����QkX�65�a��J��t��=��l�j��h�i��]ş0.��(K4l�F�����i����d�p�	��ի+�;��,�u]�k�_�`��U�;V纂�_�O��q�$}�ώ�;�:[�'�8�@�+o����t�-�a��	�Bc`��:��]%�Q:Ry�ͬ�*8Vݳ`l$��Z&#xN�s���#���8fj�3Ҕ�����&�8Ȉ	��,�]�vf�酤����f���Qa� K�c>G��A&�.er-��&�𤎕(�#�H0�-��2��{u��{w���8?�dws f�z��_oa!��&>!��y�\��g�%lѮd3��艟"JC�R�{̖����H������<�ŁY(�l�u
�N�UZg�_&a&�~�̹ �-d��n,��G��*�c!x��mqI5P���Ks�8����a�����������͔��:��4����{�k	�K�,�@M�A��(���͢�Ҝ#����S�:|�� �}}W��R��ů� ��]�)��5��G��6���a�c���,?&T���p�����Ft���/��o_�5*���z8�)�LR1�B�q�� �5`6GDb�y� 6t>�X�q3k�&6pб�g��N}�@����m��\7�a�Ђ��Eb���@�Xrt̆��M:�t�A:	=��)��z��ZY�#�.���J�f\NɄ�.MЖ�s�2#ᯱ�S%"3�b���UtN�l�nfm?��HI��ؾ9�5�	1��R��R-�%c��B�H�쌊
Q����Ew��G���<KSW�����4�xF�N%�^p"����֘$�3V�,`�c81>I���~&)������R��H@Q��VIm�r!��b� �5[|�d�cgwǞ�)�[� ��f?��`�k�Q���9��a�R�!����nIAzHk>@��v̀�Vy�$��sl���-u��v H�O���m��F�d�~b6aB����ѵ[p��ly4_m �ZP۱���O/��R���6_����h��4�k��\����Mo�1����о�w�8<V����͞�����:"��ZeB����D�LRV�5��&���mCkL�z�M܍Z��+�1���R��P��I��k�j>�qxaX�����C�f�>�(�BX:f�W��ĶuF����,7���b鶁וd�δ���넅S�SQ�Mϲ��7++����������S���EL��)��S����eC�߶P��]]*�n12������?[�U0K����Xd�W��>��A }TA�P+�=�����I܏3�}�]l]��Yz�u��m�?��3�iЖ�Slj�T�O�:�y��L�#�f�+�|�jS��&ӽE)�;��6B��3(�%�h�E�Bv.�;�⫳Y[�*cϷ�"B��`�N��w}���c�Vo��2�ڮ��|j&g�����:�fAF��Mx�H�͉i�a�=���+�������I(���*�W��.�On��-68�[ܶu�Ar��'�ͽ�	#��Bu�QO+�K���+��bl��$fn�J��D���3m:�Fq����Mzꖬ5��������TO���˭����qk>�ւg�������gz'�M嵎���:�� 6�|X�.�i��X�bF���z�^�D��	�$h�[��U$����hg��5���E ��@���%�G�T�Ҩ�!��.��@� �\�7�䳢{l��o|b��� 3F.�t~?���u(LWҿ+�hM�����l� ���/���_{�v#����ZX!?U�(�N��6y�R�R!0��Aq��j�ɯ�J�)mm&�:U_���^n7Ȭ
��A��GU�ߢf�}���7�4��yn���
q��/���ܙ�F;�FV
�K�ҷ.�Ʃ�lu\{����h���6E����6�K;T�G�mt�F%f2�|��}Q�=E@��v��0_	X��d3c��8���(h�׈1Nq�eG+�������*�˰dI*�]��(a@�r��N��-ů���nOmk{���q/�����8C��LVt�;��-��WK�v7Le�Y1s�M��uF���B�x��T�5���f��M譗s��J�����+8�j�\:��|�3aOy1�;_֫ݐB��K'-tǾǧ�������a�����:xO?F�iw|F��LPv�i]��$)���J�T��Y��r�7�i������%���?��E�̗��0��L�-Vҡ�ǘ-�'&e��u?p��~������A�Pbڙ���/��1�F��/�����'�D�)t%x�zX�h]՛ ��� �������#Z����$D+&�r�l�aV�]�-H�a Ԅ)n�r��?kh�JI�4�ŌKCkFzL+�5}цH_�n-�����RFټYώ�M]k���W�L6���c8����4��*���[�)�6�N�K���O���/s9-=�HnD�"���'���"�^����'����� �:d�T�mR�N��Ϻ�!��}��I�)���Q���Y�sK_}��$��7��7�6�oQ���4��_���Z�����2��1T#wՅ�ۊq��Gԓ��Ų5�ٓG՜)��S���KM�d���i�񙓺�v�oa����Q�>�
���GKҋ���Z�_�~�oj����/� ��3��a^���8�<*K�7$\�����t��+cgf�c�=�Hp8kL�����rјx��|��"�WJ��p�6��cT������_�����Z/j?m����O����C�&�����'<7�9߳�y��H
���B쥽j�ۚ�uW�O��o�0[�����\���Ȅvz��v"5�V,ίt�*j�bL�����Vw��R- �M&A���K��ܿKCI�t�3��qv�u�5@���+w.�����YzYr�SgHċ�~���/�Q�>M��i-��i�?�_��P"��@pY��<�x\����k
�<���
���v\:���7��[8��_��"��'(@y�m���m���Ie2X�+2��DjP�Q|�R]c3ד��/�t�V�_���ٵ��}5��Қȏ�HԤ���@�}���mtv�!j0�ҳ{Mmj����3��g��$"@�G���5|���s6�5�#��#�P���KN
�[Q�'@���2u�']�؁}M�l���U��w��.���h��:��U��v2�ث��]$��:Pv�`i��܇�8#���7���h��Y0����LV�%���[�p�-�b�~ʻ�yVr|H�#����1r����F1Խ����[6w�����:���0 ����J���3^�=�LҐ�A��.�t<'�(zC�8��6�9F�_{��
���W0Ħ��O�H/�]ȼ@9���'y������T��}��/K�G�ä`ߑ��k����U���ìz�@R|���e��5��d؁9s!@����y��{h@�ɔ����0[���,�Z�4��d]�F����0�l����L���zT�F &�ꓜ�lɏ�e
B��[��V��?r��Ǎ���b5���l$ttV�3������-��8^+m�U~ѥa�k?�-���/`��0^>�]w�1�ｿqX�&�� ���[��0���-�
�ү��ۖ��a0����"!��ʐ���{m+�����z��������esZ<�E�)�ں�{%��~�Q,�t��k|tx�����R&��Y�&��b�I@������v���ܢ��/F#̐�E�p���ʠ�
}½tu�"�ɳ>ؒ M�2g޿`�E��?��#�Rʁ�K�,�JI�<c�AB�@(�
����iqҪ�c�����][�rgwph���&�x��V�q_t���`�`״"�eY:��DȤe�����8{��/���LڠD%��"�Ո(�9��W[#Ί�D��Rb�@����3�mi���0���T��~��הxfW���Ͳ
(˧�JA���Ȅ ə@��^w�:����y(�-���@�'�h�T�ڜ>�+�98(���q�lc��o0Ha�k�C��� JCcVm�v�-��g��Qe�(�#?�)<���$���� \ц�w,�ڳ�W��6����Q�Z�B����4�����z ��hJ��9�b��9X����s6������,V����xx���S���H�z����]g��� V~`P6{���%� ��z�������腑��z�/�E�17]lW ���E��3��FW�ü�� ��|3�^�g�ED�D�9Ux��x�0�펝��D}���pe���G���\.8�P���B��?�hډ-�
0<��L2k_���`�I�i9���;5�4@3Zϓ�.]����a�O�bO ^J&�w��læ[�pcꡉƊF"�����q*#L���bV�e��ף���r�#����ʕ0G���hs�p�m���/F�`�o�jc��YI�}��	��;��dPB�j��v9�Lg�y-��g�uc����K�o�ā=�ޘ/�i C�:[.SZn��MU�O$&�W�	h�۫�b�l}��j	)��өU�~�ÍW��ՃIWb>X�t��N�xtW���M"�[���"B�׼�Ǭ�����A��K�xˡ�)���ןgj��r�/��} u����8���� $t���G�H�(��z��gl|���L���D���t���Q��X޳)�� �<�Qzi[yrUH䍃��%t�k=�B8f���Y`��6��rb/z�T�Z�c��ZlZ�/,{��O��Fx�GWpN!7VqŘ &rY�W�N��No���"�����|� �^*tW�7��� ��l½TLj�*��b��2]�<v?z�>6?۷�,1kW��;yk=W�����`	��bF��|�mچjc.�0�Ӧ������±*Y&�k���Zbd����Jޜ�,haK���4�R;Θ��\)�"�����?��lZ��O�I	y^p��g�a�9�nԇ 	�E�<Oiw:2^6����S\A©�����ƻ���n��[F͞C"�#0n�x�*v�-��7���D�&���(#��f���r�F2��=oO�6"bw���i��
']zә�����P����o7�-�L��j�$:��n��,��{����M�g�%�Y���RE��GN��֭`^��rd��4Y����u? ����؍-+�i>}z:�Y�Cj>��,��o�ژ�|�%�� ��.��:��7��,�l�B���2�7��v��M�E:���[��y�cA^�&�"0%�x�ܟƉC��܄^��J�c��#)7�<��z�nK@�=����G�V��2c:L��c��Q66�޿��9f�G�1���K����[���Yrh��E|\9�!Y=Y	ڧZb%� ,�'�u�I%\�B?o�Ny|�9�&���@��D�@��^sF�ŇL��j�HA�?��,��S�C��9bG��8�9�a�>���g���Ԁ���{
ע&E|l���->w_ ]o�١hβ��/��i��Q���/�T��q����"��w���K�Y����[_�0��&��lX�s�Uj ��U��E�%~�v~��󦱹�tړU�h��@���~�R�����Yz(�=/`d�>{��X���_�B�wf� ��O=ubxŤZ�������o�%��|L*I���벝C��*�J��}pe9�
<�7��ͮUMkU��:t��#�-E�ዮ���	s����
����}��J��(�}|��Q�#㬞F�lS��
:�l�M��1(UO;h2#�v78�p���bC��ē9��1t�s�[�
��¼��7���٩�;�}5��~�tY<_7P�����np`m��Cj���d�ݑa| �g68�5j;9A������4��H_��=v�ۜF%p����@����}D�]�!����9Tӝ����8���,a �O T����bcx@����D4;`A=�z�܊d$:��5iÆ�V���NT$Q�@\�H=ƚfº�������1si���$���?��3�+H�������zf��vW ���Ӗ��O:K�-�m����w	��X9V~L�'��^� TɎ;3ť��{Ss���Ze㍲��u�k��^o4	���G��$���ºj���b�et2��"m%)�}L�=%��3��c0�[�*�
�-��s�M��Y�\�ٚ����H9�e�v��+l�鿈Lِ_˼�o�!�ɶ(6���� �(��=�W.~�����/���d���?�]p_�qo���Z]�&C�n�|G?������-������!׼� �cm��Ú($	N��E�L�����>c�K�O��Cܒ �c4���SV�\���09�:r� �S�|]�qc��0)���7��Iݑ���-�Q�Kc�l1��z�[�j�{�BsM��6��ֻ�-�>a��c[:Ɯ�`m(� ��x����?��^ �4:P��6���y^ -fLR�Z���>1�;��1x�eF��q^'�FMv�Fe���<��n����a���p���ֆ�T�h�m�mA,�!~L*� :���;^d�$u^>�=(,Z�J���Ha�i�Pc�݉��V�3�י\��衕	�:��Z�rz��*�
�0��L~�W��\�1ds�y��6 ��H@�&J%�.p���l���taOvZǌU�c����%�@I�w���T�=���m���~9�y\ӠN4DB.Nm&Mϊ>����QL\�{>R=���W=�D��B�\(=�;K�iܟ�d��-6h��ߐ0 ��HA���C�l9aF�,�>g����N�j4����d��y�}��{M2l��8X�%_��<��h��f�Xqgy'�fh:�iEZ�h�=��!bQ%��I+�6*.Q��<��e�VL@���%.osty��D�h��p�s����Z
�i�ܳ��&���'���L�H']�L�����Eб@�&P�+ҳg.&�����u ��j�d�5u�)! F+j/ B��g�N���T~,�=��2��ĥ���pG ��+�G~��2�bvچ��YR~�3����U�@�a�V�ԙ�|�%Xh�l%J�Zȓ9�S���.~�>*�;��t�zC<�r���%�,>ƨr��N��ye�+F�{���>�����Gs���3|�#����h��`.H�B)�_��\�~��y�b�u��'�&%�d�~N��oW�\���M�Z[����s�d�hB�� ��2�wJ\�k�+S�l��b���_HA�����v_1��P	P��n��Cvu?<.}�z|�+sUİ��LQ�:w�bݤǛ�z����:�w�$��� D����5��&G���:�s)�]��d�_�l	*U��O��.w^� ׼v>7LL��(�&|���?�'�\�e̿g�!��&�"f���K����=��jb����YBC;%/�������u�M��s�1���[K^������E��,@{����6L6k��)�����\�@<��#E��ϤW�τmOi�y�"����g�U���Uϣ-��p�<*G�F"Z����"3E�g ��w[*���C�� p"mH�u�����գ�.�ݕ�	���O�_�A��ܠ��^Ò���+��	9�͆p��O驉d��.��<���h2��F�lm|�#<79='o������6Ψ�T�Wa]�0(F#�Lrܪ��e߹�8��誚��DP��&k��Й;�H�}�J����^ p����Q�f#�|������oj�[m��b�? ���Y���+3�^�=�Gp���]���a������.?8p��8�w�������ry��}R5��b��HPΠ����y�C��db����f9��`��8)�԰�u�����`pU7��]\�iJ��-�Vv,L,T�k������4��Wy޵)?<�� v�"��h�3��|��!��!�#���u�'����/�ΤFG�nˬ婫�&�l ��8���ES�x�a�D^�� R�bQ�#�ut���uZؿi_
^ֵt���p�sk�6����i|���]����K��#
e�"�F~b�/�i(YV���U��T̻nT��1� ��Z��1�K�s�&����A˄���"�G�N��3u��ȝS&0���H�����Y���ϖ����n�u&I�7}=Q�j��Ev.�,�}_X,�L�e�c�c�I���*�Ό��X�SUjo++��%Ha �t �N R�=k��@���D���&C+��@ +r�G!x�,�M}��c^��,'� [��+�n@>�Fl����fɣv�{�Nb9 �J�)L�u����8�U��:s=r����.IP.0n��8�
���](���̢{XY��e���Sc.|m����TP����+Yi4e'�����]g�3����!n4��L�@F���������ˌuZ�umG�e񤬛�Jw����%]�YI9���v���=����F(Km٪�!e�������+��!i����zu��4w�&�Uk��[�� p-ߊH:'�g�ċ���*�N���VyJ���O����1��q��ňH��b�����TO�)RK�9�����>M����#_/|eM�E�D�ml��Ry�-�|0����4���}UZ�:�������*�����Q�z�R���pa y�-��^.���i��	M~�*��E�H��%]tq2��uh�f��d�0BSr����\/!�A]�=MA�J���Һ�ܧ�j����읨����{�����إB>d�E {w:h��M�9\R!)%���F���D�-RA@�-J)ӽ�#�N��aW\�/�C�\=bM2f7�u�>��)d��'s��eÛ|�m2�D�E1�� ��R�z���ʡ]�:�v�C>�z���S�%�h���%���UNomU��ħ>�{O�
�Z9m���zU��4�?�b�km"~!��@��&�E��]����6��:b+� mҡp,���5P-�Lwq��5��56��rƘ�Hu3\�N=\`���~Jh��Tܭ�8�c>�b�E!G/��Z�����=�`�U�Zp�-�~�*UΓ|z_@.I�QQ�-5��
 ��a����C���PVV��ОsF�*%���hURQ����4I^H�'hY�݃,��i��4,���{a�Ş�"�b�7��%�!~	g(���%�r	��@d��JlS.�R�x�颛A4~���r��zh]0���~����U?��'��4U� `�(��dտ�#^�i��o�`�n
���>SV{��"u��b@�RF�e��V�u�û~��Ż���ۭ/�oK=�bZ�]k7�'A�0d�ё��H����$x*�i::2��E�NB_�6�s��Kp�g�j�an���ű���~�C����6�J�J�����*���#%:����斢?�I�y�r;J��$\�K\�Ȑ~dł]��٘s�xdC�ƕK�hU�U��t�Av9�׭ӠF���NP9�ŝ���/�Ӻ�}��e�M�����~����A��W�[���U�4T�Ke,�l���:Jſh;�X����x^�{?���V��~d2�y db��a(U��f��'Ů�<�������OM�1HcG�K�*��V���谊`q��(�H���*P��Ѕ�J� �!����\!�i#�o����m�s3"'�����i�d+���;r�}݂��|8j��[������AY�ٖ�����%�:R7��� R��2C$�
]$.U���r/�#؍=��5�4�����e�1�w��1dc5������Qg!�� 0hS�ȉe���S��`�4j,��b�~����A��U~�C�����7�Ym�?�ɝމ��wX��~	�q���M���W�˥�r[_���!�^��g|x��e2�)��D��z�Bx�gM�I�.�Y�I�CT�$h��i��L����7K�*���P��Z��чAC.;Sa����05^��ÿ����4�I]h���
��l1 �.��aE�9�a�x={�N���LP�ղ�b{���R��k���Dr��'����J���$�d#4��I~���z�j���X9����Ғ"m����Ψ��EMyC��yH_9"�Gѫ�(�װ)�㢪,�>'��pݾ�y�����Yѧ��9\S}��w�>v� .�g�����h��������' u8��2�H�\�4��y9����?=������a��s�u�@͒�U��93�ؗ���<�WA�b�`�7ӣ~���IZ�^�E;J����A�!0J�(���;o�[A~I�$��i>c����C
��A��Oh��R+K[\�:dǟn
X�V��&ʞf��FB��y�	݌˾�}������Dm�8�.���@�8K�i7qC�}���@��&_j���� ���?}�)I� ��\Rj
}�:Pm�e^�7ũ���bk���F�A�w���
��U�j�3梼@'����=!;���\�";�]���|��W�z�RF�lC0��`��� |��6We��
�������������o���!�Y��/��4ʹo*X��ܟ1M�n��k�:{��qC�ߜb��m,�8'�[|rxF����6�X2�מ��!�hh{u	TQ��q'��Nȇ6k�ĸ	
��q� s�?�9��$&��Y�YG���1(���4��/A��\6t6�۩�ݍ�"cfWӗE܄Zk!v�N6�� ��~j)�T�p�c��i��l�5Y�3�L�I[�j��x�9]�͆�*B������ ]/��ʓ�
��2>���Eߟ�;qcgU]rR:���34�v��������9I%L١��ݦO����[�����6��@
��9o���1��Kb��5TX-MTb�!�+9��@�j^�x������Ѫb	�N�Ȟ�U�h��	���w&��P�8⍉.�?о�J��B�Y��M*����X�`e��(�_8	����@87���4�BB��Ӱ�Jm�5r���X$]��ˁ�M�ǂ���G/Ly���@�3g�\���7I��Ҕ\>%͵F��� S�o�A-�v�E��g.�6
���T��K����Z���jM���)X�J���������ݔQ8�<p�$W_�|1�.M���JrM��Z���p��w�A�C�ػRT�
�@.B'�NyA���i���3��R1�#�\�a$���NvQ_eV��:Ac��&�Q���`Z�IӋ�&��s.yH�n�ͳ�8غ��	̊������	�4�.8�壮�;����ҔgͽpZ/ZI�Q���Y:q�V�PT�]"��#���.[��E&��k�{Лa ��\��G&���=�O�ȀQ�C�`��ƙ�u�j���{$���qZ������ڑ�mN���Nh<;,�³Hr=_4�fq��fL/K[�W��i.�6$V7<���on�fw���_��V�TS"Mc�����'�����\�j|�W��ii�R��\D&0���g04�K]W���� 6���,��H{�4�46IQ�ɞ;č^ɐxi}J��iЬ;��ǎT)�ц�`�w�⳰ё�暜7����$gc�Ao��_���k��b)�ȷ�6;8½~V�0+������
7�sXUt��tPvί8�M�2\_�ܳ�(��4�^��Ĺ��7?#3����ư�����"�A��_���0�>t��nK�E�b��ka ���Z�	3|3�G��w��dQ��}��6���w�_d�앢�2-G]5�jTjm�Ȟ[��B]�5;��&7�t���-��m�֛��6�0A�y�'1?�S�	�֪�2�� [��!B�	~����OX5Ǘ`�bV �?�1'	d�h!3���H�2�x^͸�02b��b�X�Rܱ�1�䵵��9�9&���tX��Á���ϟ}x�>T{dwP�������?_��S��� ���F��uO��}H����(G�5+�L�V�@$.�/��?��K~m���P�� �0wԯ�z�P�P̴y,h������Y;�4��������'
�l}O;~#x�s�A�P��iH�h۷:��k�ȴ��-���&)�R�I�B�B��1�I'���};/��J��M��� ���JYc�MS�H7������p�@Y��(���T�	�����e����s�Va� ��9".�fD�bЬ��+��C����0�77��ę|��7�.�
4M�ٿK�EIT-'j
�dN����;,:t�Y6U?����] =���zb�DXx�ºd1�c�/�͝߮��I�L��h%2��g��������:�Ȇ��4�$�����F���g�H�Ma-��TJ&����O!���eN���]��"K�'G6?��\]��MQ'�5w�j`���*F�7�T��ZtƑ�T�̦�YU��<_12��Z�mw{�]6ن�X���٫>*���������[��qQnr�2�M4��CH����?Q�!���0pN4�70���g�{��I��E �����7owa�Ü��e������A6��מ������t���:���wQ�a{c�c���VpP�@����[i���ks�d������^^*uRF��E�DHxϥ��i�<��c�W�жk������d�-�H�~_��4�`5:����D�C�HoB�qr����vn;*5̭��bM��*�?�y#�ҍ<e#��
��.$��4��{��/[�yco�=�k�d2��@T��$�?��ㅷSI6��$��;p.��a[�"�'g�B�*��VY�Ǝ��a6?�S��6Ty������;�bo��b�I|�X'OhS�Ϻ=�
��q���C���0l���@?~r!~Wu�/� f�ng�[��V�_%`�J�
T꘬P�Ԙ�5h��/�[��3�O��U����I�*A5�Y-�8���`�(���-�^����(�d��.��LG�L�'A��������ŏ����oc���*!�y�+�χ�0�]tf�1�v)
AqWmV�2Պ�{R\��z��l�c^X?����A�'Rq,��y ��j9a�M�l\:�"Qe�t�i�,����Y�S#ߺxkb}`��lm�����N}������1��5Ȍ��^V=�����y ��2#H�5*�6V��s6q*��Z��`#��b�)3��ӂO�����'�}�i�*��\���G�j��l�d�}�r�F7�����������
UJ�ū�\�(��!^8A��D~=�sC�a\w���< ���i����iN	]�g� �D� #
�i�*VF"��О��_�����ې%���{��j.= ��2���%�ҙȳ��g���H��H�Iʒ����!K�|�߳��J�N��V�'�æ���"_�E/p����=�JN0x�!�Q$ <�D#+C��c���Z���욡j�0$WEM~�dM�,�j��/@MUU��xo�R��������'���|��禰�ƶ����<�QJ5;"p:��}^eL$��2��63dQ�-��_	ԩ�$L�m���R����m�>����	� ��%{�K!��p%#L�m��6��-�"\R�H~�]�Ka��/T�`�6u3���� _��ȶIS����~��Mѡ/Ԝq�`z�s��|i�j��"��f�u|��y߱@�\!&*z�m��?��%:Y�y��@�r��&��f��W3�K
�X�����hE�m�k���+[�lQ�F�ISB�]B��F�����G��L����hw��(�Q
,h4r��v{�m`�M*�̚^��
[���ɜϗy�-�n��d4�v�#�����4�[t��C�2hN	��^;�W~�$,H�;�őI��{קf~C!y���`�����o��
�4��BD�|��C��t�7�d�(ݦ��\�˿̨K�@�o>4����>�ҳ!�bP��P�Jh�f�״@dw�fʶ< �ϕwb�,*&�>ʑ
T��6,�=ov
+����8�����?/W��������=��FV^���2�7+�����vx#͙��LR/����xUӧ��Qt�O�hT6�4�ov�0������
���K�%�<w���	�8����$O�Vx�M�`��>dzA< ��ԏ�O1)��V��@����ShE�^��)�3����p��/r�-��@�ʒ�Z੘|i�8�Q!�DA�(r�������$��Ur*�'�o���A~7��?)�h{"��<�f��s=Di�F}�H��>�j�?b�$�4�yHS�]���]����H;���i:gwY����C'��V�Y���%{	ҤZ�2�>�O��k��<9(R�;�	�a��.�m�h��eө�R\�-q�_�]r<�ª�AHϬ+Cs�M>��F}ЯC��k8�9�+%4�9�9B]c:�G3A��I��K��?>�:<���7lY�Mό���w����kҪ��$�~���{� �{��ʂarO���Vn]�ڠ2�	7��+���Z|��uz,|k�B��/*:��LrgdG����]B�2�N�b�yN����䘻D��W�V�"��v:����=�B�a���i $)	7��5~��G���h\��2�A�ߐF���1_�;'wk�	w�� ��:�	Wj��>��`j;��9]�Ro1cU] [������ү��́2z$���$�0[Q����H����s�h�zP3*��������l�T?�X�^.��Ȇz!^���>�9�ª ��É[�<��=���������CB�Hl����k�B�r+�he?՗��8z���{�ŇW���S�L;5y�m�w��PYfloCmA,�8��,h���m:Z�Jm���HP��Gq���V�gѐ�l�*�7�KT]�z��b�UX��,N�������7��P����;F.�r9��eہz�<I��X`��T_jLw�(�1�W�%������~�)V���̟\uq��̒"�s�G_۹��1٨��ץ����������XC��H����zmA���>�Q{-��Xd�a��Μ����B��;V��Szy����]k��H�^JZ�� ��v ���!8U�8��%��0���2�ɢ=?��@z3��r���F�����j��͞v5:>����~�	MW;pm���<�T�
��PwM��O����}�m�Y�Z�/M[_83���F�DWw��2DIU+���Ή�Ss���Kq�,�K'��
�C3Ե4]d���Xk�Q�C���CS��O�_ў��r�N��P���R�m|�2��Pԣ�v^���AD���rbY:�B�	zR8�f�4�ka�/Zg �ō��#�t��m�Km�����\���🱹������e��|�d��{n����S<�gx�b�v0�3I���IPM���%��r#U��@�����)���2O>%Y���}|���F���"vY�+�s˶S�e�kB�y�Zc�Q�׃����ģ�̫�wiW(���(��8�#:tjE��h��*:���>��g:�h���6��3-�7�62�$�o�J�*oe�>
�pc�z@!��oYM����G[8�(>�қ����V����^,A�U��!F�22�����:C"g>�/�yĕ�#ng��~~���T�d�&�Ae��s(u����=H����8�ZL�������6��9���?�F�����������s�Q�f��F4�u8����9�;�u$X���� +�o��Uϝҳ �#���2X��M�{k�K���EE/D�K�t5�G{�����x��K��D��c�a���i6z��:i]z���������G�	���%�堨X��1�V�ut��O��!\�U`�Ό3�r(�v���7�����^��T�:���D4Z+;揨�j�lU�ȭ��/x���L��8]&��춃�,���'Vk�.�̪�iD��Pr��#��E�e�N�(H��i<h�B�1�*�GX�tD��9y�tJ�Oy�����=��._��B��fe��RiIv�̔���l@�`�ͱ�S���G�B�ߧ�{�������}8�|�Z�2�#����&���T?"�Դ��� Q�΂|�����zK�M���P�z,ި����^����!�gK F��[�}���x��r�}�+kZ��92�E1*�7ª1��T��A�������Pl�G����L��o�g�v��6	A�?KؠY��@-�r�g�[��u)a����X�����$���_�G�^�'/1�t��������z5Rv�yaB��=PN�S��/P��?�E|��C+B�s�T�	�L��!V�!�+AJ������eM&٪=��s��p}�?�Y���R������Km���  tb�*}�"U@�V��VƘ������b��9��1�Á�&�?av�e~U�8:�R"�b�&YI�N�M�a��x�b�xD���z+�o�K,O.sn�.��ڤ1���ёN�~�ZhY��3Q�������/F��F	���Ty�����?ΎK����v�4�M��?��o�����U�#�&S��4�$wT�i$�.Պ��~�-~�����4��($���?T��Ȋ�3�ͧ�u�ac����ry&���%3HXM۩R���v|�����~:���	.��<Y\kﳋ*{�!ng8T}
��&�����O���&0��"RL�"[���N�R��C}k�񚇩T��fH��#�EHD�yK��Ȓ�|��g�@�k���A��zO�.�z,��A���G���K��;X_g�g����B��#�1���_�b-
��L�g:��u��UO�}B ����'����.��_�W�˽�b.�m�uq�A	��Yk(��+�w9��)��e�z�ât�Բ�"3�����bF-M��R��NE*[u. �	i�]����[~s-��eD'x��:g�o����F$e�qS���<o��>�h_n�X��8���N��Ϩi��J��<�4]wQ�R\�]�d�-g+�P;e�Q>Z�����|4��z�9�L.
�.9�m���W:K+�����$�5��7e<�+zl�ê���}R�*r��y��� \�c�.6�k'8Ys�O��Y�}
1�5�0zn17�Ħ��R���p*&l�����;w�_ђ�kE����fd��I����mVV���Nk<� (���3�5�JT�8U�Q:ϱǃ�0 ��y�d���qs�X�.�/	{2�4E�3�%�<?�
����G���G�z��/磆[������RD�9��"�	w��� ���������{U�%?f?��EM���_��� F
��H'���[��H�D�B|����S��J�L���&��F�3��4�oM���SR7=�������n�4����u��kרa�$��(�etZ#Ѯ0�����S��`���AM��F)/��ì�*EfK�l�j`���x��`���Na��^Q�菚��QͯW��s�
��y��a���uX\�?�����a`��>|&�D<���*|O*lŀ��&���q�+y%G�/0�0^y�N�+�8�99�G�~�� �����2�nM]�U@��V�ݏ���
�w�`ư8{�𱚑���9����~u8�ix+;���'���w�r��rB*��ȫ�����K"�y���=��XY�H��o��M��/W�E-7�i,�~���|�CȻ%�Ѵ~�R�ƃ-$[F*R�ZD�B���k5�a���_�1���D5���a_a�p�n����Kd�Wqb�W��K��&?���oMY�-3��+ܨϙ�	 �L���M��k��i*^tQ(�v��h��D��>l������bd�WET&���V�R���:��I���r\\v� ͮ0�8-��R���m��BEUS~��_HMŴ/f\i5����.a������K���m�B����@�������c��&yCZ�_i"��P��R3�H��� ���y��Ґ<��l���z��'�q��<���\������<�>RD�9[t�%�w0 K��u��Ƈ�OS���pT�AQ-��$�^h�Q�e1m4Ǯ98�u�������>��9�Q���yQ�;�g	��3���e&K`t|N�V��~"��Y#��-�D��U,�<Z����L0
j4Rc݋���RT��a��O��V�[�3)B�- Wm�f�����$L�f%8[�bF�-w���x?�����W�ݰ�R�^Ή�m�������b�%� 4��)O'�Vdj��`����wf���e�Co��,��=��2z]�N��nP����n�v�w�Ԟ���7�y�ͤ�zQ}�ɳ3V�0�fq�y�����y&�+j�2J�7��6����0�xi�&�����+�5x�&�vj�8=�P���I�ݽQ�VQ��Mڿh7(�)˯��!ϥ	dP�G��0$.-�U+�LD �[ۯ1���4��!ρ�j(��G=*V����sLE;_�+>@L�G3�|�X�FT���)Y�tw�ݚҲɪP�p�(bs�y���~T=T�X�p�<���2!,�{�~�Q��7���B��*YK1�»Z�﷖�C���'ɿ|x�6�'�䔦W�l�))���(��XxthQ��|������W78I����4lG,�*ِ����XW�V�'.r�����F�UX��+\����&��Y��ˇf��:�m���Ǉ�oo�E�^8o�ɧ�@[�����!�^�`l��dv��x�clݞ}��$N�1�΀��R��|�K����^.צ׋����b&��g H��e}�����ۦ���f�E��Kv:�1�4�M�l�m��[^>G`h^@�Z����j��T�12!��Xs�N4���O'㕎0%U���M�؈`^�5���E�mK��{jx�Aʉ�m;Ė�O�yɥsk�o4Г!�����(�"���9'᳠e&���E%��ļ�[f9)�z8=b���~�1���ݨn��*��JNV��.�;[��"�M}3/�n�M��-��L{iv�}���MEC��'J�Ih��:�H��V�7��)J�O��:�*�����GR���KՋ�� ���s�s S!KUˆʠi8,��>��E��P�.����=Z�Y�4��҈��ԅB+�uŗn�?�S��H����K�����@QԦ���8BI��>�=�����O��*98bK����-��77���d�	;�H���[�<Ϸ�#��!�%"��{VW���Vb������	�)u0D��)��&ھR���ٜ>�zʈ�C��X����ƑIc	n;\}�(lM��Wv�	�k59+v����q��J�t��G�ܘ����yF��f:��m����(�Q�Q��v�u�#��7�d�-؞�����׼j�����;���1\���u?
Zǈ H�x>��8�h�NaP7�U���W�(&L� �R�ƈ�9ҹ0lL�3I!��	D�{�tO$LRR���7�pX��l�vhV��K�s��v�w2�M�I���H1�opR8i85�8	ĭ��]O'���w��*d&�xĶfU��c�
�C�����<{��׋LW������S�'�$�S�@�E,�˗ S㺨y"֙(�фj�I�g�#�<�Q|c�6�nVPz��q�X>=%�7E��K�W�4Z�_݉~>��XzE;�	�L��ӧ�ٴT*^�Z��B�
B�}S��$6 �AtN�]���Q[�����X��F@i��4>R&�> [��ޥ���lgܓ���ֈ����U��%vl�@�7��I5�OK�r
St��Wq8���%h��5`�v�{II�|QĮ?�ֿ�3Ё���3����|pirIq+m1,h9s���*�i���ߎdp�%P�K+��s\��AA��)�$[�_O쥹�y[�A��Ӳ�n$��ٝ��eQ'�R�7���|�V4|�J (1�(5�`��S6���8�Fa��5��w[a��h��G�|=4f���f"\����r�3ǳfB�/���rUu�P�KWAs�-�X$�	�9�|�����>De�-�U��ָi��C�|�	���5S�^{K���h�|����o��R?Gp�m(Z-n���y�O���r���ؐ��C��=x�Bk���sY�y;�+H0ॷ݃��Rk�$�\dx�Ҋ�ȘE0�B��_�D!b�(��D��v;h���|��U$E;�B$oo��LV����k߯( 3
��T_Wݗ�R��P�|���շ�Μ�%5����v�x�Uje�̤j�o�בKz����m3�l�x+,�������_x
!�����"��6����;v�?����'7A?��$������>�82k�}�N����a-��4�E3�$�Z�r;|0�o�o���y7���xi�Ꝉ��7t����j{[�)_�ûp�vrm��݂���Z�&�h���h}���n��a��˨�l�R3x�Hu���_�@�w�q��"��d��5gJ>�b�ΐF��Q����yU�0���K�KVB	��5��_�.�߷��^�u���(�k�n�1Q$�W�b���?<.�o��ݗ��]���Gޅ	&�F��w�y�V���A� xt=�U+ilI�	<`:���9g�=SHAX^���������c�b8�)n�	�R�nĉp9&ۿ1�\w�sg�O���- TB�!��Zfg���[��*Z�bR�eI��	Y<jM`寏��6q��K�#�X\�?P�bL&쁚��,��o�+�C�x�j-��a�����{e��+è�k�*��0M�����@�cI��gyP�$�YW��S�������{͙��OH�6�fJ5�i������y|T�$��a�z���78�/��{Umڷ��V$��S,?;t���ȞtG]u�}O+�hp�7O�qf�Y�S+��Jr���_��Jˢ/����X�p�,!8�u7�mL�G�<�@13p7N�2ۧo��=�<��1G"!I��z���Pfu9��86km<x��%�������ܝY�n`25߸��"���.�H	J�?�2�W�a~s�$C�û'}���W��k�+X�HX.���X��+�8�H ,�NV�xS��	c%�����d�:J���	՝	' � �P�)R�6��6B�d�i;�FF�����8�˚a��$���E�A%�f�!,��\���a ;�8�t��8|�)���<�f4���<�o*��q
4w9�sm���U|z9�d��!���#
bE��L^���l�Moٹ�I�n�_!ŝ��6����+�/�(A>�֊�������1`�k�ICt���Y������Q�:��v* =k����^��;��cM״��S����Ӂ� 4�ˏ��N}�1�b��+��5"*�ȫv?�&g����g|�j�+)g�O���o[�z�re��Hc�б�舶����v���`�)ʐ�O�ڇhH��sb�g,�Wؽ^NE�
�T0Ů�bG'Oo�7�"�������
�+���÷p��G�e0��Dc幵�i���
�簏^��m˿��q�§��Ι]���d�|zϘ��f̧lO��9B��j��zlC�8q6.^RSI��u^{-kL�X7I�+W0%�1rw�pP�Ӂ0�ca3��Բ�1ŘZ²���h��հN.}V�]�\�1�/���t8�Nc�%4��hDU�Sc�\��˫�Iy�k����G��'�C<�%=2���K�]��R~T�1p9&z��L�YU�$?��� �� ���5����?k���-us�/#ɔzV|��Y��P���]S{G:�HV���Ć���*��c��.b Y��n����aZ��("�����
/G(LIg����vJq�"��r���=�N�B������|���lNkM�9涭��&�L"�4��uٔ���v����sxR�17�'��^��P�g�����yڎ�X���:wL�sG��J�Y��&MO�$H(`���4��P _*����{G4·LcS���X��0F8�-�<�%��fW��N���D�������U���v�0߯'Ey�kUN����e�t����`�8��k�a帐?":EA	�Ѩ����έ9��L���{�Έ�t#� m��|��~�c����,!���^������h�h�8�f]��Lg�uy|0Oe��R9{+��E?�%Š�*����k?#��k�Z�E8%P�������I��K�D@���m�&"	�j��o����C�jU�f^0CB�i�ȭ��mG���&B&_���:�B�]��~�[%�?k%_a�d��my�~�@��C��YkH���c��s�H]�6|�T�U�_8?;p�u�]���?��3OX����D���-�=zi����� �;�fx��ޏ]-�%�#?<{����o�({��T2T�CM��h�������CY11F�I�N�E�S^�?RB;�-l.qtP}�h׵�;���5T[U�A��>��C���O�L���U���LL���l0���0ʕ��l�*�p+�{���P~U�3�`��SϮ�������l*�?��ϥl	B�Y%�~~�2��Z�oߍ�
�,^��\�?�D��£2Tf��fC�d�<��q�������ŗ0yjw���[x�|)Y�{�n�U�	s.��/�5��s�3oٞ����Gr2E�#9�2������w��� �n�Cm�|t���i����)��5>n[�i�N�5���6��g�a�'j���.XO��~�;�z�Ӫ�����hq�O`����|���o�hoഏ�b�u�����������G���b��j�8�o��B� }@���X{��R\L��LL�z����A5�s�㟵Νf�7�[
l$ч���n] �{Ч�E6�m���>�M2x��ɞ��j8.\=�5DT!?�*\`W���c�S�+��u-;~>0����9�t�����"F.j�n�Xa�+�{�ȱ͠®�P��x�5�-&2��[�G�Ë�+�l
WU�=J�׈&?�F%S���%F<l�T�aU�lx�yM�F�g�z��
�Dd�$f���_�c-��Ux�-g�P>�ނV�$��8[���Ř�w`��y��Z�<W�q8�",���7���:��p':7� Q��d�
�^�΂��xXyK�l���`IF���y��uv8�x����L�#�ᐸ��Z�=jy#��$�h	�iPo��aY|D:��<���ؒі��6�2.ßA���F_�c(.�;��G!n����[o�9������K%�����/�
�u(��;�F��a@9��yV��靁����&Ox��T��?��5�x8 o'��s��b��i=��|r����V�����`Y_�
���@���-��e��iVc�Av���b{(��&���/�p鵫�"�9����v�|�T����>$��t��˲�A΃]���]�h>|��)���������@5����"E�*.uA���m��Ԅ�����C��x�Bl~���������)B�#�r���c2v�5A�:��vQ����ʕȺ��	P���&��ݪe*L�\���E#P�m��&{x��B�}�.iH���-M7��=ruX<�wVG������A�ӕEo�����������&��p���^���h�ى#p{=6�B�"�k(!/)��fPr�����˭��2S�E�tj��lbt��u�I;�|�b_6�Z���I��m�.?�W�*��ݙUa)��ČTה�FY7;����DȈ�-�7�s��ݍʣ":s��cxX�D:�,�������V}dUc_i�3����D��u+B�B4��3�T�!��>�!�Xq�T�=�	CWX���%���x%#��O@�!���hf�8ǯE�������ue�ϕ�J���U�آͿ�!��o�?�ٯ���l��@�r�H�_��8<��r��7����?o���� Iٛ!(V�* 3a���>�gJ'1��$ʱW��YT��\���aAI6��l�5�닕�' �p[N%D��G�2��y��z����ͬ���6C:�~Z�{F
H�x�.��z@~��^����
S.�d���fB���'-��'��u�)�)��և����U�Xr��3�]luD�~]"�~��1&�^d�L�F�r�ir��^p��b��R����A�/�hC������2�1��A�9Lv8M��Su�K����7ύ҂�W��_��i�cF��~�����<�2���e�'4F��,F����E�_>v�:��q��m�	�� �@lJK	�zCxJ>W�5y�kЦ#Nq'�k�zu4��w�O3���&n�<���.ڴ���@�c�E���@��N��}P��kcK���3�]`AK�byץti;�p��O���׬l���v��?)��J2N`�<l�����ؓ�)��D��p��[ p�s!����j=�'�
��H\����;/��H�l J�v;cl^�ҀMD\�>�l�я*鰵��
I�j{����y�.���9�	��T����N�k'#^*�2s��6���U�����~f�3���5ʸ|2��i	�;�>��������'��8G ��CŴ���U]���ŷԏY<�7�tә���魯^S�~W�f�ߩ�բenF
������ӳ����x�܎�!�Tj�2�^��k����ǭ�d7�P���H�1B۷���oSjhU���2O��VT�;���d��A�X����!�g�.'�;������b��2?���-���[{9և8�i���	�� ��"9�z��@)�yPR���?��i�-�ԇ�c�� ��7M�Egi�A��x�{2"<�>)5=��P�R��Ŀ��L��C�F�����Ty*>�7���v>��1
�y�ϵ��G�mH<�i�@\!�(@�U�G��� ۈ����Z� .G����M��%�Y!��+�a�zf��1��+�0�x���su�/��|Ti0GH�nS��׃�<���!t}�7�߸&x�rL�d�a��(ι�����0bV�"#�mt�=x/)&q���{L���m,o��8��%K�Q45�lUe-(�ο��9�]I�(�U�(��=#��J�����tU��B���>u!�u�NB���*�8K���VinO��8C���sm�{	A E�ES6���G���uG��A3n���� U�[p"
|~/a�S���B�U�{��݉}�Ty��⒇/�'���J�02-R���_l��#}�9"!�LԾ��C���I9ӷ$�_���|���d H�3���¶?l�X��X�'O�X�!d�e���5]պ;c|�����*����3�[ӄ;J��I�΋:!�d��Fcj�*\�쳛�p�4Fs��K3Q0�������/�n
^�G4G
�z�t/��Qf��{4�gJ��H-�EV�����|�����,~G�f�
�����n^�A�
�zm�S�Թ��6�������·����4��Y��N�p��W�߷w{���N^�9�>G�\\�yb�u����k��+H����]���W�d�w�VIk5DI�ARǓ�֌	��w$���>�W�ǾȅWOs��r~�F���;�*�]	!����|�]�rw}��^�H�`V1�;k�5)�{��?!���D9D	�k�F ��5�,7�_E�ZS)�?�e�z�A�? z߅6L��i�q�X���~���tI�ǋj-u�hnX�/-�j�c���"�2�v�]۔c"��]r5�j�iA���N��)�!W�$p�gS*P�g�z�+�cM���m��-�1Y�V��`��W�l�E���q��p�;x]4��Gച����t��H7c�Â���`1Z����|o3���M>�_��+L���T��[}�����V^�F.�N%��e%�K|r��r}�^� oa�[�g�W��`�z
��Fd��4�X��������������Q���K�m����j�Ad�9Tz���x��u��ԫ�T@-�^�hI�8`ℱUr��x@S�(I���*��mj<�k��祚�����	�e��ś��x�J��u��r��|�0؉C��ê�nʢ	����9!!� �g{Z��	b3,���bhE��q��حѦNwKύ>:2WƑsv�l�z�ٲZ{8
.Qϫ�?��_�Lɶ�r|�$��sJb�UR��z.���]&��%3_��&+�ۨ�_am6ߜ��͂�UA2j�����k�s��'�\M'qA}�h<���N��
�kd5,���S�҃E�3%ώ��6��ڵ�k ��,X�ȼ���y󳞃���R�x5�ek[}W���x�a�D�j��2�G����`�ѡ��[g8��U��U��R]b+<N�ǿ\��q�Eܣ�$Jd����ZG_���u�E�1��Ѵ2Ğ�' ���xb��.W��q͢ӿL��A���t�IPF�h�,\�]��?Ez�� 8�MzX������$�D��7!��[��`��~mf�c�5�A�1o�^�iVAk>]�2���+h
��ߖ��ܗH������)���"^��c�ב%��v1Sn��."A��-��$�ƞ$�DTjBN�A�rɢ$4�	̟ �(�{���D;���/I[����~���^������́]��B��@9���$���K�J���,���	u?����;�J	b9]��%_�/��_�1)�b�/�*w�v�vV���8�SBv�����Z_�d<�8��$I6�m�!���J{dļ
�
�XJ"�1P�{	h|�' c�u��?{� �#��	�;�����l���,7$t�V�������B��*�	w�=�k���s�֛�LЬe�&{���hE?���[�h_NK��<�9�#U�T}i�R����ߌ��$j�"D��$ ]�#>��N�r����Q�ߌ�;��HՆ�qļ�CP�~�`ڰ���p�?8��b�[b
՞%#n(�GK�Р�.� ����YA�t�3������;V��N�dx��<)W)Sh��tg�0j^rQlٙ_�Sпj�;) ��\��;�cY�[)'����!��#�z�j�&Dh�M-;����t�J�𩩧3s9�#�-���E��`�L��?D�n�h���q�3����EC�|��k��F�W�s�b��^?�o�����I�z�|ÃX��%����+����/�$�(��=$j����J�)֙'�%̊�������8�
P�2�Z6�=�@�(��#��`�z�]���h,�:U�[Q�_�z����}|��q�H�~f�`��{ �g�g�۪=�n�ٖ�0�;s]WCL�pCA'���)yB5��~NP`�E���A[��v���S �o=��{�I)�V�#�Z��ބ3�� �jjJ��|��1@�jΈօ�r�J��sv��qkWȷ�9���u�U���y�tap�p�vm�IX�gF�(��tYJh~9��A��T��Q�l�z/d:k���HsRq��jq��S�s��d@(�d��o�{�)z�ח=�*yR h�}���J9�M5�	��{�,^L���\v���>_�I��j2�&4v���S��xA��/��K֓Z�³��9��C����?���ă1n5B~�E�.���q����'�~e ԔC�Q[�-,�Z�B#w�1[�x�
Ȃ-tC�FG�Ju���U�cX-��K��<s\˒|�������j��B5�O����dh�4;LYJ�o�s����P�����S\�Q�e&-+ӳ4=������p#���p��bOM�h����|)�*�]ʳ�TF:�ӡ��a	˴���(�ع�!ָV3сh�l)-�Jʾ�t����e����O<7�[��Т%��Z枖fU������{���;���,"8��.x�=�"�B�KFDLY�%g�`O�YC�`�p'u/�T�sZ�~��A�b�m��D����	1q���:ԇH
�:���8�`$����V�N������C	_8Yj�@g�)p�J��q�a��2�@
,}p��(�+HFrz
��4���9��4Z'I.��~�i|�KkL$����3Y��OV�$��绠��u6"�D4�i]��LxQ�+�$�RyO���WE�k��c�p�-�%��u}�Le>�:�=�	sכ�Z��u�h����Wp�}ї��L�k�xQ���n�%�pP�w��٧��������{�(5��oM���xi��]�H�~&$_��$\�������ޱ�+�2��LR-9x��䃘r9��s�pUiFF����F({9̪���D'l�rų�>�i���;9fFLT}�O70���EȆ_�򉼪�%[㲏O��14:��;�d����T����Z1e��^���3�'�$a0dp�M��P)H��ّ�"�Hasz�����pQ��I������E6�4��� �
x{6u.ZD�+���^l���_CY�!�+*j�K!�=���`~�k̂�O.�Q�;���Y^x�fl�)�Ǐ-�E#�2�p+;=SE�fL�y�է#�j��@V��S�)��g��������R���%C��?olЋ�p��d8���9�,�]�4ۆDP��M]h�l���,�����+��w���wR�>�۹�b��3��n탈uG��3/3��$!
Y��3�����V��\c|$���"�@�l���L ����r��n�~)n�|�v`�t�;:��ބ?Q���<Y��
���t�%/YIA\�#�GLY���u�-�2����ԺVO;;�K��c��4n}�ׁ+QFO����6h"$�5� [��#���*�b�j]�\)���8���e�dmiGj���B� �h��.���v�P�W�S6ǽͺ��\�kÑ_'��"������;󦦗�PX�4���@-N�2�T),�1u̯!~��p!W����Zv�g�)��Ȥ�@�TYc���<���B�P�<(L��[~!
\��Ђ>KVz��O���Zk��E�%�ր�认���ā͵9� �k�}?���Z4ft�fe��0�]�������[J��h@�N��&|-�!�"����n�@�0��I�����������  �4�[�X������Wx�������B]�]�W����۽i]��]�����Ĥ�S`���� <zJ������� �u��}��}�<`qFR��;�,=uo`qK?Hc/4Ԋ��	����j��/p@۟��Uâͭ�vIjdIt��s�ur	X��vm���:����O�aG�o�KU��Jظ��<��x�$E�R[�!@c�ek������x��&���h�@��~t9<�D�����ǙP.Ƒ�/�]%������bw��>EH]�%%����N����X8o�'�~�z�ـ.�ď��i��Ms^��������m
Ѫq~ �[�=����RwaE���Xdi�ύ'R�p͜�/��4�L�%25b�a�.O4���Ѿ<!J;�����/1�_Y�awm��=){EV}u���e,ܥ#�N=�ׄ��'=T_��G�c�A��w��j��?@�(|F����|�B������M>�p���,������iS=�!6����ѯ�#��̡?ܫ��AH��Y�vLO5�"��n�*+HJ/�� 9�s"��h�������=ړ�l�����z�6�B���ҭ�ϒ����[H���ǋ�)���#"�j%5�6��a�Sy��C�PE\+S��c~[�A�Z�I��j2��%^�v�`ӝ%
�K��p�B%MUK�� q��@,Y��t�í�nKS��}����Y�T= Қ;����!1��~AL�8ˊ�I�еZ��?��k
/�:�bQ9W,t��敪����+g~F�c~T(\�hg\=x~�Qƍ�O�7�T����\�����sl���C�t8?Y|�(ڀ
��!�aԕw�ʾ�؍- W�$�脱�^&9w�'���VoV/$t�}����6��%�h[�|x�4a�����֓�:�i��;���v%.15�� ����la��ZGw�`�by?���������G�9_��[�b��[M�	�6����_�@&��@����Y-��Zeǩ�q�H#�S�E�����^8 �A_�#Vb��Ag= d���ސ@�5Ј�)�V�5n�v�|�D��N�S�����o�+V�I0Z�g�iQw�RV
��H�XK��L��[�+�-u�W�S<�2m��Q��6�Km�/���*��5Њk��]{g�K� p����!aբA��Ĩ�Oz32兣*Ӧ sOQ�,pL�,i�gD]99��~@d�l��l�V�5ą�YC-T]�������-W�7�H*߷��
=��Q���;sßWN�tʤ@T(�_�Rb9���a,`8�ރ'��_�ѵ+{a`�����ij��Bϫ��dn������I��3Mj���A��	٨�9n6��J���U ���x�����j���P'�m�w�-D*6�����)+���A���b'�n/�~�6�QrB�B"�6�jeSĢ�9��,��CF$7�yeS��,I��}3{�Fj1K�R� d	����S:�|�+�FN�{����CeϢR8��jB$�!^
�2�ͷ�d.�w4��CY��?o�>�h��H!�oU��� ����{4�9�@��mU�;e���]���^Z��]�h��_ ��]��ў�o5�ˍ�C8��Ӛ��9`7ߛ��� i<�4pC-j���T/|�Y����kFJ�[v���i�`���a�JX�EQ�w���z�߯�v�V� ^���ɊWB(�§���][��w^X��_9��2�`���Sa	��s}�w�#߷��M�\G�˹����'�6�zFGw�c#mm�*�=���ت~��}�#��C�v���w�E��}��U���}�����4���A�!��\L�T��;�.��KӉvԇ��H���][��y})�;$�_ٜ�N�X��qA��^���.9���x���/.�7M�tf�u��kav�WTѣmˬ-3�<y
��X�{ߔ%1Q�71J�Hk�s�	P0�`CG���4n�P�/���>��_ת@y��ȶ>��,�o�M��wذ悺�on� ��c��-�i���u�y�X^��1g)�x*;�{��𔺴g���bm��O���Ɠ�酳E (��s9J���Le�19����a��_����/$+���Xn
j�7�=x���W�H�&7�JKxVZ�0����~1&D~o�|����:��}|޴����R�\1�%&�?\��n����Z�ȫ�a�e��Љ�
=!t��p�Џ�є�R�I���2��'�~f�1�j�w,�co�!)9��p�{{�$ ��C7�0�7���ɚ7�>Eİ v�-�6�������q��a���z�-n*�,�����ve2�#��1&膊o����uˡ[\B�˺������@��H.����A�6��#�|�=��;���x�u�N�o�f�p��2u��\ߓp�ڝ��B�r������4��GE�����TQ��dO������@���'I�N;��\a�֤�_o�d�㧶rpX0V�m8zG��ܡ�,�F(�9��`"c%9OWL�@��G�%,���B���[�o����(�զ�8�TސW�ar�,�M��^�fh�΂�gɼ�|�ۘ�ăq��P~Ĝq��c�X35����ޗa�F򟌑cJ��.;e�/�Yɣ�d��ZDũ�,��O���V4mu �b���ﱄLz�Z3%�� �l�-,5��e��O�Sʆ�݉� �u��1�U��n��(^����3=[ �d�y��������&����������V�I�������a�Q�K�0�T�#,D���o�)_/��-Bȟ�w6�v��'�Jh��{�o�(����8Ī����tir��b��%�At�O�� �HQiu�ǥ�&�n�_���y�,�Ԏ� ���gҞ�BՉ|c���o�&��R�Vq������!ʱ�"pV�Jl�!�5[�1m�~K[�:27����@vk/���!��>�o��bR�a�[=����43
r	@{E��(�|�$���S�Ҕ�G��;��������aB�7鰈�_�
������{e�h�60ͮ��"XƅE���K�f�ʽc���˱��A4�(J}�H�&T
P��Xc��
x�T�=?yu:�	�%�*�ukӉ�M�(���z��QFFu������o�����Ϗl�.FłN��Hn6���0���A0k*��%(/�������e�r"�;#�K����ק�ia[2=����c���yZ�A����"��$�e�%��i�2Q3��~��U��.�T�n<٣�ޘ%\	���oF�����pX�9S� Us���C��b�|�r:�B�L�@߳�^���k/�ۇ�6�K�Z���������($J�Z�cH��L}�����.o��b�Z��_�Ȣ&=w��"H��.�^��HI�����8��n�5�.I&�����d�U6��v�C�gG��Ѥ3�t��<�G��:!/�zH�˘��}f��@�q��v扻'�GP��i�ς96x	8��ے�D࿜��3�-���8%KK�~0�>D�Y</�p��J���.֮G�f5G|�7��u����R�o������N8�c�_-rȢ�|cZR�i,dx7>M�U���?��su�xG*W�-Ae�K(ْrUs�:�>��B.���.d]V u%9v�����}��`hUk$���+{Yf�����{6N�ɇ<�l"�3��P8�1\�>9GKՓ"�|͑@�A4��l��$`�	y��o��H�γ*�Ȉ���횫ެ֫`E�	��_�3���м	�s��Jı��؈ALy�#Zq�����K�a�^:ޣ;����9yx��c.Uс@F��
�8����Y��q�aR'��!	�mtc��/��؜]�I1�畣k(}GM[|��#��.e6�^�]�!�:����pN���ނ�>�*�7=jB$n���c���3�G��IwFE�f���eŪ��ݺ�G͘��Wz�|��3�첏���� ��>x�!�_?��h
�� � ��܇8�mw�0 �c%�~+����:v��;{�Q͙}��3	E5��\�G��T�
X(�U�WXI�$T� ����$���dU��/e@�\���7�Dyk��HL����x��w�l��ܫ����r��O�v[T�1��2%-�UR}nm]em��)�o���w8İ�����f$�X���^�Yg�Z'�q���)n�-9Ɏ��١9��-���M_i���2x��dJf T59�3��/!����Qtx�x��?�?��P�B|���W�挱��s΁�qG>�څ|Qd�����`���Q	�7����VZ�q�WuuѢ��
�[`���#�?����E�vk�9в�@���F|[�-Ñz��I�� �`�����@�C�'!�S�)_����
}�!�4��d�>E����:e����l"�8;_���O�Lh �ͩ�Џ����p�K�3i6-���4;Ht��ȁw�w����pSg��m0UkZ+9+�MIּ�4&(4%����g�ё'�w(���N��r��H�:B�,���"��yvo�&����P�8��
��g�>e���sx���QR@g�}J2�ަQ}��8�$H��!������0�W~�y�\�6F�-�P5čr0����iB"�%��#��,�r�[4
s7p$B��.ʬ���Kڎ��|���0�w!��2Yw���:���Gl�N\=kQv�qئ�2��&�Z̰	�u���f}�,��!t����Lx'KJ|o��4�z���Mwߔ�U�[��N;-+
q�J���~ҒȂ� ���b���/���y�������bZ�q��.�'��\����8!�q�(bn�}������L��%tEu�l��?�����~F�Q�����hz]�������)Y��D.Bt��բ)ai!6�PR�)�*�|��FZ��G�S�A��x�sH�#�q�m!AT�kBB1(��1���7v8ʩ��-���� ��
c؃�(�>�4���^
��p(��CQ\p�|*�?V�;G���n�"���������xQ��i]��t�����%�P`P:Q�is~r�����%���PH1�S*��F�#�5�Aq�m��f�,�R7NZ�j��J�l}�u�9&��`���}�����C6��I[��Btac.FS*՛2�\RG��z(A�� J�撇.��fS��T���Ax���p�ȯ5X�r��f\.���	� ��E�R!��ӬܴHh�2� @�����o���$�ꭀą������	��X�k���(n�R4����~��Uo��z^f2���gĲ����X{�qxq�9�^���i��B��( ����#���5���*��w�W��)E��B�(���j���y0��R����'�e
!ǫE&U/8`tAv����S����A����S�@�Bׯѩ��D�(��W'�i������kp'�5�Z�z��^��0�ξ��s�2����Yk��c���
C��Tl�dֆϲ}\�t�&O�a�?��U�'�?E���R�#"��Rݍ5 �E�j���H�Lb^S#Q�e5�\��Ha������;�VI,k^6�+g��{>�O�g���Z�����d��NA�T��L,�����YB :�pY�j��Z��V��ȇ�_���C��]I�вxIF����",m�w��G���~a8���e��f.E>���1뎬�q\��"���Y�Fj�:J� c��{���=��D�-IA�@"K�����%���1��b��V�̒�c��!ƴW��qܰ���ֱӨ��0���T���fұ֊��P�ɝ)K�d��&��r�˼����8��)��޷�o���j�5��R�X���q�)ר���sN�:)2.�+��e���󮎢MA$A�"�s��a���\b�k�|J�9%%�&U���D�� �вa�]��|��=z�>?����9Q��c�n��l�]0�PS�@H�;���X����	���uW@��T6�#�á��+'
d(�up>�1�
�M�;��̹Q�}r�8b�;�-ʍ��f��-�^M�K���S�ƯJ�#x.
be�f�n�&�;60�_��7�G5`����l����ɬÙ��+�=��k�Nf7�O��?�7����@��y��'o��"��R/������:�>�O ��7��0�	w6#^�P��g�U��8 �$P��A����'�F,4��Ϊm�O�v�1ī
���}�E��Z$�y>>���e�]��-/�g��G?�A�K�h�,���s�޳���N6�ߊ�u��Fv���<�ŒꝹ7��i�94��*�����f;�q��W\�1p�$g݄���8%�D������W��+�nW~ vw4ͥ��;���8ݨ��[�(��He_C�7b�ᨸMƃMqО7z&)�}���$WK��)�q�pS5���&��AI(5�[
DW��Wn�9ox��jF$r�*/�ĺ�Av|�Vc���y�]��O`��b��1���$�.'� ��fz��N��ot�ty'�U��
�,���?��U�9�S��!Z��k�ͩ�#�?7���q0��r��ڥ/�i���t�_U�����؍/���~��Q[TB�����?��nj�-�?'��Q2�󠭃�OԒǓ��3�Y��)m�7d��St$�r����L��|6m)��Ξ/��X����R�&��3e�]{Mg��=m�i�%�&U�@[�Ȋ��>��>m����Y̥�"�(I�j�ȅ �t��+n_�"��%ǊeY�`��Ϥy$
���b�Oh���'�GدF���2/;2m֠�-�����H��Ob�F��s��"zQ���M
Tu�^��B]ς	�
q��d6��uP�9�{Z����kN����K��ЃHs��e���q�z�1;�UM\Ɯi��_J��ʕѹ���K$�NرFy�|����'���#K� �UG���Ƣ���)�� 7޴�d���ܲ����Ȝz���{�}�D�W\г����N�^���U�9�&x 2��r�gi�G�$0Nش?�C�l#~��r��E���_"���� KC��)#S���HVv.s�]�{c �B"�ݗ��ùˤ�u:k^�(쎗��Oh���؀�Z�xh��܊�z=R���|}����t}��f��S�L:O�%���Ackp��;�|"�T�ծ���$�CD���1sIh�{˱t�
I��f��ݫ��g�ٯ$��	��ڶY T�����`�Q��k�T�Yd
��%�۔���HjO�
K }l�����d|�
�U�w¸p�0�ˋ�'��rk ���.1�(�S�79�;���f��p��ۗ��+"x�V�j!�y*��Z�����u!TY",�S�켞�X;g[�
�0�.��Ke�Qo�Ō�(E(�����^�bu4�ٵ���O</�R�Ĭ#��I�A��*�-���p��=������Z6�_Iz�L��h"�}�ŵ}c@�G�֜��F���&-6���.����x^?<���C�ҼLܳ��~8�'v���n�,y��"�� `O�M�y!IIU_\�� "[����.4��k(	�q�Hܲ�ئ�u�������>�;1l�K�jXH��dU��ށh�s��v|0�^ڡc#�qPp��k 7��5gVf'�d2���y�)��_3E�\���0���`^��L�8d_H����*��t#�����x��wQ,�J*B��.	�����C]� �|Pb����s5�Ƚ��W%���ZYa[4��q��y4��	&��5�{�C+�V��X0�,�e�[M����<k��hby����"H�)��H������g�ld#�dLB��}��/!�
=�QɌ�Ƈ���<7���0�.�,N���3�v���H��h�HA9�k�������	t�@����5i�w-�`%��JJ;�n�5!Ҭ(_xBv�H�t6�^�G��@�mt�J�[>Kj���TSo�������+��n��HY���G�/���YS�2_��WI5(�M��ܲ4N��U��U�ȴf/���g�2H�A�XA��%f��HI��>H�Hy�sY��ő�6�XMA���惋�m�L��.��ʌ��	�:U���b����%�Z�$X����H_�A-��."����G��C��4a(�A���KO8�����]�Om���w��$� �׋ �Ӗ�
�f6;7-n�l�!B�������w5����X&��8L�&����M����A���}����P�|��v�t�2� )3�]��\d
Y��r�{���aq�	��Ύ߮�"��<��}��{Ӎ�)�Z�̘���@q	aծ2;����iy4/R�;�-i.�=�p�`��Y�}�G���8^���ԗ-�#�s����1#N����[`paҒ�V��	�QX^ӫ�6�M�gV��G�:�b�<Vn��n�`��</�\��Ma�y{��4��G�0��d�Yi���]84K��,(��qώ(_��Zc�I:�N)���'�xR�#MS|R�T��Ҟ�����2�Yy���TyV"���TQ>3�JEɡ�m�,_G'�Q6M��cK�����4`b�ø�(%��a��6!-�v���O���b�_M�:�8�x=���p���rL<��\Ԟ���dj����4@�9t?�ר��&�zof���u���X���&r���Gi)	2������#���i)�)M䍏b<Ղo��������.�Z��P��)('��x�%�!6�x���tg�8����=2N�Z�IR/��&3X�&��P���?��K�>|32�hFA���=L/�N�l�5�ܲv��v��B�Cu�p�Uwn�)�~�9_l?�2nD��&�c��k3T�������"l�b��T�
�6��lƉբ��ݑ�q�!�z�콑ʘ܌�\���������K�E
Ẃ jJZױ��J�ώ^kks[w��V�h������Y���~���7D7z��L���Ҫ�p����_</��P)_|0V4�p"���z@4"U��[��{���kÂ���Rp�]q̶���"\l�JMp��ǐ�7~<�!3+��jހ��@����L~<��}���48�g���M�C����t��[-7]n��Πzp��NSX/�|�����l����V����x�?�nY��`�V7u����xG����P��nح�X������A6�#��
n���ף�a3�tڋ�w�o�GKv5���TmmE�&P���t�Z19���R�g4�A�qɖY/�*n�K��m���\tApEl�st�٪��K�΁�)��S�5�U�d9%9�����j�0 ��WQ]su+OJ�`�k�>D�L\dp�z1�����>���a�mj�JL��ad-	Ԍ��$�X���!�Oy�[�k�����>�Z����ėo���f'ɑ��ܬ���TܮBL��w�L��bY�>�ʇ)���[Bk��6[8��*.r�l���Z���1+:@��;�޿������F�x�
v�d��N��p���h8Y�Ʊ6CF�;n��������R��}�C|~Xf�C�ʺ�K���ב#_{1EZwA��Z7�n��A�׶'d�a��E�c���%�s�R��
LE�%�F�yo{#	�߀�/���[MٿlB��ILk�o�/7����;f�X���Z)}hq�Qv;o��_��j���'d6b`��Nc8�����֌J�<�M¨��n/�@�|��څ�B��b�=-�, ��
Lcd�G�\U�o(��b���K�=pH�G��B����"x�����Y����Y�P��[��)�*���Gi
��O��-��z�-r^�)Y��0��{�t;�NC����JA����c�P��q��ƅ��tՂ�$��8�������S��^""��V��ߨj �:Q<�*�L6�ԃ;��6蠪z�bf`�X���T��]Q��4�ܦ�xL���@τ�8���s	`'�YA3}�)�H��Y��Yk�����J��@�(��.I���D�� Q��:ߵ��$���h��CU_��K8�w�Ǹ�B�$ɕ�2�(y!�&*#��w/J%}a�/e3���4L�����㬦b�59��cf�Ov�����&1t�B8&��X��>���������2z<1�8�qo����U�d�ndه�T޺��.���&L51{�1�G�-4�H�%�r�Iy괿��g��ඉ5�5�(x�{4Ÿ�����>��C�C�%am��ӊ0<��#�d�?.F�9�kw��[��ȪI�������LP �^{�������[l
��k�u ��AbF
��8%+� }�?�c\��������Fg����,Z����-,Ah�t��p f<�}�)��ӾO<yׇI�(�ci���Bz�q� 0��:����8"C���0�P��[�3��'*ꚓk;�Z<8�wǨ�U�1,�hj��e��\{ƿ�lo��m��A�]�Z���U�C�T�vL��y�_3ud��F�@�����'u9.�ѡFJ���(���u�2�%��Z�EG��&p0��7O-xD�[#�f�W���,]�T[@��`�-L��-w��3���R�wO�?�2��	�
F����K�D��5\��BN3�7�����h*�ux��X��	�\o[�~`o�et���bZR��d]�u@�����!��;��`��N�&���gTM����X�c�v���R?�ֲ�#�g�8�Z@Ѵk���x��(��\6�+�����}�	[�*��]��_�ԭ�C�ڐk&�j�n%�c/X�� 	�Y��D� �[m�z}���N�FlH�el����/����~-vi�]|VSN
~�y��$��F�qڪ���}��e}�҃��z�E��p(4���ojlM<ys��n�{�d�R�<j]����t���@�@����P�Q�&��75뎎��u�@=�r�u.0�//[@ii2�!���hh� n�+h���1���#�4y�?��)S����1���zS��"�mi��[�ı����A2��ī�5ΟF��_���=:��n�^�Jj�#;�x�C�9�SA;���L2�Ó��H��"9j-Jv��t�a�k���Y_�\}�6?`��4	�?U=�/#��;�4Y�����4ݷ^�B�`��3om�x�������y�֋sG���5����J�gN�;&�G/ԛ'f�LS�| %(����bwFO�Y"�[Z�};����u��aNX�½��6"2"w��Z�GX66��m�tM;�ƁU�W,�f�))�#�;߾	��8h}��N�fvD$B�U�8�/��%<I鈰K�o�o1S�/`�w��T������9.�Lywi]��5J�/"��ZH�/ŗRR1/�ݑO8q�;V�2��OeXq���tU+�<f�����9.k&��������6�K��>�^��'Nw]���if�)��jz>T��a���H���\�[ގ#�d=�xO;]<��TC�H�%*�Z��[�Z��/� �?���C�!�����^y���H�ϽHѥp��ZM�c� ��L�dt��v�.��!���Ҿn�(�Hh�Pc�Ҥݑ�n��ݝ�d#�"O��B*��B����8+����t�?�6�"�G���-H��]�O����d�e�J��kl�G���3ǁ+���K����o����W��qZ�>��0sC�]����0Ec�O>�h��|�A�c�L_=����!�4�F�\��OǴ_�3�=� �&ƤDZ�r\\.�����h��芜�Eh���o����e�b�9|�7���yZ���g�e��B�\�����OӒ���
-}Ds�T�*�濲�+���ƪ���� ��L7@=�.�s��M���:jYA.�gW�q�Y��Td�q]��ئMC�D�����M4�M\hg<)�!��:=�}���.��q���l���j����p�GRn��6�V@�m§�}���'����ǀ(<9���{�W���������V�Ҁ�Q�m�ΰ.���g<�?�.��|�tQ?�+��}
�JbUڎ%�1�9�{Eq�_�=W]��$K�s�	�;�&h���=�7�9(�Oĉp�,XP���n� ~A��������A#���D�'�A^�ҿ����*�#随0��ieR4/���I��Lhrn�?8�.���\�R?���D�~�lQ:��C�s�,i&P�&4'�fʋs�C�\�f� ��]�w�"�;K�����p�N��z
���_�>pʫz52˽6����W��R/��^I�I�����5�����NVႸβ���}.���_��"^�>0�B���S�%qS:�}-�<�\%���f^l�y���u?ף��{ݚ�+D�����{BC�lУP��O����/�a����q-�*J��^��i�L��j�X���7�zE�R��8�iTS����������	�nĤ^1����d���V�Z�u���
�`��~�;�K�F�?�E��~y��N&�J웿-ǜ0;T�FޘHQZun�5�/�^֋OQ��ޱ"9b�GaDy�o N��D7��+d!��y\���X�" &� �,�>BX�j&r�>��gP��8��ĎŔ�C�b4d�VF��-��i��p�Xx	|qc?\�*wG^{_�2[i�.l�$x���*V�=m[���F���Vd��B#�%�����t�������ߏ�v4�$�G{�+�<�ݐt%�-�2�.|�O�kޅ�LӀPm��#��g��.�� �����A���/�,đ�KV{��]�f>�Q2�'Zy�����8��l?��XM���\?u�J���-5F!���Ҙ�y��A	�K*ܚ���go���J����٫������w]���c4c�!���c���-ߣ�����RH��ٹ\m�l�zoΐc��ܠEU���dJ�H�
�&n���:�������wa�u�"aa3k{�ⷢ2�{�dm�9/a�ڇHÆ�z�(^�� $�Vv;�Oz�O��yM�>�,:'H�(�,�B�}�=��!��Ȕ���>LK�x��iz��? *Ýy��y^)F�^0��:e� y�ȴ��S���ؠ���Qo���� =���WHB���6%)׮mJ�/&}o�I���Y����"I�,bf{��A}mȅ?!����"�q���W��Y{����a�?�+έ�3�l�ȯ��� �����U��s�W�sr#��v�P�ɟ\ǰ;2��q]����e�X��
"c�,�K��1�*��+AA�+f�W�B԰�����6+z��H��X�e�4�Ꮃ�S���R�� �K��?�R9eiQu�Jx��|��&�"J ���Y��KP�Yq��4Ժ�/�
(� >8�a.!��e�?I���䰫nq��s���p��a�5\�?�pǠ��o����P���s��z�6�MH�2�{�������8�}s�a�G&�p��'�|+�2����c=<��%�u �AD�{�)q!�_ǚ�ZP*RjE�����^+a�t��d%H>�2�����7_8v���h���z:��x��ߒ�=:7����_	�����7�ZnS��7��@oF	1 �<U��$�6N*���l�_zC��ͭ��C���w����8���K��)u�0�}�v�r~��i%P�{�����P����ٔ�����X�g��Zΰ��߮��H)�H����������S;T�\�0�3GP��-bՌ�򀫂�>�����o����W��r<�L��C����;����N��4�?��3�MIm��F�M�OZ���߭��5��U�
㎶�~IT�A� D0��������;=�,ā̕�^�QXO# 
�[����)�x�^�0�V�	MVv*���%���.G�'�,5>���� �?��btTS' ��k-9f�	z������zח���=ۊ#'&c��о����acļ-<��BD��O��n#��ds�e��N�s�A|?s�Tr�#��0��>��`�P�(�~k(uҬ�agj�� 2|B3������f�����P0�M'\�4��c�J۸�j���<�G�H��0����I�t:C�d��~�R7���uG�H.-M���g���8��}�P2NSp�ߗH#Ģ+D9�2����-�@{z��.c}�[:Ҳ{n�Q'%�PJ%k�����^�	�\�?v��z��ۏ&���n�ski2�7J^Y|,�a�ͫ J�C?�QTw�	]��m֎�
 ь��
�νQ��r?å&�
#��*��\�	v��h�����Nr���b0k���3�i�!.ǃo9��_1�1�d5�=�e�$�S�	8���͚z�=�b,��qcЁ�)���Hef^i����R"����g�@Va9��`A����1���˱������,Z��]Ol!t��yg=lFu��M3�(�mܧ����ä�6��x=%E����<��_�ιW:?�����.��K���W�2�ܥH�Ϲ3�
i%�6ۛU��^�[�~}�Qn.J�PM|�����h,�?�9 9Z�j`a��k/Z��O�ϯ�Z�皆��	��`�|�;�ӓ��L�N�� �*h�$�3,�;���Y��N� 9vT��נ�N�k"�GJD��^�%�E�qW��DD>�ѻ�n�#�'��ƆE���.�Kd������3C��m���Pt�v�՚& K��= ��Oe*o�A����Cac$S�v�����a�r�x���Ӣp�l�b��{K�NS6���;eJ��嘔��+f�wbl�1.3�Yn�.���)C�X���I��K�Ә=���>S80�����zIˇ�1Vg�;6��kb _A�ѹ��ep@{r�jk���!�[�ͽ��wxVX&�SV�Qu9�8h�^������?&4TV`J������(�G��DŲ�ً%na/d~Ԭ����6�#�A���`���L�|z;l)�^Ob?f���7����V�q[�9��lVyUf3d|�J���u�yc$��M�_�:���I��%j�M`�#�j;>�$�%��ƶ��n�do
�;dY��')����9-oyx���.N*aF����r��5��]4?n"���!��J��9υ
�@a��s6C��hސ��RXC���O��8_�,�Y4׎�6)f觙�\�$�Bpt����U`�u	2]gറ��	{��^b%�,�L���{ WUѡ��@�ڄP�2VT�U�.�^����5�Gj���X.�K��l�s�A�T�E���v�OXo{��۾8��E~�}���LrH3x?#�F�_fp3�;��4h�k��A�-�v"h4/�J��&;ݘ^��M����
��o����&.v�<,Y�Ud�ڤҿ�D�˒�7fw�Є5W�j�&|٢�e�n���$��7����6��?�)\�I���v U@�)<AwXrr�Cl���7��餒P�N(��eWGF(�;��Ÿ�>������O���+��u��6;��@��V�(�{s��Ԛ�+iZߒ�E2�,���E�Ì����*�a=�H5�TcI� �xw�!R��8�18(�hn����Hc$�u��E��%��f�H}`Z�����7�� ~�R�s��4�F��ɬI�	a{NEl;�S����E�9��@ϊuJ>	Zz�$�u|o(ށ[,�>(d��`�<��5��u���!����s_��&�vx�*f��ȕ��I�Jg⎋��IҤ�K��}[
�jX��1�5AK��=�Zv�(E.w)ۉ�k���n=KN�u�˨I/p���o���|u�q#�cn?SO@<!y5�P�J0�=(���ŉ�x^��M�k�<��W!x��?Rg���k��1���ṿSx�;_
β�sAc��X|�8�>�t�۟]q2�`��h�ۭ���`�a���&�Lb��L�����墹F]�hXj���:�`�b�em&��%Ki�P9��ҀJ��-F2���Qg��[@�9�@��������$`�,�<�[(Λ#皖I(�����~*�K�w�~-�d��-�V>7� ��Y����K����$\V^_��]���%����.] ǜ�)��40� L4�1�[H��+�9�$�r��5�����Ø��-�p�!�3�Q��9��+74���=�lJ��a��ǭd���[��B���4�q�k���U�z�[v���a=��6�"k���U�k�V�-�%)-�w��Z�|($��E8,���n�2(��8�T�DS@�3��k��W��O�i*׎��`d���/@Y�[�Ty����MX#ͼ#RB�s��l�}j��ōV������m�\�=^Aj�|�B�tO�>xc��H����0�U{k7����No����iqvT�~���`ƇH���\��3���<C:3�L'���<�Ȫ0����X��{gvF=��#�Or�!��t��
]p�J1UL�����{�eᨭB<���t�d��O"Ha"�{��-�t�I�}φ�E`:�I�R�R'u��R%�؊t�.?:j�ϲ��E�+YM+|����	�X��,abW/�^3)�]�B���3/�tgMAML8��39��'���i�_92I���[J���[/qs��<:~��A��AL�	�:����l����S�(܉�[3��ȿ�=Bc��Q�tu��o>���_��9��;���//�-֏4��?�Iw��D���WPI�#�Ec�t�~Z@w�a�͞V��p"g.6
��쪼O�C�y�	I g�Cu�$F?�Hx�7 �1RP�Y��.滢�Ӂ��_\��@��^M;��;]qb4�F��S�����I��L�~&��j��n��_1�_�M|lI�碛Y��A���6����yn��n��5���E�"�t@>o���b�w�s���9��[�3���g|��dM����+�1)���:Ŭ��R�n<GC�Y����4���Ջ�!��ZN���M|��
6.��2=bه����K����	�PD�冕.��j��B�6N�d�>$͈g�����ߊ���lјT�]p����{Ϩ͎��Y��,��$қ5�����a� �&���sn](��xM�m^�6�qvK�#�*x��w}�@B'���r�q�����~"r1��H�{�5`Br|���-<<�Ǎ�	��L�r��] �s��s��?�u�L�d�}�������ǌ!�� A�̺���hE#�3�**�3�ֻU�S����-�����;���\�8$g|��0�B��v$��F(�D�GሤK�G�+���y��
Ǉ�^�|�����O�):� .��c���>@�����q9<H�����z��L�����v.���C'���[2���ĒR:~?�ƪ�V(�ZMmD��t~k���U8øoL?��v�+�P�,D9�t�\G {��g�SJ��x�QS/�"L�T=CT@|���F�~�c����F ˉMs �cE����E�ܞ��F�jd�v#���*�"jg+Z��k�� k	�G��8��u�a����U5hy�_���?�ס��	_������A|�c�#�n���fga�X2㼧��l����Y�����?��hL&�����/��~J�<���a������Q���#e��ψ�O��$KQ2�
�=q�aå������x�~�by�_��1���¯,.��ȝ,�%�.�����|����Gl�B��o�
����M�=�MU�Q=�L�Ȼt�q�}i2Ѻ41@��=}Θ��RF����@2�����_Fo���0Ȫ-F�m�'����b^�e��qR�`��n5a��Q?�ޛ��b�}ˁ\M���yz��~�#(#��t������ˁf?��+1���d��x$z����K�^6��u����sCK����p��'�Tܮ� w]r����?Y� ��}%��G���ߙ�J?Z�$
�a^�b���ҦZ��i͙pG����kͣ�K^�h֭��
pT��1=�5-���o���t�=��*�=��/?��"7뼳���"aa����.M7Α��bK�B��Ix�`���0	�l����7�:���KAE����;�Ď�n�ǹ�P��90B�����Mb�~2�<�ɛ�f�*O�Y'A�ܫ�L:��]7f�8�O3W�t?L�ܵ���]����mO��9�X�+ZE�B���P�	i��>�Rl,�~%�U(˖e��{h���B@��{�m*�SD/�&�3.�Ei>#(�Y��	&�=���^7��ؾ�۞�1�-F��S���gXt��`"�?��
�n7��h��n����R�3��k+lۈ����R�f�,��ڋ�)�e�CA5�`�^۳&�Y�K���F\3N��/'&��B%��(���8jFJ!���L H߰���d�F%��d�>�;��\Ѳ�>E�%w-RJ>s���R�ߛ�y��!j�N���ќ�B�H\��m���k<V��5�hBu���5&�����݇����T=�
��Wdq���I��>�sO_���ܬЃS�W�b�<��]%?t�kM�e�� %w�-��O�du�,�~WZ#_�j�����i�.ӝ�H?坦{��Z`�#$�(�x56ZPʉ�+��'���Eu���H��h0S�D��dZ+f"d��AY+<�N����tm�&��'��vn�_��%zi���]�#�<ߩ^s��1�:�$h3:�m�ѶG�2+�9�S�z+�X�&���
�"���k�H2��g�̡rı�ѢLKK]} �븆��K�,����`V;�S�o��v�u$�J�<U����4Q�0�rב0�Z�)%ڪ3�,	����}W���*��LN ��b�(g���]�H�T+�Fd��UO�L9ɦ�Ȕ4�wU�$�Sf]J|�@�W���to�?���D,4���L}��|�!���\�b��[�CM�	��K[��Z��{v����S�!qhj����fo��o�����b�� ��x��e_��B!i�VB��s�MX{.����t�^���t?���LTN��5@�gW�ʶk{�`��l��c�)�?n���r>�&�հ3�J݃`M�~��r�[�hlwVŠ64�����d���QG�7��.�K�R��-g+�7�S��'� ���ρ�w���M��ܡ�b��ʽ�L�i^7sw�0�ܴ�
]�S��&
SE7MO���lH��"��GE,��Q?�ת}���HS�NE��D��PxL��{D����R�Փs��u{i�K)/�H$x��+p7<�.��E+���#����Un4}��\S���4u�y7z���JO7�x]�jl�iЙo���E�gz�K�U��@RɇFSNT-�������%��L����R_u�1�5���\|dY_0?�q��b�݅�|P
wN9�2k��m�Z�bKc�n�p���˫����_�!���E�)x[::�,��'�VXb'����t��>����\>���we�C�M;���ɀ���,R��kׄ��BSP ��Nt��{�	�������TgSIt����h�D �@-����k�3��g�J6=`/����=)�X{߽w�h�7uQ��տ� �����Ա9%��O�ѽ@!6!nS�	=�����Z�YU
X�/5<
]mr_���3���M�rw.�:��������%u�v�Z�m�6A��/$82풶4��+�1yŎU�}����P��p���Ʊ����5:�1�T�ݽ��[�2�=�u-�L��&�z ; �6�A�&έ�&h4=T����o�_��o�N��Q��Z�`?Ii�@\��/��Dʝ^����1(��N`�F�F��];�������H���k�z$�F��dTd���۷I	s�ϣ?�50���Y��,.ȉm<FR�k#G��D �:eXs����E�CVJ�Ƿ(w���-����>�:@���f$�Q�	E�}Y��&kU&˸7Zsz�?{���b7��h�J�P�1��1�2�?$3����٭Al�����N7� o��i�� �W���6q?obv����nV`dd�.G�i��J$�y�sunG���,YkC�����~�@L�d~�q�h.%)�F��B���EiD,eq��� L���#�#�/�pq��1�p �Qf�R���� ����A+��{d�vsga5��D������h]�#!�E��#Ȧ;G�S��|�=�C	[������4�/`#%��)��j88`-,���?����^̈�%��K>c�d�$�%/�{:�)�QA4��4�yP�h9�VX�:�8*#����	�i"T��T����:�z�1�v��7ܣ�1c�d��	y�vE��0�9��?D[U�A����\�o�?���S�E���ƶA�@�3����Ǫ�|,39�,/��kf�KzW
H<5Ô�z��xT/RgS"d�E��w��EJG:Jݭ�D���b=꨸�����ẉܹò#�2���Y���o�=�p��h���HzZ�<������5�d�u�- �LPJX4�\i�co@T�ފ�� �q��zS߮�������A.�.�%/7*�$��nUT�6�Wai�u`�:3W�m���*�+< �m^2���cB7��Yrs�z���"��ޅ��w�J�<J�A u�[#�5�7���J�f�'qgRb�:���#r�y7:�}�?>dCR�N���[��)��w��r&��ď�|���_׀r^6\�֪9З���I��68��my�U� ���#U�P��=?±���[�P�8؊�� �c�ˠp��/���:_�W�Ѓ�]8�y�$�&�)
m)&zHO[��'��b��������^�:�@����(rP��� N���ulp�|������m�	�`���I�>�ÀI��WL���W�Q�E�Q���)	��g���D�[T����.��Q���3T_�h��;4�- l�l����>,�Y'�B�x�0i�-�]� )M��Q�W<RJ�.R��r�)RQ�(�p��퉥�H�\�QR�7O-Z,�IZ�{�H?o��q��>��8uw��?3�41k\����?Μ����W��}V&���ُ�8a,C�-����.~�O�R܊�c�4m�;*��Z�F�t��
ũe���f��z#���S�v�=3���ӤΌ0e��I��s��^��L�;Mш��q��/t�bQoeD�{��u�R n�}���g|'֌>���֯C�X��fW�n�;N�f�K���yk����T�=g�熛���%a94�S��o�R�i�hsf���\XsX
~�q���Ï��x}F�,�N�{$دϵ߂|�������4�o�H�h��焎����VXZx?t8���[��Tۜ$�`D��	5L��g5��PK(�[��(D���)$ߌ"�q�s����:���#n$S�T���tF����kq>h��v!�N^�]z�B�F�$4�3�i��&.�>���UC C�(q\���������5eMm��������q���Σ3��qY* ���,]	��J��%��s�b��{$Wd�}��e�3��atT�n�b-��u��R�-D�����	�'��Qr&X�b_��a^�eH���+��*�s9�i�	��a�����^���d^�)pL�"�� #=� �$a$�8#M8,�'�綳�Y	�yQ%�ym	��KF��6������mqe����3�S���oq|c(cp�@�/�q�"h���ƍf�%a [��'!���'fQ�Ш���~���]O-�Z����_b���f�{����[E�9h��.���*O��l�4�f^�V�y"����JX�V�ʌ��l�M���χ�!y /s� W�4�E�W;v7��'�����O@"Z����;�'�z�P�dM@v������l��RD�������;�[�0����:�R���uk��#��T�k�@P��{W�P,�L:����\g^�(B���z� �}}���5?wL�q���/�M,N
+_��|������H.!5����D��nc\$q+��g��+�������Ĵ�G��JH���1:��f��Y_햋�otr,�P�:�oK�y�0���*hF���z�yœ��ȷ�;B�4��������I���v�I�
�G8@�q8.�Gϳ�����Cw
�C57i8����(�yc����9'u�c� Um�DCs�k[��=�I!���0�E��(��1�R��9�,�޸"�^Ob/�b���|�n��ť�N�s���ů�3��$H#|`�������N�ύ!6�`�Д�OPb�Ƙ&�1Xn��p�R˯sݴ�gr%��҄I�.'��N��2H�&��f��8x���`Os���D|;1y�h�_��r;VR��x�@��؍V��en�e���:�@�s����O
��6��0
�%��
mif�m���@x�l�j��V�az9�VX� ��6m5�c<����G#�߹�7��#5
��=p�fj��ʋ��߯��T�-�S�rQN|�	ȶ.�z��Zv�8�J-|��ղp�V��89�f������~����Z{��;ˉ~7��`��ޫ�����_-H��	{�o�{*����s����4X�
M#-P0L_���*y��ϋ����6�[�q�9�=�+cCU?d+&�D��� .y�GE��!� P��\��_�;�$׍;���Q�TU�����ճQ�������:%#+�ϐ��$���T�=���4A��v�$��͸�ޗ���N.6���~��L#�ƚ�F��ꈾ������Q�B�,�a8�D�$��"r�Bb�o�Yy>���A*�
����&�Kup�w��\^�@�	��^d�"N�J���L���`#�?������0@K��K�R���)3M�G� �Bl8��l"���.�뢨���ݸ�g}�`��sń��`r�w���(�ӯ������R�v%ὦ_{�%�S�з��Ȳ��05F?�ήF�yq������x�t9�d�3���y6��O��I��X�Ɣ>�[�����b�JB=��1ƶ��l����\Ե\�P�7u0V���珚K�Ű�1]Np�=xyG��+w��X�ۉ\j�V��U��T�v�eč���M�0�`:���e���k�$��2���A�i_މ�"���;S���<���CP��(�S�����Oϝ�p�AUbOn*���V�V��|�#I�����GpG�#@���`��Do^�Y�� ���ۙ�x�:��� NN`���%�/g4�FcU�pN��ݡ����S�"�7��Q��w.���q�ɹF
�d��*T�W��3�0��Yv��7�?g�m׈0纭�N1AYs�Qj��X"O>I.3�H�N`�̗T��v�LC �V��/�Ml�f�18/+Z�⮓�BE��K�ͅ��?6�~��V�C>gB-���x/K����=x��y�2����S��1�#�3ϸ��{�TW���,�:7����0G��8���T2�4Ĵ{èA������iY�o�Ko��3R9���V�������2��F=���5i�9�8݀F��־Y���d��~]��0��K�.��
��+��$��<���uf���o�ŗ�Y���1r�uY����[-���b@.���$	)�k�D����'���v=�=DZGW$u#d��T&ɍ�dF�!**��Q#���7&��D	��x�$b������{��(�H%���a���bKUp��х����{9n���Ճi���V����=l�Uj����1��U��b����EӾc�Υp�UϏq�G���=��WvI�Mj?]�����{��+�v��MepG��vsV՗��dҦ�3�M��������ȅ����z���-�&�l\$��m�!�����������,qҬ�ph�u�ѤS��!����+�4�]�I'���K�HЩ��0}��`��\�o�fk���R�R3"�4�*��T������UNWyT�%��Bph�!�gB�d&���I��5�����V�#F�O-J�7>��m[:���y����>w3<��f[���T�,���_͚�W���^q�ҍ�h��]H���:PV&El�m�{Kl	}�膳Y%�zE�ߕ1K_7V�+�oֵ�I(�������&UC�(��X��V ��~�붕���Q�οa�3Z�G��(�o�Tk*LFe~�GX�GK�l�1��0�W\$/q)�D�^���p�4+�I���+&m�I�hޙ4�g�@�FR*��JU�9@%�m��x+,h�� EVe�i���z�5����,��i�����^ďp"�o����@����������떁,�D��O���K�	�!a�0=���h����z^뷗P�Q&$��Y&[͐�y�B}-�OH���?�)��Ϟ[�l���#>��a�{������5}���Q�nI�=��	����!���X����?(�|�g�^��V%��c�Ԕ=�+'?�_�z���~���$�\6it�������KTu4ʃ��7�>���C�(F1Yá'���w��Ω��;n�tS̄`�AݼB@a�g���=�TQ����5��:M�i�K���s��װܬڔ�܌��I��a���8�B��H��ۓLƓ�˾e�9��kߵ�:]I�j��'��UDԻXfS���Nu�:U�t��$�"g�W����ۻ��i$���(�@i�:`�<�����ԭi��2�g�:Cé͓:٤yM��TI�A@3�mT �.����Jb��@ S�g�,M2��M�cM���.���6�{�Z\t�aS�x��4κ����?[��(���-��n�)p3�^h��7��)�c�3�pk%UۖT(�(�Gq�x�u.&���������v߹^z?)m�(]G�9٦t����/��`�����ib�D�i�ϹV�*%>b��i�˰�+��ՋSf���4i���Wj����B��Z��X�����6A޻��.�~�io���G�u��Xd�#�#
�XȔ�[%�cb�c����#h��vSu��;}��sCE���&����C�r5+�����[�%�Qz��Y���Zn�(>�S:p�B�%��N�oe�:�	=�" �~X#fU���o�C��Uc�E@٨�(��7$��ɼ�A�����;Մ����v�S��F������/x�^�2��,Vmo�X&?�=a����]��m���c7��Q�Izf�#'���f�6k�|m�G7��vٛ3�$$ox)��ѿ��iC�c�_�݊���o��h6`;�ΈE6�����ND�}���x�G�� ��>X�ŕ>�IA��5�}��W_wp���^�����z%�ݲ�S`��[�kL,�6���A:��VA�!V�M5�Lg@�S<�8M����J�R�#Ⱦ�r=�������\gm�p���/����e}�r��3����FH�&!t�E�hes���~����l)	���t�=�6��||�F��z��jJ�X,�k�>~fr�����-2�f{="��h���>39� V�^%r���t)R��3[�6p�QǽTV���,.{�g_�g��-�a���6�w����c(��ir=�`^�U�2����y�����8L�a�*|>XM��^�"V"J�����VH��zĔ����c��b]��xR����)��r�Ӕn�1�Ȫ��=�S�� �����^B�(�<o�SM�h/7\���H}��tL��l]"�=_"�?ki������Z�C�S5�� p�oU~�,O�6�����'	�@�1+jk~v��ƕx��c�ҿNF��>A�X��)��q�Q���4����h���	#%*,j�P*p �)ˑYA����{U���;�bS����dVG�H
ql�\%�Hi�e�k�?A�;��ݙ���d�!
p �;v��ϋU����v�KkV$N������4��q��ä@�����<60�и����V��ʿTz�4gFϰ�4�@ؕaWOI�b(�iuz��j�|�g���G#�l���@1��(� 7Đm�aJA�S�H�����
3|l��	V��W�����k����h�G�ė�[��q
�Z��fc���YRJʴU�F9-���(�]�i�;��N��_H6Q.�̃�a���U�|�*)Lel#[���B�+,�CѼ�*��8\H�b%�6?�+8�W�ȗor����e��qi��ެ��LO�zGw�i9_�b��°tݵ�=���	�c;��NV�چ\
[B]�;�2+$b�&\�d�Jz�\"��t��^�Y�Zm���>ր�F�I��d���*��������je\�X�а#?*�l"��ӟ���7���.���j��=x��"���}�{���ӫ&J�'���]@8��,�+��"�� �p��{Ǉ�����[\���	,�����X�t�ULQ�$(�3�9��3p?�D���0^���.��[���~]��w,���eM~�НrP���jH��V	�A�*Mޓ���U�g�j��?����j�nתK>KG]�.��4T�����D��o��Ւ����G�/�^Τ������WZ�R7q���4��?�t�X�`��PǦ�g���L@ڇ�|��XX|�gW:;��>��Zd�����$6+���'�m����g�����{�����Va��H��lkЕ�ӏao͜�x:n����Bn��#y֕kޱa`�s n���m?�MrR�.9�Fg�9l()O�'ab�z2 ����N�J����w�NH���2�좗���XŬA��Z��c���C�{����i!�ۇ�������{��8"� ��|��Mn��Y��.���ǮRR\�l���J�,i�^��5)`�AA�y.�N��Ƴ/���˞_�I�0�V+y,m�gp�:�NM;��s�|�K�Do�O\H|_Y�n�g�"� #���|�5���F��?�� ���4��������ta�����de��Z�e�����D�Lx�E��HV�V �M1��X�v�3AT����X4К-�Z)w��Qr�ցѱf�SJ��jN��x,��TY����]�8��������w�a7�_@�6�Q�C1Ԏo�7"��8����A��S
���*^�hA��m�h�H5�[�T/�8>c�(t/���
�5Vɶ�hlW���v����s@+oeh�����җ�u�U�JC�j�פ"y�]&�m
�:d��t���=`�v+��bd6ן���ro�
m,Bb�U��07�!˞�XIa���jBS!EI]��&��s��4Z9��«���[9�wSXj�D6C:�w9x9�N�� rz烗L:��p�U��?8fo
n�#r3c�=-�)�� �㈿�������I�IP}LoѰ��Q�v8E�\���*>`@=�f����t�ᛴ��Nk߱�%)A������NQ��,���Jڪju�g�^Mz%�4��>�M����p%0{��O�[���*�:E��Ϣ�`!���𜵸��Z��)^���xc���z)E�N�[.�sI0��2���[#Wi��5E�^o۹��i�ԉI�`?{7������dV��]<!E�
S_@�TO#�l�l�Nu�QT���J���RB�2���g��͑��j#oE�ޠeH��	*�[:#N����޺���c�ԥ�˺!��p�*4��D܃zNn��Q��<�ό�s�{x4- �����=��P�P�V�)�����L�5>xԌ�󊾜l�ֻ,I�@��Ci������F�j\�+D6R�Z����أP��5lX�[�&dhM��Q	��]m1���#�đ��>�SV�ir�[�2�0�еO�L4 ��8bij-u-%�R���~����"�}��ei�]m��²}
�i�!��t:���C�Iwh8�R�[�YvY�Ӿ4�ʩYdU�X��0U��嘃�	��N��Nz�1~�Eb����؇���`d\0	5'���/L����e�,S)��ۃ	9L�eg/��>�f��#D��o_�#j?��b�S��<"!͍��MG�Xv�HP�Ң�8qF���ļ ����٨Ha�Y���˻����W��آ��<�*��-c#�GzK��;圖���st���+m�g�-�DSi/~��ѡ����K=�B�Ղ�Z�L���G� �7����y
��
"Y�+��6ӎ�z�O�S"*�R� 6j��1��$fec5���m�XG �V���� �H��������3�W]�DGB����Hr*Գ,�B���t4D��w!��x��؛Rۖ�V*�	\��]2䶟 �ɕ������բ�#��6g�ٗ؊�<w~�bI��"l,~t�C�I�H�f��W��"p�¸ZIs��P��BH`�����f���Xh��:���h?��i�8V��i^$����P��jr����o�?�y�Df��[H�xgp���FM�X"��VO��k�O��FN@����ZQ��O�6=�%��p�sJ��Y���2�<�F����u8i)�X9���x�N½���.���RQ]��
	�����8���//"Q�1�	��c)k�!<��"�ߕ��BVC�;�{�oע͢7�j�0[&�T�BD�Mj�r�#yz�:��-),���bze+ѢJG{ئ�u����[�����Y�������������h~S����]
���F�d[|<���F}���[�N��r����Q*�>�T&�e�� ��6�ӿ�7�J��7�����u#�\�3��1�S�´l�H�z)aj�ߎJ��_+����4��!=���-J����◎��K���f7��CHK.�4�؇�3���qX2�w�A)��#�'8�� Q�W�"Z�7��.�˓	X��x�ZOH����[�c<�n�l 3��Qq^�m�}�>�����TM7�zU�3��0��vxv|�}�eIV���)��`[���$�k-Kk1w����ov��(�.���)��[��:�
�:�T�^s��l�ڝw�Fw8��A�Jwݤ�8n�E�p<w;�-�ޒ��b�D���d����0G\�	Z��̭��7��"���&Gf����]�^�e��{��^�̂��2�l�OU����q�[�y���q���B{���G�����&�d���&vu,`�N�J%n�8���;K!hĝ��-=��ʥ	uW�!���2��1�UM^���*�6�/�D�f��x�c��
���^�J�%u���X�zT�������@�!��I\m=���y$~[�%*C7���x�g��y���9"q"���$�̙�yqی�G���W@ru|K��*�d5�4��)���4�,%Y�ҵ���k��.�h<OL�	�K�}Jwes�h�j�ˬf�n�RB�:��E3�.j�����dbU$#<>��Y����"����T�e��vd��d�zF�z�1#����粜���zeqҍX=&s���*�Wr���V�w��`2����^K�"Z���B����9�Y��a���`"oSj�~F��B3,UK�񦺹�p�Oz<����r��C�O�RfH���u��9�e����3�&��}����O�m�5 r�3�@KYi;F��
���[t�5(�|�N��C%�?��	�2�ڷ�E$u`{�Q��)J@N^!�y>&5g�ü?A(��0�}�{�v5��녣&�щ�cb�&T��ջT�rk�B~.?A�ge��J5�%r��k����&w��D�J؃ ��������+y���"�Mod�\�Hj�*Z[��
;�Ei��6�V�7H{����2��ܧ�f��HH�
�~9��'.hDJ-�'9��k�!b&�P#�a�C�"�c���!Q�
���*�{�DtF�G�=�G$�����qF�,cQ]��?l���Qg�}�U��6 j0΁�����	�Lh���R�q�F$N�c#�1_��Ʈ��\���hӛ���;n�d���� "�s�>���֚0�����I,�U'�D#�.����p��󟃧Ewf��=�4�3JR;���L�A�Y5�����(x�Ӆ;ɴ�`���|N	��J	�k�N(n�t\�|�^Yט�ME�a�nx�����3�Y9zO��](I
�Л��n���i+t��V66�����-<�&W��s>��7yzD�����<�hZR�$�w�K� :�Һ/�K�� �Ƚ�S��cxR|�� <u��^M<�o�`�7����+D.�Hۊ�K=n��l���Q�.j�;��ѴP�"Ix�Z���7M ����"Y�hX��ij��� �����e �s���%������kW��
Cn��Y�]��w߁w��7`��(=����Hľ��Ӷ�mD�N�ՊD�C�BHZ��K�)*1�T	$�^�&��Q����:S�vO�R����P[��M,-�Ό�Y�6��d��!����)�}�-�B�#D�x�/(��" �+q�k�_A�[����� 8ȶ70"J�7jE�
�����h䵹�=QVĽ�@�Qv�2$墚XX�k�����<r�����(l�S������9�g��t\�k}\���Z��PhɃswŜh�<�Jp��I(��_������= �>K Jx_�i�HՀ*"��_r�A@-����D��\��0�=8X���>=�K�;8D8���M���tb�A����6o!�Eh)�G���W�K��`N�l*CTnA��`�kP�˘�����.)4�A+��z¸"�F�ޑ��k��v\P�5�~�ے:����4�ɇ�d��a��gY�U�.^`o�'��a�fH��J�,zd���)��)<�������J��7mVE�3�t瓱EhkLF�;4������ 3���|���j�	XB�^n�۫ k3JsY�v:5���	?bW}���gKֶ�,ŗ�*Mڨ�-�Eڨ���d�E�>�C�-�36�^�U�8�S��LY�Po�M{�[��Ĝ#�����]6��"�������y>�n{��*���+L��"	�/n�j�����F�QF?�5;�0�E��Q����8!YL$�9Z�8����~��nx�	]js�3n���4�8c`7��>��s�L54'QC�`�<!�y�h�i	ɴo�5|��
7t��
��H:/Y��(g�Z`��:j�T4�%�]��U8�^��>]"Ij�.�����Tp`��?��{A���,�C(��рT"c��6�L����A� �(I�9�LL�Ud����Gl��`8�1*�f #�[�{Z}F=���Jq��L��N��Cg����T���I1��APG���`Q�8�%��\N���n<}����6UOWu��:��A޸o1���7�HM���ȫ��͵������l������ ������4��R�N�4Lj/i��wٶ���(�P���_o��;��]kmmzT�*�'"�c5�1�ش����[R�K�#8x����஫?�I�-�P1�ִG��J9����'I^��#]�y�{g��f���z�A����?��
{�(<5��Z]��]��5zJ��% �
L��3�@����"�l+��2�?����������yUzpN�M+�tU�qu�,�R&I\�����K�g���h�M/�<�����B��U��hA�I�(�u�$څT�sl������f`��I�B�q���)Y-fs�!x���G��72v6~MB��9J_�� �|:}+�r�hO�T�!���A�Ч5e
��k�d,kG���A��|�Dp�4�^��"u�Ii�!�[��:Z��gDH�֜K�X8�`�8|�qՇv��v�٨�	�W�S�	0�gA�d�t����X�D��M~������C��e�N�{r~ҽ`aܫ�h���������-��|��� ߘ,�AO�J���Ȉu��b�t�)��`Unlp��=ݐ�sT�Q#:����R�B��N�r��WjhŬ-an�y�����Y�[CNe#ǸԮn����yd��a05�&@<j��q���f¨y=��7CD&0q��L
`��a�V�^d�N�v Ž��{�c�@|"�ا��? f�0knO������b�7hQԄ�_@��F!3�$t�<��0L�R|#��nA���c__A� �	�Ձ�E:��O�Բt�.Pj����J�2�Vꦆڴ�0��S�̱hy�>YnB�`8��[�f_d'�:��:-7#�1_�bzX��K�y���·7���2rJ���p�Ì��8N�� ��S^�t�kT�C�0�!��|� ��R���m���;s�I^Af���LO� 7wݨ�9@�����_�Wh��as�V|���>��I�A.������4M�廥l�n���W�ļ#�_&T�_r�W�k>�Ԥb6b
�}��T�����P����2���������y)���r�Vr�s��yɲ�B��J�T泆�܁@Z(�ȧC
l�(�G������K5l��;��R�Ж����f�b�'���%a9���p���^�n������>��l��܁�|�NP�"��h�D�A	�u���dL1�#�tP�wZZE`0ߵ ���,��?�4�"��R�	[� s�8���y(9tFG�O�(�s;����aQ"����D�uYL�d���O.�[ž0�$ �3�Z.�A��u�d�+D�Y�lߒ�\b��8��y���(|�v�P�)�Z�����kX7*�{Qx�A�]�;
�ĀH�7<���f���?5�I\�s����(�6<���xԺn��� �@�oF��ֽ����'�%�����6�	V�؁I6q��|�X�M���b�B҆���/<[p묂�	�dvuM�I-C��RYfJ�'+d�����*u�:�]��-0+�QW���4��6_W��̮�K
39s.M�71��ݢn�u	�e�2�vo찇�'�٘`�\�P��r��h�B'w�Q��2�e�	{*�n
UC�PT���@c�z�,H�z-�<�;v���1Jd���[�E�fHu��������㩍�(�͸��IyxQ�z�����9hч.�r^ӛ�ﺙm��fF�x�*v ��˕z`	�x� {Ƽ8�1�فQ}�T1�策�)Y�j��� ��	��U̪Jп�)�J_Ұ�7?"�JD�&i�:d	������3� ���4K�I���%{RIk鵙�OM��&�x�R\������Xf��^D�ϐZ�k���^_�H`r�Aw%[�	4�r���Y>�t�F�9��_�j�)��(F����2�xb�ӌԙbT)6U��^40��3�8^i�F΃����7���L|�:�M�4D[h�g��t���u�{9���d�qē�ȿ\؋����cY� �F����A��I�Ms�F���s�A�d�5�)0 S��P� �D�FJ���|�}�N�6&-����/k!�%\� �y�r���w�?𫜢 �	�h�^|�$SW��RV�:��0��VEB���&|㩴A���Z��]�̍�|z(�YJB�a�L1׹0�b�B���8{��X��$w��!sԏ�^|e_���� �hF��U�Wo��#mzb���Ɏ���I��y��KA�~#ȹ����|S2��H�"TcK&J5��	����8��a��rz']��܌���.:����\��t��T�Br�31��h��lXD�x�ۮm�̓'�LeBe4�ޠx��dJQ,k}w[���[�P�]��8�O*��f}��>��^4��ڿ�Ag�OX���$���d��>n�A��]�3�"�H<f� w�'��3r���(�:#�P����?��Wݝ	�� ަ&Q���l����	ֵڽ5�OQ�����I��S���g(�!U�}���T��>(5B��!+��j�+-���������a����W�����y���������#	=���ʲ��(���v��_ntF����W�����"�^���Cn�P�v�SFdp%�y�k��MR�����%W����_Z!}Tz����EY>�m�]��P]�gz��լ�ï���� �΄x��]��c��>�3��J���ԡ���FqK� {4C$��q��+��-@�q��u�öBK̜f�<����;+��H�V���@�j�J��)��`��.@�"G�(�{�݋�h�m.�dm�MF���fX��7��O�M���x �� ��5/%�g1��r�t����a��Lz�xK�� ��tݓ����E����6�.s0���e���.�2���z�>F#���{=3�˦����=c��M�	�Ο� c�� �dB�4	��{h5���'B��~Ӻ�?���d=�pK��5���kJ4�@࿠�����Ģ�E��o:$�q����Ls��T;*2ʇ����]�^v~�(\��6��*MF8ƙ���d�c՘��|2�6~Tn�o���~C｟���b�A����G���,���,����M�Cl�kƘل���+�J�^[p�)~��T,+p8�d�ƶ�4ʻ�ϱ��O�#~���E� C���IZ<��`�gKߵ�X1~O·��k�|a�Mh.�u�x
�fJI��3�;�F��/H�~I�t5 mVw��A4MJ"�����ʖ�2L�"{��>+E�;Ƽ-�y��#�( ϑ)9�9����Ok`��~ܽx�D��R��6�H\W��^�R��ׁ������8VeS�Wh�>x�m�4��>�ƷM���6���H�8���\0({3}�aa<�:��TfU32F�<gwP,D�X00ph{����q��g�ke�����Ƕ�I��v�3+ǽ�Cc�/Ddˁ;�8��l�c�s�X!�.L$,	ǹ�Et�%xa|j�����n��9�����;3��&xR%r!?	B�=�B����#�C)���}��I��lw�W�ۚ��mRx,u����=z%d���rTUǿS6�;	�Z`N�Ϳ��?v��C-��>fG�݇�]��ޚ�
����:�Ed*h��ž���L��L%786:_�K�fC=y���1) �_����֢�io�[f���F@�Y��@{��Ϥ�*lJ=�t�_�H��I-�H��u;k.tdj(~@��Ȕ��T�]���.3�ߣz���jTJ��N�9CC+����Q���a��jm�1��]��n��F쒕=������qJvB-�V�t
yz��x'x��J���e�'#�9� �q�ii��x��[�ëމ�G���}Y"�JB��_X��`]���aؕ���2Ԡ�~0t�j嶪+ұ��+���Ge��s�7E�l���O=a8��7M���p"�(�.l��#�H�ȇ��ɇ�>���ˢ��Da�'0eRW֧�K�$���)��âH�i�4#27sd�ƴo&-� ϗM��1�����޾�{_���$ �aG�4��.`�tCza��F��ҵo�-$���H6�����^�/|(��Pc���(%�+�u���ŕ�j�LTM{r�KJ}#X^?���bcT�b3�;�*,��'9bLF��Pc���F��� ��:|���ɴ��D�@��^��<�7�l��14��-q�o��fJ�Mp�w��ne��R9�����&�ՙ�LX,���� E
KXv��ߗ�G��zz�~�������h�����iU��5����0%�\�~nP	^O�c�i7��� 8Yak���,p��;�F����ю TΩ�Y���%q�T�жК<�2(�0��������<��'ݟl�v�\���_h%���Ҏ���PuAM���t4?M`�\�@5F�dV"��S��2���\���®��`)FJ����w���� &�1�BX�뛿ɑ�����wu�ߥ��Xf�� ������pX,�����d�N��\�ߡ�M��Z�Џc6�Or���?�Y(xQ������% \oI�͵�[n�7�W���jvLu�ټ�T��]�%b�>�����W��W�:b���<�&���P�z�5�C�U(��*a�d�C%�8��l��gI��D��Ũ��g(�bRgeCu`�L;p����v�� ?*�[:39%ut��΃������9踺R�y��NK����\��'�\���h�������&@�{4�LԽ2����ng��3h<{*�vh ��h�U`� ��r+���k#���o{�~�����{C���]�$
�#oP̏8
���g�HQ��uv�8d�/N[�,�HB��h�Ȣ:'� ��+\S�����JK�m��7�_u{� *�Q��DH;���,�颖5d����"6,H�%%="���\DЕ�&c�V)���x���:o��#R����͍�Cq��,!9ݚLƳ�,h
Q_���ק��ˢ3�)UK��o�k��|WS��X�����s����d��j-#*lRu��#��)��l0k���\�� M6��#ᅸش��=o������y��o��"��2EH+���+�ﵯ2��k� �z�z����)GEFK`V���s��(Ò#����	E0����.	��T�'��r���,��E� S~:<�岏he�������W��֏���5*��o�k�TjV'��?�	2l~����:PP=A���Z�Z�����������Y�G���F�J��3~�'5�����<�J�h�\�0��8�.�H$����=`�c�i~�2�~F�;@c��Lx���B�w-��گ�铣'B�Ց���e`G� P3��T����PH�:���;��{��(��`�Y��e�&r���g9G[��'������Zʧ��
'�����g����I2*-�����.Ǘx�<+�ؚ� n�Q� �#,Y�"������|�������:/��/0�&�!�G�v�;���-z�����H=1���"]��5S<hq�z	0�c����Š���=a$	��.���D����gN���J���M�oq�&ֹ�.p2z���ʒ�S$<�uQW�RI
Ϲ�9%̖ Q�FӞ��ދ�baj������b�ԂK�8A��YB�Pj��Ď���_��#���� ��G�&��7y��Eo�2MA��!�"E�'O�q'7\W����j��#��;�Ky�*RFܛ���T}b���-���`����7\��g@���r�</R�1(ࣀ���m�_�J�h�{V��	0s����#C����Y!������b7� �
n��}%�@�ش0[ͱ�w������O�N{X��I�m~��a�;�I�V��FǢg��ݏ\z��Xh�q�F�Y�	mJ ��G<�@�_0��T#fG���(B�P��Ζ�pX�_qo�!��⢔dR�y��+0mBi���wA.wZh���eA�g��?���&@��0� ��V����@X��N��[ۗ�Qk��7`w�9�L'^j�H�� D���Q3�屯xH-8�����V�vHV<�,�� u�&Z���nFMw��g
� ��Εl�]�噷0���u"��;wS������>%�c>c����!�o��z����U��Y+#���u��fv�ɍgr+�s���T0��-:/�I��B.7"���[7�#��P����?�����K I��2z�3`�g��q]���u3;U����'&����S���� ���R*��"X0���������i��{��.�*X��OU����d�7��u�&�/Lyw�8�U���5ϔ� n���N|k��+�N�@"�bt?�pDJ�Jk�'�?Q_��YPލڃ�3L��=ʹ�%Zb��C�m`�/J���-��0����9Z�	�o�I�J���3�T�f��D��~
k�uznY�1!�5ק���Ms����3���w���G�7C)��J���_�p�HVs��K���%
��0�=vE�ac��f�i6wVŶ���e���	Bkmࡂ����,��W�M�`��p�$w�7mH�Մ�X�q��t��^d&��ri���WGj+�Aa����(������ü�&N?��pb�ǒm�G6�CxaN>��	�W�Kw/aG65�m���?*6U�@��|I�&��S���e9	��}�)q�zb�
[���R�L���#Ը%�Fcj	�QkHb2�Ú����k_���(e�|S�9	̀vp��+���Oۈ�I�!Ĵ<T��k^]X��/���9��R���!C㭟�஝41eR�T��&x7���\uvhh;�f0��>FdM��x��e?��J�V~8`T_3���:]��I1�W-�t��`���m_��� -p�,�/ھ{�#��ke��7�=:.�dM"�9o��Y�fN��_�,QO�z��Bd�&K�XC���gfQ�e[4�}���w�} �w}�c��r�)8v�a]<bI)�l���2�(�2���qg�\��|����s��Q~�u�d�w<����N�� ���TI�s��P"`kz�&ї��غ/[�/�9j����n�A�ѐ��=ޠ$��8Ɨ0�@U-C��"��ˮ3I|��:e��s����S�.�/��=U?+h]N�Drq��#��`?��4�v۲(a�0�{�����!!R2��u�7�"e�8������5H؟y	�GK��J�JI���l���;���w�^s$�㗁%+�cӔ����h�hb*g3��*�O������'Q�+)!�]���q�_�`�p���|��h|�K��~~�S��!	X��!�FE<�ӭ�2Q��I1�'==�kY����V���E1p��wz���!�b#X���K���^ K���� U�����[H���=�Ns�QхĖ��.��H�l~�T�("P23�8M/��$y:�t~��Z���c�`P��t��/Vٓ��)�rB�q�yx��]ܡŻ�J4�FP�	�Nz���͔}���U`�Ϙ�(sgV��5�ǹ4�e�J�˿���YH��91�G<�u�/�C�
+����*����z+w�w�7#&�T���z�4!NyG)+��o�g����֜��d�흾���J({ۄ��Jg
Y(K5��w�����ӄ��U���ڭ�%����fe�7�U�����iI�ޣ�a�*��1����6Ύ���f�i1�N�Vy���F�������p�ǎ�5��l��ɷD��������%BK�����@ʪr��Z8�'���E^J���&�T/��;�{Zt[����U�#�^�4����?D�$��RF�O^�	M1}i�IV���04�3��ܭx*!N��+$�hD+� ��CB�r��/z��Ģy��w���l��� ��R}�v�J�>���:��@f�04C���������&�W�f�/��2&���*�����c)��GN��{~�b��0VOW�Z�R&˸�����'O�1)�pAAV�&�i\�3f��� �_�6�����Q��.ue��LcQq�j��{�6,S��.�m��T�'E����2�}��el����C'TT1�3. �*�oSgWgO	���'2/0�7��-ll
Jpm��I�������cB��F��f���B�ؔ�Bk��>WY���(h�t��q�&SMv��́ 3�l�X�0�T�c�:�R�qk��%�'�����Z�woI/hV��z'H:��e���s������"M\�<��l���U`���"�#�W��zL�>r.�)p�,���r��9��v���s)*����4\5E_W=j��˘�'�	%�i�y���r���dN������u������^7w�jw;30��q�J�f�*�����z"�5��z��;�'x�B��B�ϭ5H|�;�b"W�ϭ1��V\���Q�����pҔ�{�/�rK6c{	λɭ���J��K�������4AK׆:�堬hۛ����`'�����o[���\~���_T��]�~RZ�An�4��o[�C����7�[��%�2֠�kx��gծ�a�������)<�M�����������o/q ���_��*��־�r��% ��[�����1m���^6� �JⅿFy#@03�T��r|�4�`~Dj�b-�=�JV��伷rQu*}T`�$�CBG,��"��o��3�료6x���F����ߋ���rY���"
���m~Ҳ����{��z˳�fL�0/�_�۶94ƙ���>#1w�C	�R����)G"	���kg���)����}"�W��s<����\ ލ���Z?��f�0 z��f���e�a��.�7�Mm�&S�5z��^�~�d�E��s�JD�s&�8</�H�[�W�c��/}?�N�E�o���L(",HB���k�͈2�������Nb�g�3o���)7���$r�c~�з9W��e�yu�����xĩ�&I�]�z��p����� U���bJB��m���l�9��-�P=�{#c���=݂D�Iة�J���0I�ϨRKv�id4�j�l3����q��b��RJ/Oo���\r�S;�C�!���4Q�><�@Tz����&t�faX�ԴZE�6gA^�I[C�1Ԅs�����A����F�@L�������Qn�6R��0�"�R��v�����+څ��/�`�]�{��&a�>�>X�7��J]B�Q��Z~�<k�~��|O��ɕ��u�#"	�9�����u��-�\���yo�t�,Գ��y���b���!��0�~�K�-��~2�XJ=�xA%�O��1��H��?K��c�`r����\�r .[x(牾��#Kcj��靃%V��G�z;żk��p2
t�"_�5����*�<��p�֎@�Yj��;��Q��𬃩�PiO����hE*xs�5j�)�0����K,����;m���q��X�Mɮ�-��/��-G��A>�'�:h��X&o��k��v ��°��� Iw�^v=�J��<�\9��I��-*�����ֻɅ;���Pl����uqa�h�� �Y����t�M�=7�Ͷ �lc�0`���;D�b9��������|���$:B�ⲶZ2|�A�L��͗��NY1��L�'1��%�$�uF%��yn��z(I@��	*�W��q��鍌�*�2�$���7GO�'Di�4ԣ: +xQ��������R�s<Q(oiH��f��s�o��]��OҶ�E�3�����l�Ҫ ���Б���F�`�;a�7H�nzr^h5ώc1j.�_85pՒ�ݥI	�,IA'z�R���\(#��Y*����������_
�����F$ �yO���gFE"��_�#�p]�-���>i����0����.��R��U�e�q��(�C�w�%jp�� ���nu+X�&�|�]��V���J'��4NM`��&IQf�'�7B�U�:�2 :Ԛw��{y�`@�[db��ɂ��V�����{?6��	N�;_,i���=�ތN)�F'����@9� n6!�hɽ��S��LaNf<"Q�O�^�L���z�B��KEk�>��e�x9�4ăJ���vZ��m.}�!�2 jX]`�� 	+��-,%�Z���+Õ�=��Cd��X�*[#6~���q��3#,��6.��:�_��rߚJ��2�)�k���tJ9��G�.U�Q��
Y����Q?bH�|^����D=O�Namf-��τش�e0�ĈT���5.]ӣ=�U}:���+��#�)뛳�U����!�tLt(��$C^.ٿD��J��ސ��&_����k�i�
}�"�J��p�0Bۭ=pa��� !��4iߢ/�Y���B���J�?<g�y�I�1T�ܫ�6�o�`	)��,�Pc~����7_�[���æSǺc�����힉�	Cn�|w3��߰o9�{桞WU������Dۑ��r����a�"{��Sgd1����Yb�G��*!�1�9ث1���D����m�y���,�(�~y��r�w�s��.�g�h�n�+�E�E�p�eZ_A�Q��M3�E�Z.��R��RO+",���\�g������t��ժs�?C������@K����c��J�U��������UZr��%-�w��[���G�Ӟ�m��Z)ޝ"�sɎk�^��?bKlb��~JS�7 �v�'��FцY�W�{����"�����5}`}�%K��O_���j�<����%���p���v�CȚIЌ������2�gI֣!0�5׽�7b�}���;4������E3�	���Z�-1�؏���++��$9���\���
w�P���0$�;%q0�&JLqХ��fE_�3Q�V:-��r}9{��U�-�)=�::֘-���m8�z0�����/�7�<P�(�E� ad�n��	� �ث� {6����U[�ލڻX���,-M�����}YXև'��$���$,�3�4�k|����+�v5�康�Hś���T����i%�U�tV�Cv��뫳�U͂l�K�Z���.���.h�����e��#�e2V���0��wෂ��m�2c
1��c��5��]����e�gf\<�!aw��	���K��1������)�+ɳ���1�<$�V]��3q`0���+w/�U���_����ߛ6E����
�l�K�4-!���#I����΍`-Ӵ* Z��?�u���+��(@|�^��&&Z�n�0]|% �TB2�I�0��fS��TA��`y��ɮH��DG�R��QT(���#ݨ�W����u��;_Ԉۺ���B:W��=�m#����YSϴnK�#�Z��λpkT��n�#6���ޢ�I���}B#
�Ń-;��@�tBq=R�?  ��=;��Ftb!� Ą��>yO�G�����o �uND��:��M^ ����t;���^6��Umn�F)�5��z�! q�*��[�-�P�=�AA��_+9ȵ�B��_�^���<Zs����S|��F��-ҾW<"��S�,��v�e�룆G'L�� F��!֓�Up��RTEH���n|��n�L�IsƔ���V9��b��o�	O|9�&m�V̬�����[�h]�"2��r��T� ��>�M�)���J�Og���z]l�Bݶ����`�mƱd=;�X {���k�V��eD��^�[���4���+���D��󷮼��E������M�����2�lQ��ĹD�}�2���twFٹyM,u���f�q�Y00)Oһ�)���@X鯟("I�����6�w&ќ�_Mg#R��<�ˠR��BJ,;���X���0��!vv>��H�k'Ó�e���J��ڈ�ž/�PL��cc7ƥ���*�\��_kq;�2 �����J��f�hFH^�wn�D��N�@�����0��FEE֦�p���L���r<�'p^��VL��	�XU	�V@�D�ы��nfY���,�@����-jzv@x,������i�/a����p�a)�5�sM�~ �\̲��w�/��skgx�ǃ�M�Z+ɸ�񺝘���HU%*zSRᙻq8�''��qt��Z��i���$g�K�0
�`��p�
,,$Z����S��o�xtG�	�ǐ��LVy(���p2gK�0������繟d�r��=^m�U���o���g ������$�W��֞Mܱ�(Q�tZ�~��\*T��]�!7͗Q�ǰ��'�ږ%T��0�d���n�P��s��=���%=�*O����NB%C�`=@gt�	�F��KZ��&�.tT���nT��S�	�T���)UN{e)I��5�'u~��w�`�]�?t���l$@j��%�/���tȐ����.�-�'���7*�*�ĵ��9���d�R-ыJD���n�+	42�!��A�gA�<�b�w�X�i�w�W~	p�|��HQ�k���4g��fv�uߢ�~^G4�j����b�	t��S�O
����1�+U��>�m�Af�=��B�� ���݁r�ȝ¨��?|ߊg�w�ڡ���.��RA��w;�\����%I�}��xR`���p�ʲ��X~j�h�����;#��Y������^�]��AXZ�僝�	_``�c:��v'�����*f�>�A9�wN��2bd���u�������j�^��%��1��/1�g��洜�����c�Э�1�M�&H�VxK7Q�Gӏ����d�����59���1&<�����'��������t� �\�+4D��f�H��k0+ �ϑ�$�⒠c���Q��uE�6+�9�ry!\&���bcƧ�{I{Cu8e���נ �]-�����@���h/Vw��$�7�ۛx�
�yo���A7�(��1��Pi�R'#�����G�\��J C�����{�ax�@:Ù�G��9ERMť2mI�#>�Ê�z7/���j3 �ab%��Ig�]��K�H�[|�x�!B�D��%�Û'��
�=��j�7�U�"Җ;N2��4������v�w�B��	h�8�E���q�-s�9E���\��T����� ���vy��a7�R~������ � �+ �W���s�m���m��7lf�iZ5��Ŀuh~+�;�^o_}���_�8x�y������Բ8-�?��-@$�D��>03�b4�� �.�׿	���n��U}�7�¸���Q c ���s��6�J����}�:b�c0�J��p��)���tn|i�S��<	�`G����F�--67�Q�m�4ζ����򪓞Hp������F��R�{��O��Nx�l��ȋޠPh;?��ըi����akVςw>��8ހ)d���kyk��]*2�|����5����4R���8F�*?҄ȭs^��U���T*eWx/��i?	u2x	��m�t#�ƺ=�q7��g>h���v|� � a���,��k�w�G"H�#��-�V�L͠s��7�KgK�c.nI�-?�?�y�������6�h/��+V��n��5 r�;��-1#�!����v���m8�v*��h���-���c��uC%&�H=i�0�(	����TR;�/F�5�q�����(�����HP�#�cg�����w�ҳ�-�h![�8�5 "���o.����=DI��T��A� ��UZ`��Q��w:z����jVgȳ�`D�N_�d��Z��J8��a�����*/ޯ8i��A�	����!�q��LG0�ի(Ǒ���pDn�w�9yABh��G'�x��V<��Ý�����C3����֒7{xP~�q�&��ń�|H�]Ȳ��
��hi�GP异�t�.D��wv����Ls|[�5P��?�$;������$a[ӰZ���go=��΢ׄ���!Ǝ0>��d9?a>߬m�hm"��m�����fr�]ħ�H��:7���b��n�?�cR�������꒧f�<�(W �)���Pn�u�
�G�W`���!����g/�Hj~{
���y�*2 ֪���kTb�{���{��.��9�U_`�4��~7��Y3���/��ǁ��J0h8}1��O�����כ�&5���z�S����g��Cf���s��4���A�O���K͕�w2�A�z����ۊg�l�#��Xurq*YÕyV��8�l��%g�H��	�,�﮹#_�9��Qjzb�vzU>��&1�+B�P�*j���"������-|�]�#�-�g$řUD����'8Χ�a�h�>����8US�ݐ$��3�p�e���m�H����Hj-��x
�����)^|�$�+jglG�
]�"CU.�=3�n۰���� q�N�2���;����:_9بU�2����Y2HccX���χ��(�G����m�o��;眼5�d��k���g����H/���K�r]k*��sӪ�Z��(���$����yc��� �[���HJ�'��"1G���a=˽$�R~�C#�bC�ˊ �Y�8T��/O��"f�v�`U�M�U6_� ��3u��g(�ލC@�}�s�=Z�rw���C�S�h0���$��G��o'kyF]�b�� '�֏L�q�r��'�<AS��h��BiIl:1��vU}��é-w�S���,7�"��!���*!�e�zL 傞�йx $�Y�B�9Ldf�V�<�l�C���(�=�#�/��5�3N�u���ƽk�)#L�9-�%"f,���쪓�>��?�Ƶʒ�d�##Mwٸ0Ó_���pr��|<�@kV�|0��Q_c����dP?�W�!�2��Z�s�Ք�دQ���򔑿����Z�p����E��J�Np#�(��5g�n��ek D3BM��%y{�Q��rRS�j� �� s�d�M�IVh���(���{����o#!�K,��[�p��=��{z��G��R��<��	6��\4'�0h:[Bd�"�w�����x��n�L�M<�=׋RB�%M�����msl�[��J��wfi܏��i�ғ�gn�Ԭ q0X
��6�o�5�~PJ'�7�zUW�G�1�T���85ƙ��iaɻ"�O�q
|xax�Kx���ȹ����O1�I�̜��(���멇*��x��m�����f"�����3b�ks���jȒ
����O�C�"�
���=:��/��Es�Q������o��p>+���_,���u���T��^�t��Ut��h��AB��9,&����T}{�N�3���(�7�9WbU����v㫫 �Ǝ�N�u^��~ �.F�Y����� b.��[f[%>��e�2[��?6�dN�6O�����U��;{�v'E��WCN �`F�u�#/��ȃ7f�Dj�z�����N�zuٷ�X`�I;g�������|��/O[�����K�x��0ϑ�H�2|�{�q�h�wװk	��[$� I���g�����u	���W�{��]���/E~��{`1iҦ�(�q����rA�h���rb[���B� ��X�Å��p�����T���q��&T=-�-��ڞ�-�`�)=u�����A���r�}=e5ޙn|i���{���A�u�����l�Vk��^#����4�<2#T%P����\��8J��Ѡ�r;�\ؔ�r3n5���^z9IG��$v`�~�5��T���d$��AV��<'�rv�">"J831e�KRL[;�������o�D�cN>�%�Z��?礽�`�9���<��|	�> -�ᣓIڸ�b��1�V����}�j����K�M92���z�� 0|&���$������q+�%S�P�5�lO$r�?�,��EO�2)r�'sjv䗰́ZU��}J9�����0�t;���|����Up��o!G�?��l���O[������E�X����q=�CL."�5Q:I�?W��}����w�f2����D�0��m�ŔJ�?�#3gڡҩaq��G��JNܮ?���w!k���UB�02��+�P����j��w�aѧY��dǋNXj��'*늯>OVkF���%2ֽy&�
��L��~zUKA#Jl�x>�F�г]J��KpII���9���#��W6���3��o��_G���s���32{��
 �Lm��6z��'*���dE�$jb+�ݹ��}Vn,Y\�k�-�uQ������3����s�b$'��?�X��~j�r��<9,����Й�ʜ'Ǌ�h�H��yf����ü���Άu�gg��|е��f>p����-!0-��jh`!���AC&S������^��T;	�k�&�i=.�fA��9�T����9#Gf�ut����-��'��D�cܕ���B��n����%����'�4J,{XutF��)ij�Ӽ��b��B�O�}������5Y
ŗr4��W�m5�Oi�O���Aa؀p���T�k3��l�ΊSU�׵z�g��ͷ���f+���v�L�hэ��`{�ĸ�<x0��5h�%�0��ψ}�Y�����P NEON)d'��?uZ���p��?�4W2R�����y�kH=G���n�/M�Ir�L"F�(��O-@��#�+`�$6��nέh�o �̆� �*���ݹ�(f�X<�uB�ZY�	�����q�yO�8����!L����$~�$�Ru��1���	�h��[�b�ZG�^c�-K|���Hc?�1��-��������z.> �&���� ��}4e�u��V�?��0I�7O>�b��H�l�"�H{GR�9�c�ܵ�������M�����Y|rxJN �\	h,��`@��b������l����BlO�܈������8�c����P|�����Vu�C��У�P~���r�a��j�U��� ���T	'���8�	z[\^�t*��h���U������������w���!amnSro����8����eԿ�lg%��υ��;�q�����X������G��D �j߅f���~~��A1oa1�ޭ��(ۺ�75I�^�*�q���./���Z�'=�o�1F�K��b�K��(�{=��X,��M�e���}� y�}&�*9Y��'̏�ˤ6y0�m��O,_GYD���)ܨ��,�0��쉥G~=���"�RW�pY��jJ�RS��]hŴ�~��
-��}1y�?4|�ƢZ���w�/��T0��/��